VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_silife
  CLASS BLOCK ;
  FOREIGN wrapped_silife ;
  ORIGIN 0.000 0.000 ;
  SIZE 894.870 BY 905.590 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.350 0.000 294.910 4.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.140 4.000 633.340 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.990 901.590 34.550 905.590 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 827.980 894.870 829.180 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.190 901.590 43.750 905.590 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.390 901.590 328.950 905.590 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.470 0.000 466.030 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.030 901.590 367.590 905.590 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.550 901.590 833.110 905.590 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.030 0.000 275.590 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.180 4.000 380.380 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 813.020 894.870 814.220 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.540 4.000 857.740 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.590 0.000 200.150 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.990 901.590 471.550 905.590 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.750 0.000 428.310 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.510 901.590 63.070 905.590 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 109.900 894.870 111.100 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 644.380 894.870 645.580 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.550 0.000 856.110 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.660 4.000 506.860 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.150 901.590 262.710 905.590 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.910 0.000 104.470 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.020 4.000 576.220 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.220 4.000 127.420 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.030 901.590 528.590 905.590 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.350 0.000 570.910 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 770.860 894.870 772.060 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.820 4.000 549.020 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.670 0.000 38.230 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.220 4.000 365.420 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 236.380 894.870 237.580 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.830 901.590 243.390 905.590 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.910 901.590 81.470 905.590 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.190 0.000 342.750 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 901.590 671.190 905.590 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.070 901.590 585.630 905.590 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.630 901.590 234.190 905.590 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 883.740 894.870 884.940 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.510 901.590 776.070 905.590 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.100 4.000 478.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.270 901.590 709.830 905.590 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 672.940 894.870 674.140 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 702.860 4.000 704.060 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 405.020 894.870 406.220 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 0.000 95.270 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.510 0.000 799.070 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.990 901.590 195.550 905.590 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 490.700 4.000 491.900 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 209.180 894.870 210.380 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.980 4.000 183.180 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.270 901.590 433.830 905.590 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.510 901.590 339.070 905.590 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 0.000 351.950 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 0.000 257.190 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.790 0.000 761.350 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.420 4.000 562.620 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 489.340 894.870 490.540 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.870 0.000 875.430 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.230 0.000 675.790 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.300 4.000 267.500 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 546.460 894.870 547.660 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.790 0.000 209.350 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.710 901.590 348.270 905.590 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.310 901.590 766.870 905.590 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 560.060 894.870 561.260 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.630 0.000 418.190 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.070 0.000 884.630 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.270 0.000 180.830 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 194.220 894.870 195.420 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.070 901.590 424.630 905.590 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.620 4.000 759.820 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.100 4.000 70.300 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.590 901.590 453.150 905.590 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.030 0.000 827.590 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 447.180 894.870 448.380 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.310 0.000 237.870 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.900 4.000 43.100 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.350 901.590 271.910 905.590 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.430 0.000 684.990 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.500 4.000 872.700 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 475.740 894.870 476.940 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 897.340 894.870 898.540 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.470 901.590 443.030 905.590 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 659.340 894.870 660.540 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.470 901.590 719.030 905.590 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 901.590 871.750 905.590 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.670 901.590 291.230 905.590 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 167.020 894.870 168.220 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.710 901.590 624.270 905.590 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.390 901.590 880.950 905.590 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.500 4.000 464.700 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.190 0.000 779.750 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 180.620 894.870 181.820 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.390 0.000 627.950 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 901.590 157.830 905.590 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.030 0.000 551.590 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.190 0.000 66.750 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.710 901.590 72.270 905.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 320.700 894.870 321.900 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.470 0.000 190.030 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.270 0.000 732.830 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 589.980 4.000 591.180 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 885.100 4.000 886.300 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.830 901.590 519.390 905.590 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.230 901.590 652.790 905.590 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.550 0.000 143.110 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 743.660 894.870 744.860 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.150 901.590 538.710 905.590 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.630 0.000 533.190 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.870 0.000 599.430 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.070 0.000 332.630 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.390 901.590 604.950 905.590 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 504.300 894.870 505.500 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 124.860 894.870 126.060 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 901.590 310.550 905.590 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.230 901.590 100.790 905.590 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 901.590 148.630 905.590 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 687.900 4.000 689.100 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.620 4.000 351.820 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.740 4.000 238.940 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.820 4.000 141.020 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.230 0.000 836.790 4.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 617.180 894.870 618.380 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.870 0.000 47.430 4.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.300 4.000 675.500 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.550 0.000 304.110 4.000 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.870 901.590 852.430 905.590 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.910 901.590 357.470 905.590 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.630 0.000 694.190 4.000 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.470 901.590 282.030 905.590 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.660 4.000 98.860 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 264.940 894.870 266.140 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 800.780 4.000 801.980 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 855.180 894.870 856.380 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 901.590 6.030 905.590 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.460 4.000 717.660 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.190 0.000 618.750 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 0.000 742.030 4.000 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 433.580 894.870 434.780 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 901.590 481.670 905.590 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 0.000 866.230 4.000 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.710 0.000 808.270 4.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.310 901.590 490.870 905.590 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 40.540 894.870 41.740 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.420 4.000 154.620 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 54.140 894.870 55.340 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.180 4.000 788.380 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 901.590 109.990 905.590 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.020 4.000 338.220 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 0.000 132.990 4.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 0.000 476.150 4.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.790 901.590 738.350 905.590 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.230 901.590 376.790 905.590 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 531.500 894.870 532.700 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.540 4.000 211.740 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 701.500 894.870 702.700 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.790 901.590 462.350 905.590 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.900 4.000 281.100 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 901.590 129.310 905.590 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.950 901.590 253.510 905.590 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.340 4.000 830.540 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.700 4.000 661.900 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 462.140 894.870 463.340 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 517.900 894.870 519.100 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.380 4.000 815.580 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.030 901.590 804.590 905.590 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 349.260 894.870 350.460 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.670 0.000 314.230 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.390 901.590 52.950 905.590 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 901.590 700.630 905.590 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.780 4.000 393.980 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.260 4.000 112.460 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.870 0.000 323.430 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.910 0.000 656.470 4.000 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 588.620 894.870 589.820 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.950 0.000 713.510 4.000 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.340 4.000 422.540 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.230 0.000 123.790 4.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.380 4.000 169.580 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.350 901.590 547.910 905.590 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.310 0.000 513.870 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.510 0.000 247.070 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.790 0.000 485.350 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 96.300 894.870 97.500 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 898.700 4.000 899.900 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.110 0.000 504.670 4.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.430 901.590 661.990 905.590 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 0.000 647.270 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 251.340 894.870 252.540 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.590 901.590 890.150 905.590 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 138.460 894.870 139.660 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 645.740 4.000 646.940 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 728.700 894.870 729.900 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.150 0.000 722.710 4.000 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.150 901.590 814.710 905.590 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 0.000 608.630 4.000 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 901.590 576.430 905.590 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.510 0.000 86.070 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.870 901.590 24.430 905.590 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.710 0.000 371.270 4.000 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.590 901.590 177.150 905.590 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.070 0.000 171.630 4.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.590 0.000 637.150 4.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.190 901.590 595.750 905.590 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 799.420 894.870 800.620 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.190 901.590 319.750 905.590 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 901.590 186.350 905.590 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.590 901.590 614.150 905.590 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 892.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 892.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 892.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 892.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 892.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 892.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 892.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 892.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 892.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 892.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 892.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 892.400 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.310 0.000 789.870 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.510 901.590 500.070 905.590 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 25.580 894.870 26.780 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.350 901.590 823.910 905.590 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.750 901.590 681.310 905.590 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.310 901.590 214.870 905.590 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 532.860 4.000 534.060 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.110 901.590 205.670 905.590 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 419.980 894.870 421.180 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 362.860 894.870 364.060 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.950 0.000 437.510 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 293.500 894.870 294.700 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 11.980 894.870 13.180 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.110 0.000 665.670 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.630 901.590 786.190 905.590 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 785.820 894.870 787.020 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.110 0.000 389.670 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.150 0.000 561.710 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.350 0.000 846.910 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.750 901.590 405.310 905.590 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.910 0.000 380.470 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.390 0.000 75.950 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.550 901.590 557.110 905.590 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 307.100 894.870 308.300 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 686.540 894.870 687.740 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.830 0.000 266.390 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.070 901.590 861.630 905.590 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 152.060 894.870 153.260 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.500 4.000 56.700 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.060 4.000 731.260 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 0.000 523.070 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.990 0.000 218.550 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.940 4.000 28.140 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.750 0.000 704.310 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.190 0.000 894.750 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.630 901.590 510.190 905.590 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.580 4.000 196.780 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.550 901.590 120.110 905.590 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.470 901.590 167.030 905.590 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.950 901.590 138.510 905.590 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.470 0.000 29.030 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.460 4.000 309.660 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 278.540 894.870 279.740 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.430 0.000 408.990 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.990 901.590 747.550 905.590 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 870.140 894.870 871.340 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.870 901.590 300.430 905.590 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.180 4.000 618.380 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.260 4.000 520.460 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 841.580 894.870 842.780 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 842.940 4.000 844.140 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 573.660 894.870 574.860 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.140 4.000 225.340 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.060 4.000 323.260 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.670 901.590 843.230 905.590 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.950 901.590 414.510 905.590 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.110 0.000 228.670 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 391.420 894.870 392.620 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.670 0.000 590.230 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 67.740 894.870 68.940 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.020 4.000 746.220 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.670 0.000 751.230 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.030 0.000 114.590 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.590 0.000 361.150 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 222.780 894.870 223.980 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.830 901.590 795.390 905.590 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 715.100 894.870 716.300 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.990 0.000 770.550 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.860 4.000 296.060 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 377.820 894.870 379.020 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 0.000 9.710 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 757.260 894.870 758.460 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.110 901.590 757.670 905.590 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.830 0.000 818.390 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.590 901.590 729.150 905.590 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.380 4.000 407.580 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.540 4.000 449.740 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.990 0.000 494.550 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.550 0.000 580.110 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.580 4.000 604.780 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.060 4.000 85.260 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.430 901.590 385.990 905.590 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.940 4.000 436.140 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.750 0.000 152.310 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.990 0.000 57.550 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.670 901.590 567.230 905.590 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.550 901.590 396.110 905.590 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.230 0.000 399.790 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.950 901.590 690.510 905.590 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 82.700 894.870 83.900 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 772.220 4.000 773.420 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 630.780 894.870 631.980 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.950 0.000 161.510 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.150 0.000 285.710 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.070 0.000 447.630 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 602.220 894.870 603.420 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.270 0.000 456.830 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.110 901.590 642.670 905.590 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.910 901.590 633.470 905.590 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 901.590 91.590 905.590 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.510 901.590 224.070 905.590 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.830 0.000 542.390 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.700 4.000 253.900 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.670 901.590 15.230 905.590 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 890.870 335.660 894.870 336.860 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 894.555 892.245 ;
      LAYER met1 ;
        RECT 0.070 3.100 894.630 898.920 ;
      LAYER met2 ;
        RECT 0.100 901.310 5.190 901.590 ;
        RECT 6.310 901.310 14.390 901.590 ;
        RECT 15.510 901.310 23.590 901.590 ;
        RECT 24.710 901.310 33.710 901.590 ;
        RECT 34.830 901.310 42.910 901.590 ;
        RECT 44.030 901.310 52.110 901.590 ;
        RECT 53.230 901.310 62.230 901.590 ;
        RECT 63.350 901.310 71.430 901.590 ;
        RECT 72.550 901.310 80.630 901.590 ;
        RECT 81.750 901.310 90.750 901.590 ;
        RECT 91.870 901.310 99.950 901.590 ;
        RECT 101.070 901.310 109.150 901.590 ;
        RECT 110.270 901.310 119.270 901.590 ;
        RECT 120.390 901.310 128.470 901.590 ;
        RECT 129.590 901.310 137.670 901.590 ;
        RECT 138.790 901.310 147.790 901.590 ;
        RECT 148.910 901.310 156.990 901.590 ;
        RECT 158.110 901.310 166.190 901.590 ;
        RECT 167.310 901.310 176.310 901.590 ;
        RECT 177.430 901.310 185.510 901.590 ;
        RECT 186.630 901.310 194.710 901.590 ;
        RECT 195.830 901.310 204.830 901.590 ;
        RECT 205.950 901.310 214.030 901.590 ;
        RECT 215.150 901.310 223.230 901.590 ;
        RECT 224.350 901.310 233.350 901.590 ;
        RECT 234.470 901.310 242.550 901.590 ;
        RECT 243.670 901.310 252.670 901.590 ;
        RECT 253.790 901.310 261.870 901.590 ;
        RECT 262.990 901.310 271.070 901.590 ;
        RECT 272.190 901.310 281.190 901.590 ;
        RECT 282.310 901.310 290.390 901.590 ;
        RECT 291.510 901.310 299.590 901.590 ;
        RECT 300.710 901.310 309.710 901.590 ;
        RECT 310.830 901.310 318.910 901.590 ;
        RECT 320.030 901.310 328.110 901.590 ;
        RECT 329.230 901.310 338.230 901.590 ;
        RECT 339.350 901.310 347.430 901.590 ;
        RECT 348.550 901.310 356.630 901.590 ;
        RECT 357.750 901.310 366.750 901.590 ;
        RECT 367.870 901.310 375.950 901.590 ;
        RECT 377.070 901.310 385.150 901.590 ;
        RECT 386.270 901.310 395.270 901.590 ;
        RECT 396.390 901.310 404.470 901.590 ;
        RECT 405.590 901.310 413.670 901.590 ;
        RECT 414.790 901.310 423.790 901.590 ;
        RECT 424.910 901.310 432.990 901.590 ;
        RECT 434.110 901.310 442.190 901.590 ;
        RECT 443.310 901.310 452.310 901.590 ;
        RECT 453.430 901.310 461.510 901.590 ;
        RECT 462.630 901.310 470.710 901.590 ;
        RECT 471.830 901.310 480.830 901.590 ;
        RECT 481.950 901.310 490.030 901.590 ;
        RECT 491.150 901.310 499.230 901.590 ;
        RECT 500.350 901.310 509.350 901.590 ;
        RECT 510.470 901.310 518.550 901.590 ;
        RECT 519.670 901.310 527.750 901.590 ;
        RECT 528.870 901.310 537.870 901.590 ;
        RECT 538.990 901.310 547.070 901.590 ;
        RECT 548.190 901.310 556.270 901.590 ;
        RECT 557.390 901.310 566.390 901.590 ;
        RECT 567.510 901.310 575.590 901.590 ;
        RECT 576.710 901.310 584.790 901.590 ;
        RECT 585.910 901.310 594.910 901.590 ;
        RECT 596.030 901.310 604.110 901.590 ;
        RECT 605.230 901.310 613.310 901.590 ;
        RECT 614.430 901.310 623.430 901.590 ;
        RECT 624.550 901.310 632.630 901.590 ;
        RECT 633.750 901.310 641.830 901.590 ;
        RECT 642.950 901.310 651.950 901.590 ;
        RECT 653.070 901.310 661.150 901.590 ;
        RECT 662.270 901.310 670.350 901.590 ;
        RECT 671.470 901.310 680.470 901.590 ;
        RECT 681.590 901.310 689.670 901.590 ;
        RECT 690.790 901.310 699.790 901.590 ;
        RECT 700.910 901.310 708.990 901.590 ;
        RECT 710.110 901.310 718.190 901.590 ;
        RECT 719.310 901.310 728.310 901.590 ;
        RECT 729.430 901.310 737.510 901.590 ;
        RECT 738.630 901.310 746.710 901.590 ;
        RECT 747.830 901.310 756.830 901.590 ;
        RECT 757.950 901.310 766.030 901.590 ;
        RECT 767.150 901.310 775.230 901.590 ;
        RECT 776.350 901.310 785.350 901.590 ;
        RECT 786.470 901.310 794.550 901.590 ;
        RECT 795.670 901.310 803.750 901.590 ;
        RECT 804.870 901.310 813.870 901.590 ;
        RECT 814.990 901.310 823.070 901.590 ;
        RECT 824.190 901.310 832.270 901.590 ;
        RECT 833.390 901.310 842.390 901.590 ;
        RECT 843.510 901.310 851.590 901.590 ;
        RECT 852.710 901.310 860.790 901.590 ;
        RECT 861.910 901.310 870.910 901.590 ;
        RECT 872.030 901.310 880.110 901.590 ;
        RECT 881.230 901.310 889.310 901.590 ;
        RECT 890.430 901.310 894.600 901.590 ;
        RECT 0.100 4.280 894.600 901.310 ;
        RECT 0.790 2.875 8.870 4.280 ;
        RECT 9.990 2.875 18.070 4.280 ;
        RECT 19.190 2.875 28.190 4.280 ;
        RECT 29.310 2.875 37.390 4.280 ;
        RECT 38.510 2.875 46.590 4.280 ;
        RECT 47.710 2.875 56.710 4.280 ;
        RECT 57.830 2.875 65.910 4.280 ;
        RECT 67.030 2.875 75.110 4.280 ;
        RECT 76.230 2.875 85.230 4.280 ;
        RECT 86.350 2.875 94.430 4.280 ;
        RECT 95.550 2.875 103.630 4.280 ;
        RECT 104.750 2.875 113.750 4.280 ;
        RECT 114.870 2.875 122.950 4.280 ;
        RECT 124.070 2.875 132.150 4.280 ;
        RECT 133.270 2.875 142.270 4.280 ;
        RECT 143.390 2.875 151.470 4.280 ;
        RECT 152.590 2.875 160.670 4.280 ;
        RECT 161.790 2.875 170.790 4.280 ;
        RECT 171.910 2.875 179.990 4.280 ;
        RECT 181.110 2.875 189.190 4.280 ;
        RECT 190.310 2.875 199.310 4.280 ;
        RECT 200.430 2.875 208.510 4.280 ;
        RECT 209.630 2.875 217.710 4.280 ;
        RECT 218.830 2.875 227.830 4.280 ;
        RECT 228.950 2.875 237.030 4.280 ;
        RECT 238.150 2.875 246.230 4.280 ;
        RECT 247.350 2.875 256.350 4.280 ;
        RECT 257.470 2.875 265.550 4.280 ;
        RECT 266.670 2.875 274.750 4.280 ;
        RECT 275.870 2.875 284.870 4.280 ;
        RECT 285.990 2.875 294.070 4.280 ;
        RECT 295.190 2.875 303.270 4.280 ;
        RECT 304.390 2.875 313.390 4.280 ;
        RECT 314.510 2.875 322.590 4.280 ;
        RECT 323.710 2.875 331.790 4.280 ;
        RECT 332.910 2.875 341.910 4.280 ;
        RECT 343.030 2.875 351.110 4.280 ;
        RECT 352.230 2.875 360.310 4.280 ;
        RECT 361.430 2.875 370.430 4.280 ;
        RECT 371.550 2.875 379.630 4.280 ;
        RECT 380.750 2.875 388.830 4.280 ;
        RECT 389.950 2.875 398.950 4.280 ;
        RECT 400.070 2.875 408.150 4.280 ;
        RECT 409.270 2.875 417.350 4.280 ;
        RECT 418.470 2.875 427.470 4.280 ;
        RECT 428.590 2.875 436.670 4.280 ;
        RECT 437.790 2.875 446.790 4.280 ;
        RECT 447.910 2.875 455.990 4.280 ;
        RECT 457.110 2.875 465.190 4.280 ;
        RECT 466.310 2.875 475.310 4.280 ;
        RECT 476.430 2.875 484.510 4.280 ;
        RECT 485.630 2.875 493.710 4.280 ;
        RECT 494.830 2.875 503.830 4.280 ;
        RECT 504.950 2.875 513.030 4.280 ;
        RECT 514.150 2.875 522.230 4.280 ;
        RECT 523.350 2.875 532.350 4.280 ;
        RECT 533.470 2.875 541.550 4.280 ;
        RECT 542.670 2.875 550.750 4.280 ;
        RECT 551.870 2.875 560.870 4.280 ;
        RECT 561.990 2.875 570.070 4.280 ;
        RECT 571.190 2.875 579.270 4.280 ;
        RECT 580.390 2.875 589.390 4.280 ;
        RECT 590.510 2.875 598.590 4.280 ;
        RECT 599.710 2.875 607.790 4.280 ;
        RECT 608.910 2.875 617.910 4.280 ;
        RECT 619.030 2.875 627.110 4.280 ;
        RECT 628.230 2.875 636.310 4.280 ;
        RECT 637.430 2.875 646.430 4.280 ;
        RECT 647.550 2.875 655.630 4.280 ;
        RECT 656.750 2.875 664.830 4.280 ;
        RECT 665.950 2.875 674.950 4.280 ;
        RECT 676.070 2.875 684.150 4.280 ;
        RECT 685.270 2.875 693.350 4.280 ;
        RECT 694.470 2.875 703.470 4.280 ;
        RECT 704.590 2.875 712.670 4.280 ;
        RECT 713.790 2.875 721.870 4.280 ;
        RECT 722.990 2.875 731.990 4.280 ;
        RECT 733.110 2.875 741.190 4.280 ;
        RECT 742.310 2.875 750.390 4.280 ;
        RECT 751.510 2.875 760.510 4.280 ;
        RECT 761.630 2.875 769.710 4.280 ;
        RECT 770.830 2.875 778.910 4.280 ;
        RECT 780.030 2.875 789.030 4.280 ;
        RECT 790.150 2.875 798.230 4.280 ;
        RECT 799.350 2.875 807.430 4.280 ;
        RECT 808.550 2.875 817.550 4.280 ;
        RECT 818.670 2.875 826.750 4.280 ;
        RECT 827.870 2.875 835.950 4.280 ;
        RECT 837.070 2.875 846.070 4.280 ;
        RECT 847.190 2.875 855.270 4.280 ;
        RECT 856.390 2.875 865.390 4.280 ;
        RECT 866.510 2.875 874.590 4.280 ;
        RECT 875.710 2.875 883.790 4.280 ;
        RECT 884.910 2.875 893.910 4.280 ;
      LAYER met3 ;
        RECT 2.365 896.940 890.470 898.105 ;
        RECT 2.365 886.700 891.170 896.940 ;
        RECT 4.400 885.340 891.170 886.700 ;
        RECT 4.400 884.700 890.470 885.340 ;
        RECT 2.365 883.340 890.470 884.700 ;
        RECT 2.365 873.100 891.170 883.340 ;
        RECT 4.400 871.740 891.170 873.100 ;
        RECT 4.400 871.100 890.470 871.740 ;
        RECT 2.365 869.740 890.470 871.100 ;
        RECT 2.365 858.140 891.170 869.740 ;
        RECT 4.400 856.780 891.170 858.140 ;
        RECT 4.400 856.140 890.470 856.780 ;
        RECT 2.365 854.780 890.470 856.140 ;
        RECT 2.365 844.540 891.170 854.780 ;
        RECT 4.400 843.180 891.170 844.540 ;
        RECT 4.400 842.540 890.470 843.180 ;
        RECT 2.365 841.180 890.470 842.540 ;
        RECT 2.365 830.940 891.170 841.180 ;
        RECT 4.400 829.580 891.170 830.940 ;
        RECT 4.400 828.940 890.470 829.580 ;
        RECT 2.365 827.580 890.470 828.940 ;
        RECT 2.365 815.980 891.170 827.580 ;
        RECT 4.400 814.620 891.170 815.980 ;
        RECT 4.400 813.980 890.470 814.620 ;
        RECT 2.365 812.620 890.470 813.980 ;
        RECT 2.365 802.380 891.170 812.620 ;
        RECT 4.400 801.020 891.170 802.380 ;
        RECT 4.400 800.380 890.470 801.020 ;
        RECT 2.365 799.020 890.470 800.380 ;
        RECT 2.365 788.780 891.170 799.020 ;
        RECT 4.400 787.420 891.170 788.780 ;
        RECT 4.400 786.780 890.470 787.420 ;
        RECT 2.365 785.420 890.470 786.780 ;
        RECT 2.365 773.820 891.170 785.420 ;
        RECT 4.400 772.460 891.170 773.820 ;
        RECT 4.400 771.820 890.470 772.460 ;
        RECT 2.365 770.460 890.470 771.820 ;
        RECT 2.365 760.220 891.170 770.460 ;
        RECT 4.400 758.860 891.170 760.220 ;
        RECT 4.400 758.220 890.470 758.860 ;
        RECT 2.365 756.860 890.470 758.220 ;
        RECT 2.365 746.620 891.170 756.860 ;
        RECT 4.400 745.260 891.170 746.620 ;
        RECT 4.400 744.620 890.470 745.260 ;
        RECT 2.365 743.260 890.470 744.620 ;
        RECT 2.365 731.660 891.170 743.260 ;
        RECT 4.400 730.300 891.170 731.660 ;
        RECT 4.400 729.660 890.470 730.300 ;
        RECT 2.365 728.300 890.470 729.660 ;
        RECT 2.365 718.060 891.170 728.300 ;
        RECT 4.400 716.700 891.170 718.060 ;
        RECT 4.400 716.060 890.470 716.700 ;
        RECT 2.365 714.700 890.470 716.060 ;
        RECT 2.365 704.460 891.170 714.700 ;
        RECT 4.400 703.100 891.170 704.460 ;
        RECT 4.400 702.460 890.470 703.100 ;
        RECT 2.365 701.100 890.470 702.460 ;
        RECT 2.365 689.500 891.170 701.100 ;
        RECT 4.400 688.140 891.170 689.500 ;
        RECT 4.400 687.500 890.470 688.140 ;
        RECT 2.365 686.140 890.470 687.500 ;
        RECT 2.365 675.900 891.170 686.140 ;
        RECT 4.400 674.540 891.170 675.900 ;
        RECT 4.400 673.900 890.470 674.540 ;
        RECT 2.365 672.540 890.470 673.900 ;
        RECT 2.365 662.300 891.170 672.540 ;
        RECT 4.400 660.940 891.170 662.300 ;
        RECT 4.400 660.300 890.470 660.940 ;
        RECT 2.365 658.940 890.470 660.300 ;
        RECT 2.365 647.340 891.170 658.940 ;
        RECT 4.400 645.980 891.170 647.340 ;
        RECT 4.400 645.340 890.470 645.980 ;
        RECT 2.365 643.980 890.470 645.340 ;
        RECT 2.365 633.740 891.170 643.980 ;
        RECT 4.400 632.380 891.170 633.740 ;
        RECT 4.400 631.740 890.470 632.380 ;
        RECT 2.365 630.380 890.470 631.740 ;
        RECT 2.365 618.780 891.170 630.380 ;
        RECT 4.400 616.780 890.470 618.780 ;
        RECT 2.365 605.180 891.170 616.780 ;
        RECT 4.400 603.820 891.170 605.180 ;
        RECT 4.400 603.180 890.470 603.820 ;
        RECT 2.365 601.820 890.470 603.180 ;
        RECT 2.365 591.580 891.170 601.820 ;
        RECT 4.400 590.220 891.170 591.580 ;
        RECT 4.400 589.580 890.470 590.220 ;
        RECT 2.365 588.220 890.470 589.580 ;
        RECT 2.365 576.620 891.170 588.220 ;
        RECT 4.400 575.260 891.170 576.620 ;
        RECT 4.400 574.620 890.470 575.260 ;
        RECT 2.365 573.260 890.470 574.620 ;
        RECT 2.365 563.020 891.170 573.260 ;
        RECT 4.400 561.660 891.170 563.020 ;
        RECT 4.400 561.020 890.470 561.660 ;
        RECT 2.365 559.660 890.470 561.020 ;
        RECT 2.365 549.420 891.170 559.660 ;
        RECT 4.400 548.060 891.170 549.420 ;
        RECT 4.400 547.420 890.470 548.060 ;
        RECT 2.365 546.060 890.470 547.420 ;
        RECT 2.365 534.460 891.170 546.060 ;
        RECT 4.400 533.100 891.170 534.460 ;
        RECT 4.400 532.460 890.470 533.100 ;
        RECT 2.365 531.100 890.470 532.460 ;
        RECT 2.365 520.860 891.170 531.100 ;
        RECT 4.400 519.500 891.170 520.860 ;
        RECT 4.400 518.860 890.470 519.500 ;
        RECT 2.365 517.500 890.470 518.860 ;
        RECT 2.365 507.260 891.170 517.500 ;
        RECT 4.400 505.900 891.170 507.260 ;
        RECT 4.400 505.260 890.470 505.900 ;
        RECT 2.365 503.900 890.470 505.260 ;
        RECT 2.365 492.300 891.170 503.900 ;
        RECT 4.400 490.940 891.170 492.300 ;
        RECT 4.400 490.300 890.470 490.940 ;
        RECT 2.365 488.940 890.470 490.300 ;
        RECT 2.365 478.700 891.170 488.940 ;
        RECT 4.400 477.340 891.170 478.700 ;
        RECT 4.400 476.700 890.470 477.340 ;
        RECT 2.365 475.340 890.470 476.700 ;
        RECT 2.365 465.100 891.170 475.340 ;
        RECT 4.400 463.740 891.170 465.100 ;
        RECT 4.400 463.100 890.470 463.740 ;
        RECT 2.365 461.740 890.470 463.100 ;
        RECT 2.365 450.140 891.170 461.740 ;
        RECT 4.400 448.780 891.170 450.140 ;
        RECT 4.400 448.140 890.470 448.780 ;
        RECT 2.365 446.780 890.470 448.140 ;
        RECT 2.365 436.540 891.170 446.780 ;
        RECT 4.400 435.180 891.170 436.540 ;
        RECT 4.400 434.540 890.470 435.180 ;
        RECT 2.365 433.180 890.470 434.540 ;
        RECT 2.365 422.940 891.170 433.180 ;
        RECT 4.400 421.580 891.170 422.940 ;
        RECT 4.400 420.940 890.470 421.580 ;
        RECT 2.365 419.580 890.470 420.940 ;
        RECT 2.365 407.980 891.170 419.580 ;
        RECT 4.400 406.620 891.170 407.980 ;
        RECT 4.400 405.980 890.470 406.620 ;
        RECT 2.365 404.620 890.470 405.980 ;
        RECT 2.365 394.380 891.170 404.620 ;
        RECT 4.400 393.020 891.170 394.380 ;
        RECT 4.400 392.380 890.470 393.020 ;
        RECT 2.365 391.020 890.470 392.380 ;
        RECT 2.365 380.780 891.170 391.020 ;
        RECT 4.400 379.420 891.170 380.780 ;
        RECT 4.400 378.780 890.470 379.420 ;
        RECT 2.365 377.420 890.470 378.780 ;
        RECT 2.365 365.820 891.170 377.420 ;
        RECT 4.400 364.460 891.170 365.820 ;
        RECT 4.400 363.820 890.470 364.460 ;
        RECT 2.365 362.460 890.470 363.820 ;
        RECT 2.365 352.220 891.170 362.460 ;
        RECT 4.400 350.860 891.170 352.220 ;
        RECT 4.400 350.220 890.470 350.860 ;
        RECT 2.365 348.860 890.470 350.220 ;
        RECT 2.365 338.620 891.170 348.860 ;
        RECT 4.400 337.260 891.170 338.620 ;
        RECT 4.400 336.620 890.470 337.260 ;
        RECT 2.365 335.260 890.470 336.620 ;
        RECT 2.365 323.660 891.170 335.260 ;
        RECT 4.400 322.300 891.170 323.660 ;
        RECT 4.400 321.660 890.470 322.300 ;
        RECT 2.365 320.300 890.470 321.660 ;
        RECT 2.365 310.060 891.170 320.300 ;
        RECT 4.400 308.700 891.170 310.060 ;
        RECT 4.400 308.060 890.470 308.700 ;
        RECT 2.365 306.700 890.470 308.060 ;
        RECT 2.365 296.460 891.170 306.700 ;
        RECT 4.400 295.100 891.170 296.460 ;
        RECT 4.400 294.460 890.470 295.100 ;
        RECT 2.365 293.100 890.470 294.460 ;
        RECT 2.365 281.500 891.170 293.100 ;
        RECT 4.400 280.140 891.170 281.500 ;
        RECT 4.400 279.500 890.470 280.140 ;
        RECT 2.365 278.140 890.470 279.500 ;
        RECT 2.365 267.900 891.170 278.140 ;
        RECT 4.400 266.540 891.170 267.900 ;
        RECT 4.400 265.900 890.470 266.540 ;
        RECT 2.365 264.540 890.470 265.900 ;
        RECT 2.365 254.300 891.170 264.540 ;
        RECT 4.400 252.940 891.170 254.300 ;
        RECT 4.400 252.300 890.470 252.940 ;
        RECT 2.365 250.940 890.470 252.300 ;
        RECT 2.365 239.340 891.170 250.940 ;
        RECT 4.400 237.980 891.170 239.340 ;
        RECT 4.400 237.340 890.470 237.980 ;
        RECT 2.365 235.980 890.470 237.340 ;
        RECT 2.365 225.740 891.170 235.980 ;
        RECT 4.400 224.380 891.170 225.740 ;
        RECT 4.400 223.740 890.470 224.380 ;
        RECT 2.365 222.380 890.470 223.740 ;
        RECT 2.365 212.140 891.170 222.380 ;
        RECT 4.400 210.780 891.170 212.140 ;
        RECT 4.400 210.140 890.470 210.780 ;
        RECT 2.365 208.780 890.470 210.140 ;
        RECT 2.365 197.180 891.170 208.780 ;
        RECT 4.400 195.820 891.170 197.180 ;
        RECT 4.400 195.180 890.470 195.820 ;
        RECT 2.365 193.820 890.470 195.180 ;
        RECT 2.365 183.580 891.170 193.820 ;
        RECT 4.400 182.220 891.170 183.580 ;
        RECT 4.400 181.580 890.470 182.220 ;
        RECT 2.365 180.220 890.470 181.580 ;
        RECT 2.365 169.980 891.170 180.220 ;
        RECT 4.400 168.620 891.170 169.980 ;
        RECT 4.400 167.980 890.470 168.620 ;
        RECT 2.365 166.620 890.470 167.980 ;
        RECT 2.365 155.020 891.170 166.620 ;
        RECT 4.400 153.660 891.170 155.020 ;
        RECT 4.400 153.020 890.470 153.660 ;
        RECT 2.365 151.660 890.470 153.020 ;
        RECT 2.365 141.420 891.170 151.660 ;
        RECT 4.400 140.060 891.170 141.420 ;
        RECT 4.400 139.420 890.470 140.060 ;
        RECT 2.365 138.060 890.470 139.420 ;
        RECT 2.365 127.820 891.170 138.060 ;
        RECT 4.400 126.460 891.170 127.820 ;
        RECT 4.400 125.820 890.470 126.460 ;
        RECT 2.365 124.460 890.470 125.820 ;
        RECT 2.365 112.860 891.170 124.460 ;
        RECT 4.400 111.500 891.170 112.860 ;
        RECT 4.400 110.860 890.470 111.500 ;
        RECT 2.365 109.500 890.470 110.860 ;
        RECT 2.365 99.260 891.170 109.500 ;
        RECT 4.400 97.900 891.170 99.260 ;
        RECT 4.400 97.260 890.470 97.900 ;
        RECT 2.365 95.900 890.470 97.260 ;
        RECT 2.365 85.660 891.170 95.900 ;
        RECT 4.400 84.300 891.170 85.660 ;
        RECT 4.400 83.660 890.470 84.300 ;
        RECT 2.365 82.300 890.470 83.660 ;
        RECT 2.365 70.700 891.170 82.300 ;
        RECT 4.400 69.340 891.170 70.700 ;
        RECT 4.400 68.700 890.470 69.340 ;
        RECT 2.365 67.340 890.470 68.700 ;
        RECT 2.365 57.100 891.170 67.340 ;
        RECT 4.400 55.740 891.170 57.100 ;
        RECT 4.400 55.100 890.470 55.740 ;
        RECT 2.365 53.740 890.470 55.100 ;
        RECT 2.365 43.500 891.170 53.740 ;
        RECT 4.400 42.140 891.170 43.500 ;
        RECT 4.400 41.500 890.470 42.140 ;
        RECT 2.365 40.140 890.470 41.500 ;
        RECT 2.365 28.540 891.170 40.140 ;
        RECT 4.400 27.180 891.170 28.540 ;
        RECT 4.400 26.540 890.470 27.180 ;
        RECT 2.365 25.180 890.470 26.540 ;
        RECT 2.365 14.940 891.170 25.180 ;
        RECT 4.400 13.580 891.170 14.940 ;
        RECT 4.400 12.940 890.470 13.580 ;
        RECT 2.365 11.580 890.470 12.940 ;
        RECT 2.365 2.895 891.170 11.580 ;
      LAYER met4 ;
        RECT 4.895 10.240 20.640 891.305 ;
        RECT 23.040 10.240 97.440 891.305 ;
        RECT 99.840 10.240 174.240 891.305 ;
        RECT 176.640 10.240 251.040 891.305 ;
        RECT 253.440 10.240 327.840 891.305 ;
        RECT 330.240 10.240 404.640 891.305 ;
        RECT 407.040 10.240 481.440 891.305 ;
        RECT 483.840 10.240 558.240 891.305 ;
        RECT 560.640 10.240 635.040 891.305 ;
        RECT 637.440 10.240 711.840 891.305 ;
        RECT 714.240 10.240 788.640 891.305 ;
        RECT 791.040 10.240 865.440 891.305 ;
        RECT 867.840 10.240 882.905 891.305 ;
        RECT 4.895 4.935 882.905 10.240 ;
  END
END wrapped_silife
END LIBRARY

