VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_openram_wrapper
  CLASS BLOCK ;
  FOREIGN wb_openram_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 400.000 ;
  PIN ram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END ram_addr0[0]
  PIN ram_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END ram_addr0[1]
  PIN ram_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END ram_addr0[2]
  PIN ram_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END ram_addr0[3]
  PIN ram_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END ram_addr0[4]
  PIN ram_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END ram_addr0[5]
  PIN ram_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END ram_addr0[6]
  PIN ram_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END ram_addr0[7]
  PIN ram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END ram_addr1[0]
  PIN ram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END ram_addr1[1]
  PIN ram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END ram_addr1[2]
  PIN ram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END ram_addr1[3]
  PIN ram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END ram_addr1[4]
  PIN ram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END ram_addr1[5]
  PIN ram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END ram_addr1[6]
  PIN ram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END ram_addr1[7]
  PIN ram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END ram_clk0
  PIN ram_clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END ram_clk1
  PIN ram_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END ram_csb0
  PIN ram_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END ram_csb1
  PIN ram_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END ram_din0[0]
  PIN ram_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END ram_din0[10]
  PIN ram_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END ram_din0[11]
  PIN ram_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END ram_din0[12]
  PIN ram_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END ram_din0[13]
  PIN ram_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END ram_din0[14]
  PIN ram_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END ram_din0[15]
  PIN ram_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END ram_din0[16]
  PIN ram_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END ram_din0[17]
  PIN ram_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END ram_din0[18]
  PIN ram_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END ram_din0[19]
  PIN ram_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END ram_din0[1]
  PIN ram_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END ram_din0[20]
  PIN ram_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END ram_din0[21]
  PIN ram_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END ram_din0[22]
  PIN ram_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END ram_din0[23]
  PIN ram_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END ram_din0[24]
  PIN ram_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END ram_din0[25]
  PIN ram_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END ram_din0[26]
  PIN ram_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END ram_din0[27]
  PIN ram_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END ram_din0[28]
  PIN ram_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END ram_din0[29]
  PIN ram_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END ram_din0[2]
  PIN ram_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END ram_din0[30]
  PIN ram_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END ram_din0[31]
  PIN ram_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END ram_din0[3]
  PIN ram_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END ram_din0[4]
  PIN ram_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END ram_din0[5]
  PIN ram_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END ram_din0[6]
  PIN ram_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END ram_din0[7]
  PIN ram_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END ram_din0[8]
  PIN ram_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END ram_din0[9]
  PIN ram_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END ram_dout0[0]
  PIN ram_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END ram_dout0[10]
  PIN ram_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END ram_dout0[11]
  PIN ram_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END ram_dout0[12]
  PIN ram_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END ram_dout0[13]
  PIN ram_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END ram_dout0[14]
  PIN ram_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END ram_dout0[15]
  PIN ram_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END ram_dout0[16]
  PIN ram_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END ram_dout0[17]
  PIN ram_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END ram_dout0[18]
  PIN ram_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END ram_dout0[19]
  PIN ram_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END ram_dout0[1]
  PIN ram_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END ram_dout0[20]
  PIN ram_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END ram_dout0[21]
  PIN ram_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END ram_dout0[22]
  PIN ram_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END ram_dout0[23]
  PIN ram_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END ram_dout0[24]
  PIN ram_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END ram_dout0[25]
  PIN ram_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END ram_dout0[26]
  PIN ram_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END ram_dout0[27]
  PIN ram_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END ram_dout0[28]
  PIN ram_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END ram_dout0[29]
  PIN ram_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END ram_dout0[2]
  PIN ram_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END ram_dout0[30]
  PIN ram_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END ram_dout0[31]
  PIN ram_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END ram_dout0[3]
  PIN ram_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END ram_dout0[4]
  PIN ram_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END ram_dout0[5]
  PIN ram_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END ram_dout0[6]
  PIN ram_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END ram_dout0[7]
  PIN ram_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END ram_dout0[8]
  PIN ram_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END ram_dout0[9]
  PIN ram_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END ram_dout1[0]
  PIN ram_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END ram_dout1[10]
  PIN ram_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END ram_dout1[11]
  PIN ram_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END ram_dout1[12]
  PIN ram_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END ram_dout1[13]
  PIN ram_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END ram_dout1[14]
  PIN ram_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END ram_dout1[15]
  PIN ram_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END ram_dout1[16]
  PIN ram_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END ram_dout1[17]
  PIN ram_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END ram_dout1[18]
  PIN ram_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END ram_dout1[19]
  PIN ram_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END ram_dout1[1]
  PIN ram_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END ram_dout1[20]
  PIN ram_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END ram_dout1[21]
  PIN ram_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END ram_dout1[22]
  PIN ram_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END ram_dout1[23]
  PIN ram_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END ram_dout1[24]
  PIN ram_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END ram_dout1[25]
  PIN ram_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END ram_dout1[26]
  PIN ram_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END ram_dout1[27]
  PIN ram_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END ram_dout1[28]
  PIN ram_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END ram_dout1[29]
  PIN ram_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END ram_dout1[2]
  PIN ram_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END ram_dout1[30]
  PIN ram_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END ram_dout1[31]
  PIN ram_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END ram_dout1[3]
  PIN ram_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END ram_dout1[4]
  PIN ram_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END ram_dout1[5]
  PIN ram_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END ram_dout1[6]
  PIN ram_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END ram_dout1[7]
  PIN ram_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END ram_dout1[8]
  PIN ram_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END ram_dout1[9]
  PIN ram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END ram_web0
  PIN ram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END ram_wmask0[0]
  PIN ram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END ram_wmask0[1]
  PIN ram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END ram_wmask0[2]
  PIN ram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END ram_wmask0[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 12.875 10.640 14.475 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.195 10.640 30.795 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.515 10.640 47.115 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.035 10.640 22.635 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.355 10.640 38.955 389.200 ;
    END
  END vssd1
  PIN wb_a_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 2.760 60.000 3.360 ;
    END
  END wb_a_clk_i
  PIN wb_a_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 4.800 60.000 5.400 ;
    END
  END wb_a_rst_i
  PIN wb_b_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 201.320 60.000 201.920 ;
    END
  END wb_b_clk_i
  PIN wb_b_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 204.040 60.000 204.640 ;
    END
  END wb_b_rst_i
  PIN wbs_a_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 14.320 60.000 14.920 ;
    END
  END wbs_a_ack_o
  PIN wbs_a_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 26.560 60.000 27.160 ;
    END
  END wbs_a_adr_i[0]
  PIN wbs_a_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 28.600 60.000 29.200 ;
    END
  END wbs_a_adr_i[1]
  PIN wbs_a_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 31.320 60.000 31.920 ;
    END
  END wbs_a_adr_i[2]
  PIN wbs_a_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 33.360 60.000 33.960 ;
    END
  END wbs_a_adr_i[3]
  PIN wbs_a_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 36.080 60.000 36.680 ;
    END
  END wbs_a_adr_i[4]
  PIN wbs_a_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 38.120 60.000 38.720 ;
    END
  END wbs_a_adr_i[5]
  PIN wbs_a_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 40.840 60.000 41.440 ;
    END
  END wbs_a_adr_i[6]
  PIN wbs_a_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 42.880 60.000 43.480 ;
    END
  END wbs_a_adr_i[7]
  PIN wbs_a_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 45.600 60.000 46.200 ;
    END
  END wbs_a_adr_i[8]
  PIN wbs_a_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 47.640 60.000 48.240 ;
    END
  END wbs_a_adr_i[9]
  PIN wbs_a_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 9.560 60.000 10.160 ;
    END
  END wbs_a_cyc_i
  PIN wbs_a_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 50.360 60.000 50.960 ;
    END
  END wbs_a_dat_i[0]
  PIN wbs_a_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 73.480 60.000 74.080 ;
    END
  END wbs_a_dat_i[10]
  PIN wbs_a_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 76.200 60.000 76.800 ;
    END
  END wbs_a_dat_i[11]
  PIN wbs_a_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 78.240 60.000 78.840 ;
    END
  END wbs_a_dat_i[12]
  PIN wbs_a_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 80.960 60.000 81.560 ;
    END
  END wbs_a_dat_i[13]
  PIN wbs_a_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 83.000 60.000 83.600 ;
    END
  END wbs_a_dat_i[14]
  PIN wbs_a_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 85.720 60.000 86.320 ;
    END
  END wbs_a_dat_i[15]
  PIN wbs_a_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 87.760 60.000 88.360 ;
    END
  END wbs_a_dat_i[16]
  PIN wbs_a_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 90.480 60.000 91.080 ;
    END
  END wbs_a_dat_i[17]
  PIN wbs_a_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 92.520 60.000 93.120 ;
    END
  END wbs_a_dat_i[18]
  PIN wbs_a_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 95.240 60.000 95.840 ;
    END
  END wbs_a_dat_i[19]
  PIN wbs_a_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 52.400 60.000 53.000 ;
    END
  END wbs_a_dat_i[1]
  PIN wbs_a_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 97.280 60.000 97.880 ;
    END
  END wbs_a_dat_i[20]
  PIN wbs_a_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 100.000 60.000 100.600 ;
    END
  END wbs_a_dat_i[21]
  PIN wbs_a_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 102.040 60.000 102.640 ;
    END
  END wbs_a_dat_i[22]
  PIN wbs_a_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 104.760 60.000 105.360 ;
    END
  END wbs_a_dat_i[23]
  PIN wbs_a_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 106.800 60.000 107.400 ;
    END
  END wbs_a_dat_i[24]
  PIN wbs_a_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 109.520 60.000 110.120 ;
    END
  END wbs_a_dat_i[25]
  PIN wbs_a_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 111.560 60.000 112.160 ;
    END
  END wbs_a_dat_i[26]
  PIN wbs_a_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 114.280 60.000 114.880 ;
    END
  END wbs_a_dat_i[27]
  PIN wbs_a_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 116.320 60.000 116.920 ;
    END
  END wbs_a_dat_i[28]
  PIN wbs_a_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 118.360 60.000 118.960 ;
    END
  END wbs_a_dat_i[29]
  PIN wbs_a_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 55.120 60.000 55.720 ;
    END
  END wbs_a_dat_i[2]
  PIN wbs_a_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 121.080 60.000 121.680 ;
    END
  END wbs_a_dat_i[30]
  PIN wbs_a_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 123.120 60.000 123.720 ;
    END
  END wbs_a_dat_i[31]
  PIN wbs_a_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 57.160 60.000 57.760 ;
    END
  END wbs_a_dat_i[3]
  PIN wbs_a_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 59.200 60.000 59.800 ;
    END
  END wbs_a_dat_i[4]
  PIN wbs_a_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 61.920 60.000 62.520 ;
    END
  END wbs_a_dat_i[5]
  PIN wbs_a_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 63.960 60.000 64.560 ;
    END
  END wbs_a_dat_i[6]
  PIN wbs_a_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 66.680 60.000 67.280 ;
    END
  END wbs_a_dat_i[7]
  PIN wbs_a_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 68.720 60.000 69.320 ;
    END
  END wbs_a_dat_i[8]
  PIN wbs_a_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 71.440 60.000 72.040 ;
    END
  END wbs_a_dat_i[9]
  PIN wbs_a_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 125.840 60.000 126.440 ;
    END
  END wbs_a_dat_o[0]
  PIN wbs_a_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 149.640 60.000 150.240 ;
    END
  END wbs_a_dat_o[10]
  PIN wbs_a_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 151.680 60.000 152.280 ;
    END
  END wbs_a_dat_o[11]
  PIN wbs_a_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 154.400 60.000 155.000 ;
    END
  END wbs_a_dat_o[12]
  PIN wbs_a_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 156.440 60.000 157.040 ;
    END
  END wbs_a_dat_o[13]
  PIN wbs_a_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 159.160 60.000 159.760 ;
    END
  END wbs_a_dat_o[14]
  PIN wbs_a_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 161.200 60.000 161.800 ;
    END
  END wbs_a_dat_o[15]
  PIN wbs_a_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 163.920 60.000 164.520 ;
    END
  END wbs_a_dat_o[16]
  PIN wbs_a_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 165.960 60.000 166.560 ;
    END
  END wbs_a_dat_o[17]
  PIN wbs_a_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 168.680 60.000 169.280 ;
    END
  END wbs_a_dat_o[18]
  PIN wbs_a_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 170.720 60.000 171.320 ;
    END
  END wbs_a_dat_o[19]
  PIN wbs_a_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 127.880 60.000 128.480 ;
    END
  END wbs_a_dat_o[1]
  PIN wbs_a_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 172.760 60.000 173.360 ;
    END
  END wbs_a_dat_o[20]
  PIN wbs_a_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 175.480 60.000 176.080 ;
    END
  END wbs_a_dat_o[21]
  PIN wbs_a_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 177.520 60.000 178.120 ;
    END
  END wbs_a_dat_o[22]
  PIN wbs_a_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 180.240 60.000 180.840 ;
    END
  END wbs_a_dat_o[23]
  PIN wbs_a_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 182.280 60.000 182.880 ;
    END
  END wbs_a_dat_o[24]
  PIN wbs_a_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 185.000 60.000 185.600 ;
    END
  END wbs_a_dat_o[25]
  PIN wbs_a_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 187.040 60.000 187.640 ;
    END
  END wbs_a_dat_o[26]
  PIN wbs_a_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 189.760 60.000 190.360 ;
    END
  END wbs_a_dat_o[27]
  PIN wbs_a_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 191.800 60.000 192.400 ;
    END
  END wbs_a_dat_o[28]
  PIN wbs_a_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 194.520 60.000 195.120 ;
    END
  END wbs_a_dat_o[29]
  PIN wbs_a_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 130.600 60.000 131.200 ;
    END
  END wbs_a_dat_o[2]
  PIN wbs_a_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 196.560 60.000 197.160 ;
    END
  END wbs_a_dat_o[30]
  PIN wbs_a_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 199.280 60.000 199.880 ;
    END
  END wbs_a_dat_o[31]
  PIN wbs_a_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 132.640 60.000 133.240 ;
    END
  END wbs_a_dat_o[3]
  PIN wbs_a_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 135.360 60.000 135.960 ;
    END
  END wbs_a_dat_o[4]
  PIN wbs_a_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 137.400 60.000 138.000 ;
    END
  END wbs_a_dat_o[5]
  PIN wbs_a_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 140.120 60.000 140.720 ;
    END
  END wbs_a_dat_o[6]
  PIN wbs_a_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 142.160 60.000 142.760 ;
    END
  END wbs_a_dat_o[7]
  PIN wbs_a_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 144.880 60.000 145.480 ;
    END
  END wbs_a_dat_o[8]
  PIN wbs_a_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 146.920 60.000 147.520 ;
    END
  END wbs_a_dat_o[9]
  PIN wbs_a_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 17.040 60.000 17.640 ;
    END
  END wbs_a_sel_i[0]
  PIN wbs_a_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 19.080 60.000 19.680 ;
    END
  END wbs_a_sel_i[1]
  PIN wbs_a_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 21.800 60.000 22.400 ;
    END
  END wbs_a_sel_i[2]
  PIN wbs_a_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 23.840 60.000 24.440 ;
    END
  END wbs_a_sel_i[3]
  PIN wbs_a_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 7.520 60.000 8.120 ;
    END
  END wbs_a_stb_i
  PIN wbs_a_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 12.280 60.000 12.880 ;
    END
  END wbs_a_we_i
  PIN wbs_b_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 213.560 60.000 214.160 ;
    END
  END wbs_b_ack_o
  PIN wbs_b_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 225.120 60.000 225.720 ;
    END
  END wbs_b_adr_i[0]
  PIN wbs_b_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 227.840 60.000 228.440 ;
    END
  END wbs_b_adr_i[1]
  PIN wbs_b_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 229.880 60.000 230.480 ;
    END
  END wbs_b_adr_i[2]
  PIN wbs_b_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 231.920 60.000 232.520 ;
    END
  END wbs_b_adr_i[3]
  PIN wbs_b_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 234.640 60.000 235.240 ;
    END
  END wbs_b_adr_i[4]
  PIN wbs_b_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 236.680 60.000 237.280 ;
    END
  END wbs_b_adr_i[5]
  PIN wbs_b_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 239.400 60.000 240.000 ;
    END
  END wbs_b_adr_i[6]
  PIN wbs_b_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 241.440 60.000 242.040 ;
    END
  END wbs_b_adr_i[7]
  PIN wbs_b_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 244.160 60.000 244.760 ;
    END
  END wbs_b_adr_i[8]
  PIN wbs_b_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 246.200 60.000 246.800 ;
    END
  END wbs_b_adr_i[9]
  PIN wbs_b_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 208.800 60.000 209.400 ;
    END
  END wbs_b_cyc_i
  PIN wbs_b_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 248.920 60.000 249.520 ;
    END
  END wbs_b_dat_i[0]
  PIN wbs_b_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 272.720 60.000 273.320 ;
    END
  END wbs_b_dat_i[10]
  PIN wbs_b_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 274.760 60.000 275.360 ;
    END
  END wbs_b_dat_i[11]
  PIN wbs_b_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 277.480 60.000 278.080 ;
    END
  END wbs_b_dat_i[12]
  PIN wbs_b_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 279.520 60.000 280.120 ;
    END
  END wbs_b_dat_i[13]
  PIN wbs_b_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 282.240 60.000 282.840 ;
    END
  END wbs_b_dat_i[14]
  PIN wbs_b_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 284.280 60.000 284.880 ;
    END
  END wbs_b_dat_i[15]
  PIN wbs_b_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 286.320 60.000 286.920 ;
    END
  END wbs_b_dat_i[16]
  PIN wbs_b_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 289.040 60.000 289.640 ;
    END
  END wbs_b_dat_i[17]
  PIN wbs_b_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 291.080 60.000 291.680 ;
    END
  END wbs_b_dat_i[18]
  PIN wbs_b_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 293.800 60.000 294.400 ;
    END
  END wbs_b_dat_i[19]
  PIN wbs_b_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 250.960 60.000 251.560 ;
    END
  END wbs_b_dat_i[1]
  PIN wbs_b_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 295.840 60.000 296.440 ;
    END
  END wbs_b_dat_i[20]
  PIN wbs_b_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 298.560 60.000 299.160 ;
    END
  END wbs_b_dat_i[21]
  PIN wbs_b_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 300.600 60.000 301.200 ;
    END
  END wbs_b_dat_i[22]
  PIN wbs_b_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 303.320 60.000 303.920 ;
    END
  END wbs_b_dat_i[23]
  PIN wbs_b_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 305.360 60.000 305.960 ;
    END
  END wbs_b_dat_i[24]
  PIN wbs_b_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 308.080 60.000 308.680 ;
    END
  END wbs_b_dat_i[25]
  PIN wbs_b_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 310.120 60.000 310.720 ;
    END
  END wbs_b_dat_i[26]
  PIN wbs_b_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 312.840 60.000 313.440 ;
    END
  END wbs_b_dat_i[27]
  PIN wbs_b_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 314.880 60.000 315.480 ;
    END
  END wbs_b_dat_i[28]
  PIN wbs_b_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 317.600 60.000 318.200 ;
    END
  END wbs_b_dat_i[29]
  PIN wbs_b_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 253.680 60.000 254.280 ;
    END
  END wbs_b_dat_i[2]
  PIN wbs_b_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 319.640 60.000 320.240 ;
    END
  END wbs_b_dat_i[30]
  PIN wbs_b_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 322.360 60.000 322.960 ;
    END
  END wbs_b_dat_i[31]
  PIN wbs_b_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 255.720 60.000 256.320 ;
    END
  END wbs_b_dat_i[3]
  PIN wbs_b_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 258.440 60.000 259.040 ;
    END
  END wbs_b_dat_i[4]
  PIN wbs_b_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 260.480 60.000 261.080 ;
    END
  END wbs_b_dat_i[5]
  PIN wbs_b_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 263.200 60.000 263.800 ;
    END
  END wbs_b_dat_i[6]
  PIN wbs_b_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 265.240 60.000 265.840 ;
    END
  END wbs_b_dat_i[7]
  PIN wbs_b_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 267.960 60.000 268.560 ;
    END
  END wbs_b_dat_i[8]
  PIN wbs_b_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 270.000 60.000 270.600 ;
    END
  END wbs_b_dat_i[9]
  PIN wbs_b_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 324.400 60.000 325.000 ;
    END
  END wbs_b_dat_o[0]
  PIN wbs_b_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 348.200 60.000 348.800 ;
    END
  END wbs_b_dat_o[10]
  PIN wbs_b_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 350.240 60.000 350.840 ;
    END
  END wbs_b_dat_o[11]
  PIN wbs_b_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 352.960 60.000 353.560 ;
    END
  END wbs_b_dat_o[12]
  PIN wbs_b_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 355.000 60.000 355.600 ;
    END
  END wbs_b_dat_o[13]
  PIN wbs_b_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 357.720 60.000 358.320 ;
    END
  END wbs_b_dat_o[14]
  PIN wbs_b_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 359.760 60.000 360.360 ;
    END
  END wbs_b_dat_o[15]
  PIN wbs_b_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 362.480 60.000 363.080 ;
    END
  END wbs_b_dat_o[16]
  PIN wbs_b_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 364.520 60.000 365.120 ;
    END
  END wbs_b_dat_o[17]
  PIN wbs_b_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 367.240 60.000 367.840 ;
    END
  END wbs_b_dat_o[18]
  PIN wbs_b_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 369.280 60.000 369.880 ;
    END
  END wbs_b_dat_o[19]
  PIN wbs_b_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 327.120 60.000 327.720 ;
    END
  END wbs_b_dat_o[1]
  PIN wbs_b_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 372.000 60.000 372.600 ;
    END
  END wbs_b_dat_o[20]
  PIN wbs_b_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 374.040 60.000 374.640 ;
    END
  END wbs_b_dat_o[21]
  PIN wbs_b_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 376.760 60.000 377.360 ;
    END
  END wbs_b_dat_o[22]
  PIN wbs_b_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 378.800 60.000 379.400 ;
    END
  END wbs_b_dat_o[23]
  PIN wbs_b_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 381.520 60.000 382.120 ;
    END
  END wbs_b_dat_o[24]
  PIN wbs_b_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 383.560 60.000 384.160 ;
    END
  END wbs_b_dat_o[25]
  PIN wbs_b_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 386.280 60.000 386.880 ;
    END
  END wbs_b_dat_o[26]
  PIN wbs_b_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 388.320 60.000 388.920 ;
    END
  END wbs_b_dat_o[27]
  PIN wbs_b_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 391.040 60.000 391.640 ;
    END
  END wbs_b_dat_o[28]
  PIN wbs_b_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 393.080 60.000 393.680 ;
    END
  END wbs_b_dat_o[29]
  PIN wbs_b_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 329.160 60.000 329.760 ;
    END
  END wbs_b_dat_o[2]
  PIN wbs_b_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 395.800 60.000 396.400 ;
    END
  END wbs_b_dat_o[30]
  PIN wbs_b_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 397.840 60.000 398.440 ;
    END
  END wbs_b_dat_o[31]
  PIN wbs_b_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 331.880 60.000 332.480 ;
    END
  END wbs_b_dat_o[3]
  PIN wbs_b_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 333.920 60.000 334.520 ;
    END
  END wbs_b_dat_o[4]
  PIN wbs_b_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 336.640 60.000 337.240 ;
    END
  END wbs_b_dat_o[5]
  PIN wbs_b_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 338.680 60.000 339.280 ;
    END
  END wbs_b_dat_o[6]
  PIN wbs_b_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 341.400 60.000 342.000 ;
    END
  END wbs_b_dat_o[7]
  PIN wbs_b_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 343.440 60.000 344.040 ;
    END
  END wbs_b_dat_o[8]
  PIN wbs_b_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 345.480 60.000 346.080 ;
    END
  END wbs_b_dat_o[9]
  PIN wbs_b_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 215.600 60.000 216.200 ;
    END
  END wbs_b_sel_i[0]
  PIN wbs_b_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 218.320 60.000 218.920 ;
    END
  END wbs_b_sel_i[1]
  PIN wbs_b_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 220.360 60.000 220.960 ;
    END
  END wbs_b_sel_i[2]
  PIN wbs_b_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 223.080 60.000 223.680 ;
    END
  END wbs_b_sel_i[3]
  PIN wbs_b_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 206.080 60.000 206.680 ;
    END
  END wbs_b_stb_i
  PIN wbs_b_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 210.840 60.000 211.440 ;
    END
  END wbs_b_we_i
  PIN writable_port_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 0.720 60.000 1.320 ;
    END
  END writable_port_req
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 59.655 389.045 ;
      LAYER met1 ;
        RECT 1.910 10.640 59.925 389.200 ;
      LAYER met2 ;
        RECT 1.940 0.835 59.710 398.325 ;
      LAYER met3 ;
        RECT 4.400 397.440 55.600 398.305 ;
        RECT 3.990 396.800 59.735 397.440 ;
        RECT 3.990 395.440 55.600 396.800 ;
        RECT 4.400 395.400 55.600 395.440 ;
        RECT 4.400 394.080 59.735 395.400 ;
        RECT 4.400 394.040 55.600 394.080 ;
        RECT 3.990 392.680 55.600 394.040 ;
        RECT 3.990 392.040 59.735 392.680 ;
        RECT 4.400 390.640 55.600 392.040 ;
        RECT 3.990 389.320 59.735 390.640 ;
        RECT 3.990 388.640 55.600 389.320 ;
        RECT 4.400 387.920 55.600 388.640 ;
        RECT 4.400 387.280 59.735 387.920 ;
        RECT 4.400 387.240 55.600 387.280 ;
        RECT 3.990 385.880 55.600 387.240 ;
        RECT 3.990 385.240 59.735 385.880 ;
        RECT 4.400 384.560 59.735 385.240 ;
        RECT 4.400 383.840 55.600 384.560 ;
        RECT 3.990 383.160 55.600 383.840 ;
        RECT 3.990 382.520 59.735 383.160 ;
        RECT 3.990 381.840 55.600 382.520 ;
        RECT 4.400 381.120 55.600 381.840 ;
        RECT 4.400 380.440 59.735 381.120 ;
        RECT 3.990 379.800 59.735 380.440 ;
        RECT 3.990 378.440 55.600 379.800 ;
        RECT 4.400 378.400 55.600 378.440 ;
        RECT 4.400 377.760 59.735 378.400 ;
        RECT 4.400 377.040 55.600 377.760 ;
        RECT 3.990 376.360 55.600 377.040 ;
        RECT 3.990 375.720 59.735 376.360 ;
        RECT 4.400 375.040 59.735 375.720 ;
        RECT 4.400 374.320 55.600 375.040 ;
        RECT 3.990 373.640 55.600 374.320 ;
        RECT 3.990 373.000 59.735 373.640 ;
        RECT 3.990 372.320 55.600 373.000 ;
        RECT 4.400 371.600 55.600 372.320 ;
        RECT 4.400 370.920 59.735 371.600 ;
        RECT 3.990 370.280 59.735 370.920 ;
        RECT 3.990 368.920 55.600 370.280 ;
        RECT 4.400 368.880 55.600 368.920 ;
        RECT 4.400 368.240 59.735 368.880 ;
        RECT 4.400 367.520 55.600 368.240 ;
        RECT 3.990 366.840 55.600 367.520 ;
        RECT 3.990 365.520 59.735 366.840 ;
        RECT 4.400 364.120 55.600 365.520 ;
        RECT 3.990 363.480 59.735 364.120 ;
        RECT 3.990 362.120 55.600 363.480 ;
        RECT 4.400 362.080 55.600 362.120 ;
        RECT 4.400 360.760 59.735 362.080 ;
        RECT 4.400 360.720 55.600 360.760 ;
        RECT 3.990 359.360 55.600 360.720 ;
        RECT 3.990 358.720 59.735 359.360 ;
        RECT 4.400 357.320 55.600 358.720 ;
        RECT 3.990 356.000 59.735 357.320 ;
        RECT 3.990 355.320 55.600 356.000 ;
        RECT 4.400 354.600 55.600 355.320 ;
        RECT 4.400 353.960 59.735 354.600 ;
        RECT 4.400 353.920 55.600 353.960 ;
        RECT 3.990 352.600 55.600 353.920 ;
        RECT 4.400 352.560 55.600 352.600 ;
        RECT 4.400 351.240 59.735 352.560 ;
        RECT 4.400 351.200 55.600 351.240 ;
        RECT 3.990 349.840 55.600 351.200 ;
        RECT 3.990 349.200 59.735 349.840 ;
        RECT 4.400 347.800 55.600 349.200 ;
        RECT 3.990 346.480 59.735 347.800 ;
        RECT 3.990 345.800 55.600 346.480 ;
        RECT 4.400 345.080 55.600 345.800 ;
        RECT 4.400 344.440 59.735 345.080 ;
        RECT 4.400 344.400 55.600 344.440 ;
        RECT 3.990 343.040 55.600 344.400 ;
        RECT 3.990 342.400 59.735 343.040 ;
        RECT 4.400 341.000 55.600 342.400 ;
        RECT 3.990 339.680 59.735 341.000 ;
        RECT 3.990 339.000 55.600 339.680 ;
        RECT 4.400 338.280 55.600 339.000 ;
        RECT 4.400 337.640 59.735 338.280 ;
        RECT 4.400 337.600 55.600 337.640 ;
        RECT 3.990 336.240 55.600 337.600 ;
        RECT 3.990 335.600 59.735 336.240 ;
        RECT 4.400 334.920 59.735 335.600 ;
        RECT 4.400 334.200 55.600 334.920 ;
        RECT 3.990 333.520 55.600 334.200 ;
        RECT 3.990 332.880 59.735 333.520 ;
        RECT 3.990 332.200 55.600 332.880 ;
        RECT 4.400 331.480 55.600 332.200 ;
        RECT 4.400 330.800 59.735 331.480 ;
        RECT 3.990 330.160 59.735 330.800 ;
        RECT 3.990 329.480 55.600 330.160 ;
        RECT 4.400 328.760 55.600 329.480 ;
        RECT 4.400 328.120 59.735 328.760 ;
        RECT 4.400 328.080 55.600 328.120 ;
        RECT 3.990 326.720 55.600 328.080 ;
        RECT 3.990 326.080 59.735 326.720 ;
        RECT 4.400 325.400 59.735 326.080 ;
        RECT 4.400 324.680 55.600 325.400 ;
        RECT 3.990 324.000 55.600 324.680 ;
        RECT 3.990 323.360 59.735 324.000 ;
        RECT 3.990 322.680 55.600 323.360 ;
        RECT 4.400 321.960 55.600 322.680 ;
        RECT 4.400 321.280 59.735 321.960 ;
        RECT 3.990 320.640 59.735 321.280 ;
        RECT 3.990 319.280 55.600 320.640 ;
        RECT 4.400 319.240 55.600 319.280 ;
        RECT 4.400 318.600 59.735 319.240 ;
        RECT 4.400 317.880 55.600 318.600 ;
        RECT 3.990 317.200 55.600 317.880 ;
        RECT 3.990 315.880 59.735 317.200 ;
        RECT 4.400 314.480 55.600 315.880 ;
        RECT 3.990 313.840 59.735 314.480 ;
        RECT 3.990 312.480 55.600 313.840 ;
        RECT 4.400 312.440 55.600 312.480 ;
        RECT 4.400 311.120 59.735 312.440 ;
        RECT 4.400 311.080 55.600 311.120 ;
        RECT 3.990 309.720 55.600 311.080 ;
        RECT 3.990 309.080 59.735 309.720 ;
        RECT 4.400 307.680 55.600 309.080 ;
        RECT 3.990 306.360 59.735 307.680 ;
        RECT 4.400 304.960 55.600 306.360 ;
        RECT 3.990 304.320 59.735 304.960 ;
        RECT 3.990 302.960 55.600 304.320 ;
        RECT 4.400 302.920 55.600 302.960 ;
        RECT 4.400 301.600 59.735 302.920 ;
        RECT 4.400 301.560 55.600 301.600 ;
        RECT 3.990 300.200 55.600 301.560 ;
        RECT 3.990 299.560 59.735 300.200 ;
        RECT 4.400 298.160 55.600 299.560 ;
        RECT 3.990 296.840 59.735 298.160 ;
        RECT 3.990 296.160 55.600 296.840 ;
        RECT 4.400 295.440 55.600 296.160 ;
        RECT 4.400 294.800 59.735 295.440 ;
        RECT 4.400 294.760 55.600 294.800 ;
        RECT 3.990 293.400 55.600 294.760 ;
        RECT 3.990 292.760 59.735 293.400 ;
        RECT 4.400 292.080 59.735 292.760 ;
        RECT 4.400 291.360 55.600 292.080 ;
        RECT 3.990 290.680 55.600 291.360 ;
        RECT 3.990 290.040 59.735 290.680 ;
        RECT 3.990 289.360 55.600 290.040 ;
        RECT 4.400 288.640 55.600 289.360 ;
        RECT 4.400 287.960 59.735 288.640 ;
        RECT 3.990 287.320 59.735 287.960 ;
        RECT 3.990 285.960 55.600 287.320 ;
        RECT 4.400 285.920 55.600 285.960 ;
        RECT 4.400 285.280 59.735 285.920 ;
        RECT 4.400 284.560 55.600 285.280 ;
        RECT 3.990 283.880 55.600 284.560 ;
        RECT 3.990 283.240 59.735 283.880 ;
        RECT 4.400 281.840 55.600 283.240 ;
        RECT 3.990 280.520 59.735 281.840 ;
        RECT 3.990 279.840 55.600 280.520 ;
        RECT 4.400 279.120 55.600 279.840 ;
        RECT 4.400 278.480 59.735 279.120 ;
        RECT 4.400 278.440 55.600 278.480 ;
        RECT 3.990 277.080 55.600 278.440 ;
        RECT 3.990 276.440 59.735 277.080 ;
        RECT 4.400 275.760 59.735 276.440 ;
        RECT 4.400 275.040 55.600 275.760 ;
        RECT 3.990 274.360 55.600 275.040 ;
        RECT 3.990 273.720 59.735 274.360 ;
        RECT 3.990 273.040 55.600 273.720 ;
        RECT 4.400 272.320 55.600 273.040 ;
        RECT 4.400 271.640 59.735 272.320 ;
        RECT 3.990 271.000 59.735 271.640 ;
        RECT 3.990 269.640 55.600 271.000 ;
        RECT 4.400 269.600 55.600 269.640 ;
        RECT 4.400 268.960 59.735 269.600 ;
        RECT 4.400 268.240 55.600 268.960 ;
        RECT 3.990 267.560 55.600 268.240 ;
        RECT 3.990 266.240 59.735 267.560 ;
        RECT 4.400 264.840 55.600 266.240 ;
        RECT 3.990 264.200 59.735 264.840 ;
        RECT 3.990 262.840 55.600 264.200 ;
        RECT 4.400 262.800 55.600 262.840 ;
        RECT 4.400 261.480 59.735 262.800 ;
        RECT 4.400 261.440 55.600 261.480 ;
        RECT 3.990 260.120 55.600 261.440 ;
        RECT 4.400 260.080 55.600 260.120 ;
        RECT 4.400 259.440 59.735 260.080 ;
        RECT 4.400 258.720 55.600 259.440 ;
        RECT 3.990 258.040 55.600 258.720 ;
        RECT 3.990 256.720 59.735 258.040 ;
        RECT 4.400 255.320 55.600 256.720 ;
        RECT 3.990 254.680 59.735 255.320 ;
        RECT 3.990 253.320 55.600 254.680 ;
        RECT 4.400 253.280 55.600 253.320 ;
        RECT 4.400 251.960 59.735 253.280 ;
        RECT 4.400 251.920 55.600 251.960 ;
        RECT 3.990 250.560 55.600 251.920 ;
        RECT 3.990 249.920 59.735 250.560 ;
        RECT 4.400 248.520 55.600 249.920 ;
        RECT 3.990 247.200 59.735 248.520 ;
        RECT 3.990 246.520 55.600 247.200 ;
        RECT 4.400 245.800 55.600 246.520 ;
        RECT 4.400 245.160 59.735 245.800 ;
        RECT 4.400 245.120 55.600 245.160 ;
        RECT 3.990 243.760 55.600 245.120 ;
        RECT 3.990 243.120 59.735 243.760 ;
        RECT 4.400 242.440 59.735 243.120 ;
        RECT 4.400 241.720 55.600 242.440 ;
        RECT 3.990 241.040 55.600 241.720 ;
        RECT 3.990 240.400 59.735 241.040 ;
        RECT 3.990 239.720 55.600 240.400 ;
        RECT 4.400 239.000 55.600 239.720 ;
        RECT 4.400 238.320 59.735 239.000 ;
        RECT 3.990 237.680 59.735 238.320 ;
        RECT 3.990 237.000 55.600 237.680 ;
        RECT 4.400 236.280 55.600 237.000 ;
        RECT 4.400 235.640 59.735 236.280 ;
        RECT 4.400 235.600 55.600 235.640 ;
        RECT 3.990 234.240 55.600 235.600 ;
        RECT 3.990 233.600 59.735 234.240 ;
        RECT 4.400 232.920 59.735 233.600 ;
        RECT 4.400 232.200 55.600 232.920 ;
        RECT 3.990 231.520 55.600 232.200 ;
        RECT 3.990 230.880 59.735 231.520 ;
        RECT 3.990 230.200 55.600 230.880 ;
        RECT 4.400 229.480 55.600 230.200 ;
        RECT 4.400 228.840 59.735 229.480 ;
        RECT 4.400 228.800 55.600 228.840 ;
        RECT 3.990 227.440 55.600 228.800 ;
        RECT 3.990 226.800 59.735 227.440 ;
        RECT 4.400 226.120 59.735 226.800 ;
        RECT 4.400 225.400 55.600 226.120 ;
        RECT 3.990 224.720 55.600 225.400 ;
        RECT 3.990 224.080 59.735 224.720 ;
        RECT 3.990 223.400 55.600 224.080 ;
        RECT 4.400 222.680 55.600 223.400 ;
        RECT 4.400 222.000 59.735 222.680 ;
        RECT 3.990 221.360 59.735 222.000 ;
        RECT 3.990 220.000 55.600 221.360 ;
        RECT 4.400 219.960 55.600 220.000 ;
        RECT 4.400 219.320 59.735 219.960 ;
        RECT 4.400 218.600 55.600 219.320 ;
        RECT 3.990 217.920 55.600 218.600 ;
        RECT 3.990 216.600 59.735 217.920 ;
        RECT 4.400 215.200 55.600 216.600 ;
        RECT 3.990 214.560 59.735 215.200 ;
        RECT 3.990 213.880 55.600 214.560 ;
        RECT 4.400 213.160 55.600 213.880 ;
        RECT 4.400 212.480 59.735 213.160 ;
        RECT 3.990 211.840 59.735 212.480 ;
        RECT 3.990 210.480 55.600 211.840 ;
        RECT 4.400 210.440 55.600 210.480 ;
        RECT 4.400 209.800 59.735 210.440 ;
        RECT 4.400 209.080 55.600 209.800 ;
        RECT 3.990 208.400 55.600 209.080 ;
        RECT 3.990 207.080 59.735 208.400 ;
        RECT 4.400 205.680 55.600 207.080 ;
        RECT 3.990 205.040 59.735 205.680 ;
        RECT 3.990 203.680 55.600 205.040 ;
        RECT 4.400 203.640 55.600 203.680 ;
        RECT 4.400 202.320 59.735 203.640 ;
        RECT 4.400 202.280 55.600 202.320 ;
        RECT 3.990 200.920 55.600 202.280 ;
        RECT 3.990 200.280 59.735 200.920 ;
        RECT 4.400 198.880 55.600 200.280 ;
        RECT 3.990 197.560 59.735 198.880 ;
        RECT 3.990 196.880 55.600 197.560 ;
        RECT 4.400 196.160 55.600 196.880 ;
        RECT 4.400 195.520 59.735 196.160 ;
        RECT 4.400 195.480 55.600 195.520 ;
        RECT 3.990 194.120 55.600 195.480 ;
        RECT 3.990 193.480 59.735 194.120 ;
        RECT 4.400 192.800 59.735 193.480 ;
        RECT 4.400 192.080 55.600 192.800 ;
        RECT 3.990 191.400 55.600 192.080 ;
        RECT 3.990 190.760 59.735 191.400 ;
        RECT 3.990 190.080 55.600 190.760 ;
        RECT 4.400 189.360 55.600 190.080 ;
        RECT 4.400 188.680 59.735 189.360 ;
        RECT 3.990 188.040 59.735 188.680 ;
        RECT 3.990 187.360 55.600 188.040 ;
        RECT 4.400 186.640 55.600 187.360 ;
        RECT 4.400 186.000 59.735 186.640 ;
        RECT 4.400 185.960 55.600 186.000 ;
        RECT 3.990 184.600 55.600 185.960 ;
        RECT 3.990 183.960 59.735 184.600 ;
        RECT 4.400 183.280 59.735 183.960 ;
        RECT 4.400 182.560 55.600 183.280 ;
        RECT 3.990 181.880 55.600 182.560 ;
        RECT 3.990 181.240 59.735 181.880 ;
        RECT 3.990 180.560 55.600 181.240 ;
        RECT 4.400 179.840 55.600 180.560 ;
        RECT 4.400 179.160 59.735 179.840 ;
        RECT 3.990 178.520 59.735 179.160 ;
        RECT 3.990 177.160 55.600 178.520 ;
        RECT 4.400 177.120 55.600 177.160 ;
        RECT 4.400 176.480 59.735 177.120 ;
        RECT 4.400 175.760 55.600 176.480 ;
        RECT 3.990 175.080 55.600 175.760 ;
        RECT 3.990 173.760 59.735 175.080 ;
        RECT 4.400 172.360 55.600 173.760 ;
        RECT 3.990 171.720 59.735 172.360 ;
        RECT 3.990 170.360 55.600 171.720 ;
        RECT 4.400 170.320 55.600 170.360 ;
        RECT 4.400 169.680 59.735 170.320 ;
        RECT 4.400 168.960 55.600 169.680 ;
        RECT 3.990 168.280 55.600 168.960 ;
        RECT 3.990 166.960 59.735 168.280 ;
        RECT 4.400 165.560 55.600 166.960 ;
        RECT 3.990 164.920 59.735 165.560 ;
        RECT 3.990 164.240 55.600 164.920 ;
        RECT 4.400 163.520 55.600 164.240 ;
        RECT 4.400 162.840 59.735 163.520 ;
        RECT 3.990 162.200 59.735 162.840 ;
        RECT 3.990 160.840 55.600 162.200 ;
        RECT 4.400 160.800 55.600 160.840 ;
        RECT 4.400 160.160 59.735 160.800 ;
        RECT 4.400 159.440 55.600 160.160 ;
        RECT 3.990 158.760 55.600 159.440 ;
        RECT 3.990 157.440 59.735 158.760 ;
        RECT 4.400 156.040 55.600 157.440 ;
        RECT 3.990 155.400 59.735 156.040 ;
        RECT 3.990 154.040 55.600 155.400 ;
        RECT 4.400 154.000 55.600 154.040 ;
        RECT 4.400 152.680 59.735 154.000 ;
        RECT 4.400 152.640 55.600 152.680 ;
        RECT 3.990 151.280 55.600 152.640 ;
        RECT 3.990 150.640 59.735 151.280 ;
        RECT 4.400 149.240 55.600 150.640 ;
        RECT 3.990 147.920 59.735 149.240 ;
        RECT 3.990 147.240 55.600 147.920 ;
        RECT 4.400 146.520 55.600 147.240 ;
        RECT 4.400 145.880 59.735 146.520 ;
        RECT 4.400 145.840 55.600 145.880 ;
        RECT 3.990 144.480 55.600 145.840 ;
        RECT 3.990 143.840 59.735 144.480 ;
        RECT 4.400 143.160 59.735 143.840 ;
        RECT 4.400 142.440 55.600 143.160 ;
        RECT 3.990 141.760 55.600 142.440 ;
        RECT 3.990 141.120 59.735 141.760 ;
        RECT 4.400 139.720 55.600 141.120 ;
        RECT 3.990 138.400 59.735 139.720 ;
        RECT 3.990 137.720 55.600 138.400 ;
        RECT 4.400 137.000 55.600 137.720 ;
        RECT 4.400 136.360 59.735 137.000 ;
        RECT 4.400 136.320 55.600 136.360 ;
        RECT 3.990 134.960 55.600 136.320 ;
        RECT 3.990 134.320 59.735 134.960 ;
        RECT 4.400 133.640 59.735 134.320 ;
        RECT 4.400 132.920 55.600 133.640 ;
        RECT 3.990 132.240 55.600 132.920 ;
        RECT 3.990 131.600 59.735 132.240 ;
        RECT 3.990 130.920 55.600 131.600 ;
        RECT 4.400 130.200 55.600 130.920 ;
        RECT 4.400 129.520 59.735 130.200 ;
        RECT 3.990 128.880 59.735 129.520 ;
        RECT 3.990 127.520 55.600 128.880 ;
        RECT 4.400 127.480 55.600 127.520 ;
        RECT 4.400 126.840 59.735 127.480 ;
        RECT 4.400 126.120 55.600 126.840 ;
        RECT 3.990 125.440 55.600 126.120 ;
        RECT 3.990 124.120 59.735 125.440 ;
        RECT 4.400 122.720 55.600 124.120 ;
        RECT 3.990 122.080 59.735 122.720 ;
        RECT 3.990 120.720 55.600 122.080 ;
        RECT 4.400 120.680 55.600 120.720 ;
        RECT 4.400 119.360 59.735 120.680 ;
        RECT 4.400 119.320 55.600 119.360 ;
        RECT 3.990 118.000 55.600 119.320 ;
        RECT 4.400 117.960 55.600 118.000 ;
        RECT 4.400 117.320 59.735 117.960 ;
        RECT 4.400 116.600 55.600 117.320 ;
        RECT 3.990 115.920 55.600 116.600 ;
        RECT 3.990 115.280 59.735 115.920 ;
        RECT 3.990 114.600 55.600 115.280 ;
        RECT 4.400 113.880 55.600 114.600 ;
        RECT 4.400 113.200 59.735 113.880 ;
        RECT 3.990 112.560 59.735 113.200 ;
        RECT 3.990 111.200 55.600 112.560 ;
        RECT 4.400 111.160 55.600 111.200 ;
        RECT 4.400 110.520 59.735 111.160 ;
        RECT 4.400 109.800 55.600 110.520 ;
        RECT 3.990 109.120 55.600 109.800 ;
        RECT 3.990 107.800 59.735 109.120 ;
        RECT 4.400 106.400 55.600 107.800 ;
        RECT 3.990 105.760 59.735 106.400 ;
        RECT 3.990 104.400 55.600 105.760 ;
        RECT 4.400 104.360 55.600 104.400 ;
        RECT 4.400 103.040 59.735 104.360 ;
        RECT 4.400 103.000 55.600 103.040 ;
        RECT 3.990 101.640 55.600 103.000 ;
        RECT 3.990 101.000 59.735 101.640 ;
        RECT 4.400 99.600 55.600 101.000 ;
        RECT 3.990 98.280 59.735 99.600 ;
        RECT 3.990 97.600 55.600 98.280 ;
        RECT 4.400 96.880 55.600 97.600 ;
        RECT 4.400 96.240 59.735 96.880 ;
        RECT 4.400 96.200 55.600 96.240 ;
        RECT 3.990 94.880 55.600 96.200 ;
        RECT 4.400 94.840 55.600 94.880 ;
        RECT 4.400 93.520 59.735 94.840 ;
        RECT 4.400 93.480 55.600 93.520 ;
        RECT 3.990 92.120 55.600 93.480 ;
        RECT 3.990 91.480 59.735 92.120 ;
        RECT 4.400 90.080 55.600 91.480 ;
        RECT 3.990 88.760 59.735 90.080 ;
        RECT 3.990 88.080 55.600 88.760 ;
        RECT 4.400 87.360 55.600 88.080 ;
        RECT 4.400 86.720 59.735 87.360 ;
        RECT 4.400 86.680 55.600 86.720 ;
        RECT 3.990 85.320 55.600 86.680 ;
        RECT 3.990 84.680 59.735 85.320 ;
        RECT 4.400 84.000 59.735 84.680 ;
        RECT 4.400 83.280 55.600 84.000 ;
        RECT 3.990 82.600 55.600 83.280 ;
        RECT 3.990 81.960 59.735 82.600 ;
        RECT 3.990 81.280 55.600 81.960 ;
        RECT 4.400 80.560 55.600 81.280 ;
        RECT 4.400 79.880 59.735 80.560 ;
        RECT 3.990 79.240 59.735 79.880 ;
        RECT 3.990 77.880 55.600 79.240 ;
        RECT 4.400 77.840 55.600 77.880 ;
        RECT 4.400 77.200 59.735 77.840 ;
        RECT 4.400 76.480 55.600 77.200 ;
        RECT 3.990 75.800 55.600 76.480 ;
        RECT 3.990 74.480 59.735 75.800 ;
        RECT 4.400 73.080 55.600 74.480 ;
        RECT 3.990 72.440 59.735 73.080 ;
        RECT 3.990 71.760 55.600 72.440 ;
        RECT 4.400 71.040 55.600 71.760 ;
        RECT 4.400 70.360 59.735 71.040 ;
        RECT 3.990 69.720 59.735 70.360 ;
        RECT 3.990 68.360 55.600 69.720 ;
        RECT 4.400 68.320 55.600 68.360 ;
        RECT 4.400 67.680 59.735 68.320 ;
        RECT 4.400 66.960 55.600 67.680 ;
        RECT 3.990 66.280 55.600 66.960 ;
        RECT 3.990 64.960 59.735 66.280 ;
        RECT 4.400 63.560 55.600 64.960 ;
        RECT 3.990 62.920 59.735 63.560 ;
        RECT 3.990 61.560 55.600 62.920 ;
        RECT 4.400 61.520 55.600 61.560 ;
        RECT 4.400 60.200 59.735 61.520 ;
        RECT 4.400 60.160 55.600 60.200 ;
        RECT 3.990 58.800 55.600 60.160 ;
        RECT 3.990 58.160 59.735 58.800 ;
        RECT 4.400 56.760 55.600 58.160 ;
        RECT 3.990 56.120 59.735 56.760 ;
        RECT 3.990 54.760 55.600 56.120 ;
        RECT 4.400 54.720 55.600 54.760 ;
        RECT 4.400 53.400 59.735 54.720 ;
        RECT 4.400 53.360 55.600 53.400 ;
        RECT 3.990 52.000 55.600 53.360 ;
        RECT 3.990 51.360 59.735 52.000 ;
        RECT 4.400 49.960 55.600 51.360 ;
        RECT 3.990 48.640 59.735 49.960 ;
        RECT 4.400 47.240 55.600 48.640 ;
        RECT 3.990 46.600 59.735 47.240 ;
        RECT 3.990 45.240 55.600 46.600 ;
        RECT 4.400 45.200 55.600 45.240 ;
        RECT 4.400 43.880 59.735 45.200 ;
        RECT 4.400 43.840 55.600 43.880 ;
        RECT 3.990 42.480 55.600 43.840 ;
        RECT 3.990 41.840 59.735 42.480 ;
        RECT 4.400 40.440 55.600 41.840 ;
        RECT 3.990 39.120 59.735 40.440 ;
        RECT 3.990 38.440 55.600 39.120 ;
        RECT 4.400 37.720 55.600 38.440 ;
        RECT 4.400 37.080 59.735 37.720 ;
        RECT 4.400 37.040 55.600 37.080 ;
        RECT 3.990 35.680 55.600 37.040 ;
        RECT 3.990 35.040 59.735 35.680 ;
        RECT 4.400 34.360 59.735 35.040 ;
        RECT 4.400 33.640 55.600 34.360 ;
        RECT 3.990 32.960 55.600 33.640 ;
        RECT 3.990 32.320 59.735 32.960 ;
        RECT 3.990 31.640 55.600 32.320 ;
        RECT 4.400 30.920 55.600 31.640 ;
        RECT 4.400 30.240 59.735 30.920 ;
        RECT 3.990 29.600 59.735 30.240 ;
        RECT 3.990 28.240 55.600 29.600 ;
        RECT 4.400 28.200 55.600 28.240 ;
        RECT 4.400 27.560 59.735 28.200 ;
        RECT 4.400 26.840 55.600 27.560 ;
        RECT 3.990 26.160 55.600 26.840 ;
        RECT 3.990 25.520 59.735 26.160 ;
        RECT 4.400 24.840 59.735 25.520 ;
        RECT 4.400 24.120 55.600 24.840 ;
        RECT 3.990 23.440 55.600 24.120 ;
        RECT 3.990 22.800 59.735 23.440 ;
        RECT 3.990 22.120 55.600 22.800 ;
        RECT 4.400 21.400 55.600 22.120 ;
        RECT 4.400 20.720 59.735 21.400 ;
        RECT 3.990 20.080 59.735 20.720 ;
        RECT 3.990 18.720 55.600 20.080 ;
        RECT 4.400 18.680 55.600 18.720 ;
        RECT 4.400 18.040 59.735 18.680 ;
        RECT 4.400 17.320 55.600 18.040 ;
        RECT 3.990 16.640 55.600 17.320 ;
        RECT 3.990 15.320 59.735 16.640 ;
        RECT 4.400 13.920 55.600 15.320 ;
        RECT 3.990 13.280 59.735 13.920 ;
        RECT 3.990 11.920 55.600 13.280 ;
        RECT 4.400 11.880 55.600 11.920 ;
        RECT 4.400 10.560 59.735 11.880 ;
        RECT 4.400 10.520 55.600 10.560 ;
        RECT 3.990 9.160 55.600 10.520 ;
        RECT 3.990 8.520 59.735 9.160 ;
        RECT 4.400 7.120 55.600 8.520 ;
        RECT 3.990 5.800 59.735 7.120 ;
        RECT 3.990 5.120 55.600 5.800 ;
        RECT 4.400 4.400 55.600 5.120 ;
        RECT 4.400 3.760 59.735 4.400 ;
        RECT 4.400 3.720 55.600 3.760 ;
        RECT 3.990 2.400 55.600 3.720 ;
        RECT 4.400 2.360 55.600 2.400 ;
        RECT 4.400 1.720 59.735 2.360 ;
        RECT 4.400 1.000 55.600 1.720 ;
        RECT 3.990 0.855 55.600 1.000 ;
      LAYER met4 ;
        RECT 14.875 10.640 20.635 389.200 ;
        RECT 23.035 10.640 28.795 389.200 ;
        RECT 31.195 10.640 36.955 389.200 ;
        RECT 39.355 10.640 45.115 389.200 ;
        RECT 47.515 10.640 58.585 389.200 ;
  END
END wb_openram_wrapper
END LIBRARY

