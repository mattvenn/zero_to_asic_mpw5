VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_frequency_counter
  CLASS BLOCK ;
  FOREIGN wrapped_frequency_counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 250.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.340 4.000 184.540 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.130 0.000 61.690 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.130 246.000 61.690 250.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.340 4.000 201.540 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 217.340 150.000 218.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.330 0.000 93.890 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 246.000 26.270 250.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 227.540 150.000 228.740 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 67.740 150.000 68.940 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.140 4.000 242.340 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 246.000 0.510 250.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 20.140 150.000 21.340 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.340 4.000 65.540 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.340 4.000 116.540 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.540 4.000 75.740 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 115.340 150.000 116.540 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.740 4.000 238.940 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.540 4.000 228.740 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 0.000 148.630 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.850 0.000 145.410 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 94.940 150.000 96.140 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 0.000 132.530 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 246.000 148.630 250.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 0.000 64.910 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 128.940 150.000 130.140 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.540 4.000 177.740 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 0.000 122.870 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.740 4.000 102.940 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 246.000 103.550 250.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.530 246.000 126.090 250.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 176.540 150.000 177.740 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 246.000 129.310 250.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 246.000 64.910 250.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 173.140 150.000 174.340 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 241.140 150.000 242.340 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.140 4.000 123.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.740 4.000 85.940 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 183.340 150.000 184.540 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.340 4.000 235.540 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.210 0.000 106.770 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.740 4.000 68.940 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 162.940 150.000 164.140 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 108.540 150.000 109.740 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 105.140 150.000 106.340 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.740 4.000 17.940 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 246.000 6.950 250.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 60.940 150.000 62.140 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.690 0.000 55.250 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.330 246.000 93.890 250.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.610 246.000 10.170 250.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 6.540 150.000 7.740 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 135.740 150.000 136.940 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.140 4.000 208.340 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.270 0.000 19.830 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 246.000 52.030 250.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.690 246.000 55.250 250.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 40.540 150.000 41.740 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 207.140 150.000 208.340 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 246.000 68.130 250.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 16.740 150.000 17.940 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 179.940 150.000 181.140 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 246.000 116.430 250.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.540 4.000 211.740 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 13.340 150.000 14.540 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.340 4.000 99.540 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 43.940 150.000 45.140 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.940 4.000 249.140 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.140 4.000 89.340 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.940 4.000 45.140 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.140 4.000 72.340 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.770 0.000 100.330 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 50.740 150.000 51.940 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.940 4.000 130.140 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 122.140 150.000 123.340 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.170 246.000 3.730 250.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 0.000 16.610 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 0.000 42.370 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 237.740 150.000 238.940 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 159.540 150.000 160.740 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.940 4.000 11.140 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.340 4.000 31.540 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 9.940 150.000 11.140 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 210.540 150.000 211.740 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.340 4.000 167.540 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 156.140 150.000 157.340 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.190 246.000 135.750 250.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 37.140 150.000 38.340 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.940 4.000 96.140 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.670 246.000 84.230 250.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 246.000 113.210 250.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.540 4.000 160.740 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.530 0.000 126.090 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 142.540 150.000 143.740 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 0.000 109.990 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.770 246.000 100.330 250.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.140 4.000 21.340 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.210 246.000 106.770 250.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 0.000 68.130 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 54.140 150.000 55.340 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.930 0.000 29.490 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.540 4.000 24.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.540 4.000 58.740 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.740 4.000 187.940 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 77.940 150.000 79.140 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 213.940 150.000 215.140 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 203.740 150.000 204.940 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 246.000 13.390 250.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 230.940 150.000 232.140 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.140 4.000 174.340 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 169.740 150.000 170.940 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 246.000 42.370 250.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 246.000 142.190 250.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.940 4.000 79.140 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 0.000 74.570 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.940 4.000 62.140 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 81.340 150.000 82.540 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.890 0.000 87.450 4.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 74.540 150.000 75.740 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.340 4.000 150.540 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.190 0.000 135.750 4.000 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.740 4.000 51.940 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 246.000 16.610 250.000 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 246.000 77.790 250.000 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 246.000 48.810 250.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 23.540 150.000 24.740 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.490 246.000 23.050 250.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 0.000 81.010 4.000 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.940 4.000 147.140 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.850 246.000 145.410 250.000 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 88.140 150.000 89.340 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.140 4.000 4.340 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 0.000 58.470 4.000 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.740 4.000 153.940 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 64.340 150.000 65.540 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.870 0.000 116.430 4.000 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.340 4.000 133.540 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.740 4.000 204.940 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.030 0.000 45.590 4.000 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 0.000 6.950 4.000 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 -0.260 150.000 0.940 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.540 4.000 126.740 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 246.000 119.650 250.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 149.340 150.000 150.540 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.930 246.000 29.490 250.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.540 4.000 92.740 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 246.000 32.710 250.000 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.140 4.000 140.340 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 0.000 32.710 4.000 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 98.340 150.000 99.540 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 0.000 90.670 4.000 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 234.340 150.000 235.540 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.740 4.000 221.940 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 246.000 58.470 250.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.540 4.000 7.740 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 118.740 150.000 119.940 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 196.940 150.000 198.140 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.140 4.000 225.340 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 152.740 150.000 153.940 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.940 4.000 181.140 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 224.140 150.000 225.340 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 246.000 74.570 250.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 0.000 48.810 4.000 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 125.540 150.000 126.740 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 71.140 150.000 72.340 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.540 4.000 194.740 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 26.940 150.000 28.140 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.490 0.000 23.050 4.000 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.670 0.000 84.230 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 101.740 150.000 102.940 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 244.540 150.000 245.740 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.140 4.000 38.340 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 33.740 150.000 34.940 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 0.000 13.390 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 132.340 150.000 133.540 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.170 0.000 3.730 4.000 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 200.340 150.000 201.540 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 246.000 138.970 250.000 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 47.340 150.000 48.540 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 246.000 132.530 250.000 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.940 4.000 113.140 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.740 4.000 119.940 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 0.000 119.650 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 0.000 142.190 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.540 4.000 143.740 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.940 4.000 215.140 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 246.000 39.150 250.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.140 4.000 106.340 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.370 0.000 35.930 4.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.610 0.000 10.170 4.000 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 246.000 81.010 250.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.370 246.000 35.930 250.000 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.550 0.000 97.110 4.000 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 246.000 109.990 250.000 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 91.540 150.000 92.740 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.140 4.000 157.340 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 190.140 150.000 191.340 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 0.000 39.150 4.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 0.000 71.350 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.740 4.000 34.940 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 186.740 150.000 187.940 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 0.000 113.210 4.000 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 246.000 90.670 250.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.890 246.000 87.450 250.000 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.940 4.000 198.140 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.940 4.000 232.140 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 0.000 138.970 4.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.340 4.000 48.540 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.740 4.000 170.940 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.880 10.640 29.480 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.200 10.640 75.800 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.520 10.640 122.120 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.360 10.640 98.960 236.880 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 145.940 150.000 147.140 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 236.725 ;
      LAYER met1 ;
        RECT 0.070 10.640 145.290 236.880 ;
      LAYER met2 ;
        RECT 0.790 245.720 2.890 248.725 ;
        RECT 4.010 245.720 6.110 248.725 ;
        RECT 7.230 245.720 9.330 248.725 ;
        RECT 10.450 245.720 12.550 248.725 ;
        RECT 13.670 245.720 15.770 248.725 ;
        RECT 16.890 245.720 22.210 248.725 ;
        RECT 23.330 245.720 25.430 248.725 ;
        RECT 26.550 245.720 28.650 248.725 ;
        RECT 29.770 245.720 31.870 248.725 ;
        RECT 32.990 245.720 35.090 248.725 ;
        RECT 36.210 245.720 38.310 248.725 ;
        RECT 39.430 245.720 41.530 248.725 ;
        RECT 42.650 245.720 47.970 248.725 ;
        RECT 49.090 245.720 51.190 248.725 ;
        RECT 52.310 245.720 54.410 248.725 ;
        RECT 55.530 245.720 57.630 248.725 ;
        RECT 58.750 245.720 60.850 248.725 ;
        RECT 61.970 245.720 64.070 248.725 ;
        RECT 65.190 245.720 67.290 248.725 ;
        RECT 68.410 245.720 73.730 248.725 ;
        RECT 74.850 245.720 76.950 248.725 ;
        RECT 78.070 245.720 80.170 248.725 ;
        RECT 81.290 245.720 83.390 248.725 ;
        RECT 84.510 245.720 86.610 248.725 ;
        RECT 87.730 245.720 89.830 248.725 ;
        RECT 90.950 245.720 93.050 248.725 ;
        RECT 94.170 245.720 99.490 248.725 ;
        RECT 100.610 245.720 102.710 248.725 ;
        RECT 103.830 245.720 105.930 248.725 ;
        RECT 107.050 245.720 109.150 248.725 ;
        RECT 110.270 245.720 112.370 248.725 ;
        RECT 113.490 245.720 115.590 248.725 ;
        RECT 116.710 245.720 118.810 248.725 ;
        RECT 119.930 245.720 125.250 248.725 ;
        RECT 126.370 245.720 128.470 248.725 ;
        RECT 129.590 245.720 131.690 248.725 ;
        RECT 132.810 245.720 134.910 248.725 ;
        RECT 136.030 245.720 138.130 248.725 ;
        RECT 139.250 245.720 141.350 248.725 ;
        RECT 142.470 245.720 144.570 248.725 ;
        RECT 0.100 4.280 145.270 245.720 ;
        RECT 0.790 4.000 2.890 4.280 ;
        RECT 4.010 4.000 6.110 4.280 ;
        RECT 7.230 4.000 9.330 4.280 ;
        RECT 10.450 4.000 12.550 4.280 ;
        RECT 13.670 4.000 15.770 4.280 ;
        RECT 16.890 4.000 18.990 4.280 ;
        RECT 20.110 4.000 22.210 4.280 ;
        RECT 23.330 4.000 28.650 4.280 ;
        RECT 29.770 4.000 31.870 4.280 ;
        RECT 32.990 4.000 35.090 4.280 ;
        RECT 36.210 4.000 38.310 4.280 ;
        RECT 39.430 4.000 41.530 4.280 ;
        RECT 42.650 4.000 44.750 4.280 ;
        RECT 45.870 4.000 47.970 4.280 ;
        RECT 49.090 4.000 54.410 4.280 ;
        RECT 55.530 4.000 57.630 4.280 ;
        RECT 58.750 4.000 60.850 4.280 ;
        RECT 61.970 4.000 64.070 4.280 ;
        RECT 65.190 4.000 67.290 4.280 ;
        RECT 68.410 4.000 70.510 4.280 ;
        RECT 71.630 4.000 73.730 4.280 ;
        RECT 74.850 4.000 80.170 4.280 ;
        RECT 81.290 4.000 83.390 4.280 ;
        RECT 84.510 4.000 86.610 4.280 ;
        RECT 87.730 4.000 89.830 4.280 ;
        RECT 90.950 4.000 93.050 4.280 ;
        RECT 94.170 4.000 96.270 4.280 ;
        RECT 97.390 4.000 99.490 4.280 ;
        RECT 100.610 4.000 105.930 4.280 ;
        RECT 107.050 4.000 109.150 4.280 ;
        RECT 110.270 4.000 112.370 4.280 ;
        RECT 113.490 4.000 115.590 4.280 ;
        RECT 116.710 4.000 118.810 4.280 ;
        RECT 119.930 4.000 122.030 4.280 ;
        RECT 123.150 4.000 125.250 4.280 ;
        RECT 126.370 4.000 131.690 4.280 ;
        RECT 132.810 4.000 134.910 4.280 ;
        RECT 136.030 4.000 138.130 4.280 ;
        RECT 139.250 4.000 141.350 4.280 ;
        RECT 142.470 4.000 144.570 4.280 ;
      LAYER met3 ;
        RECT 4.400 247.540 146.000 248.705 ;
        RECT 4.000 246.140 146.000 247.540 ;
        RECT 4.000 244.140 145.600 246.140 ;
        RECT 4.000 242.740 146.000 244.140 ;
        RECT 4.400 240.740 145.600 242.740 ;
        RECT 4.000 239.340 146.000 240.740 ;
        RECT 4.400 237.340 145.600 239.340 ;
        RECT 4.000 235.940 146.000 237.340 ;
        RECT 4.400 233.940 145.600 235.940 ;
        RECT 4.000 232.540 146.000 233.940 ;
        RECT 4.400 230.540 145.600 232.540 ;
        RECT 4.000 229.140 146.000 230.540 ;
        RECT 4.400 227.140 145.600 229.140 ;
        RECT 4.000 225.740 146.000 227.140 ;
        RECT 4.400 223.740 145.600 225.740 ;
        RECT 4.000 222.340 146.000 223.740 ;
        RECT 4.400 220.340 146.000 222.340 ;
        RECT 4.000 218.940 146.000 220.340 ;
        RECT 4.000 216.940 145.600 218.940 ;
        RECT 4.000 215.540 146.000 216.940 ;
        RECT 4.400 213.540 145.600 215.540 ;
        RECT 4.000 212.140 146.000 213.540 ;
        RECT 4.400 210.140 145.600 212.140 ;
        RECT 4.000 208.740 146.000 210.140 ;
        RECT 4.400 206.740 145.600 208.740 ;
        RECT 4.000 205.340 146.000 206.740 ;
        RECT 4.400 203.340 145.600 205.340 ;
        RECT 4.000 201.940 146.000 203.340 ;
        RECT 4.400 199.940 145.600 201.940 ;
        RECT 4.000 198.540 146.000 199.940 ;
        RECT 4.400 196.540 145.600 198.540 ;
        RECT 4.000 195.140 146.000 196.540 ;
        RECT 4.400 193.140 146.000 195.140 ;
        RECT 4.000 191.740 146.000 193.140 ;
        RECT 4.000 189.740 145.600 191.740 ;
        RECT 4.000 188.340 146.000 189.740 ;
        RECT 4.400 186.340 145.600 188.340 ;
        RECT 4.000 184.940 146.000 186.340 ;
        RECT 4.400 182.940 145.600 184.940 ;
        RECT 4.000 181.540 146.000 182.940 ;
        RECT 4.400 179.540 145.600 181.540 ;
        RECT 4.000 178.140 146.000 179.540 ;
        RECT 4.400 176.140 145.600 178.140 ;
        RECT 4.000 174.740 146.000 176.140 ;
        RECT 4.400 172.740 145.600 174.740 ;
        RECT 4.000 171.340 146.000 172.740 ;
        RECT 4.400 169.340 145.600 171.340 ;
        RECT 4.000 167.940 146.000 169.340 ;
        RECT 4.400 165.940 146.000 167.940 ;
        RECT 4.000 164.540 146.000 165.940 ;
        RECT 4.000 162.540 145.600 164.540 ;
        RECT 4.000 161.140 146.000 162.540 ;
        RECT 4.400 159.140 145.600 161.140 ;
        RECT 4.000 157.740 146.000 159.140 ;
        RECT 4.400 155.740 145.600 157.740 ;
        RECT 4.000 154.340 146.000 155.740 ;
        RECT 4.400 152.340 145.600 154.340 ;
        RECT 4.000 150.940 146.000 152.340 ;
        RECT 4.400 148.940 145.600 150.940 ;
        RECT 4.000 147.540 146.000 148.940 ;
        RECT 4.400 145.540 145.600 147.540 ;
        RECT 4.000 144.140 146.000 145.540 ;
        RECT 4.400 142.140 145.600 144.140 ;
        RECT 4.000 140.740 146.000 142.140 ;
        RECT 4.400 138.740 146.000 140.740 ;
        RECT 4.000 137.340 146.000 138.740 ;
        RECT 4.000 135.340 145.600 137.340 ;
        RECT 4.000 133.940 146.000 135.340 ;
        RECT 4.400 131.940 145.600 133.940 ;
        RECT 4.000 130.540 146.000 131.940 ;
        RECT 4.400 128.540 145.600 130.540 ;
        RECT 4.000 127.140 146.000 128.540 ;
        RECT 4.400 125.140 145.600 127.140 ;
        RECT 4.000 123.740 146.000 125.140 ;
        RECT 4.400 121.740 145.600 123.740 ;
        RECT 4.000 120.340 146.000 121.740 ;
        RECT 4.400 118.340 145.600 120.340 ;
        RECT 4.000 116.940 146.000 118.340 ;
        RECT 4.400 114.940 145.600 116.940 ;
        RECT 4.000 113.540 146.000 114.940 ;
        RECT 4.400 111.540 146.000 113.540 ;
        RECT 4.000 110.140 146.000 111.540 ;
        RECT 4.000 108.140 145.600 110.140 ;
        RECT 4.000 106.740 146.000 108.140 ;
        RECT 4.400 104.740 145.600 106.740 ;
        RECT 4.000 103.340 146.000 104.740 ;
        RECT 4.400 101.340 145.600 103.340 ;
        RECT 4.000 99.940 146.000 101.340 ;
        RECT 4.400 97.940 145.600 99.940 ;
        RECT 4.000 96.540 146.000 97.940 ;
        RECT 4.400 94.540 145.600 96.540 ;
        RECT 4.000 93.140 146.000 94.540 ;
        RECT 4.400 91.140 145.600 93.140 ;
        RECT 4.000 89.740 146.000 91.140 ;
        RECT 4.400 87.740 145.600 89.740 ;
        RECT 4.000 86.340 146.000 87.740 ;
        RECT 4.400 84.340 146.000 86.340 ;
        RECT 4.000 82.940 146.000 84.340 ;
        RECT 4.000 80.940 145.600 82.940 ;
        RECT 4.000 79.540 146.000 80.940 ;
        RECT 4.400 77.540 145.600 79.540 ;
        RECT 4.000 76.140 146.000 77.540 ;
        RECT 4.400 74.140 145.600 76.140 ;
        RECT 4.000 72.740 146.000 74.140 ;
        RECT 4.400 70.740 145.600 72.740 ;
        RECT 4.000 69.340 146.000 70.740 ;
        RECT 4.400 67.340 145.600 69.340 ;
        RECT 4.000 65.940 146.000 67.340 ;
        RECT 4.400 63.940 145.600 65.940 ;
        RECT 4.000 62.540 146.000 63.940 ;
        RECT 4.400 60.540 145.600 62.540 ;
        RECT 4.000 59.140 146.000 60.540 ;
        RECT 4.400 57.140 146.000 59.140 ;
        RECT 4.000 55.740 146.000 57.140 ;
        RECT 4.000 53.740 145.600 55.740 ;
        RECT 4.000 52.340 146.000 53.740 ;
        RECT 4.400 50.340 145.600 52.340 ;
        RECT 4.000 48.940 146.000 50.340 ;
        RECT 4.400 46.940 145.600 48.940 ;
        RECT 4.000 45.540 146.000 46.940 ;
        RECT 4.400 43.540 145.600 45.540 ;
        RECT 4.000 42.140 146.000 43.540 ;
        RECT 4.400 40.140 145.600 42.140 ;
        RECT 4.000 38.740 146.000 40.140 ;
        RECT 4.400 36.740 145.600 38.740 ;
        RECT 4.000 35.340 146.000 36.740 ;
        RECT 4.400 33.340 145.600 35.340 ;
        RECT 4.000 31.940 146.000 33.340 ;
        RECT 4.400 29.940 146.000 31.940 ;
        RECT 4.000 28.540 146.000 29.940 ;
        RECT 4.000 26.540 145.600 28.540 ;
        RECT 4.000 25.140 146.000 26.540 ;
        RECT 4.400 23.140 145.600 25.140 ;
        RECT 4.000 21.740 146.000 23.140 ;
        RECT 4.400 19.740 145.600 21.740 ;
        RECT 4.000 18.340 146.000 19.740 ;
        RECT 4.400 16.340 145.600 18.340 ;
        RECT 4.000 14.940 146.000 16.340 ;
        RECT 4.400 12.940 145.600 14.940 ;
        RECT 4.000 11.540 146.000 12.940 ;
        RECT 4.400 9.540 145.600 11.540 ;
        RECT 4.000 8.140 146.000 9.540 ;
        RECT 4.400 6.975 145.600 8.140 ;
      LAYER met4 ;
        RECT 93.215 19.895 96.960 221.505 ;
        RECT 99.360 19.895 120.120 221.505 ;
        RECT 122.520 19.895 137.705 221.505 ;
  END
END wrapped_frequency_counter
END LIBRARY

