magic
tech sky130A
magscale 1 2
timestamp 1646921648
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 177942 700340 177948 700392
rect 178000 700380 178006 700392
rect 218974 700380 218980 700392
rect 178000 700352 218980 700380
rect 178000 700340 178006 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 268378 700340 268384 700392
rect 268436 700380 268442 700392
rect 494790 700380 494796 700392
rect 268436 700352 494796 700380
rect 268436 700340 268442 700352
rect 494790 700340 494796 700352
rect 494848 700340 494854 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 54478 700312 54484 700324
rect 24360 700284 54484 700312
rect 24360 700272 24366 700284
rect 54478 700272 54484 700284
rect 54536 700272 54542 700324
rect 137830 700272 137836 700324
rect 137888 700312 137894 700324
rect 178678 700312 178684 700324
rect 137888 700284 178684 700312
rect 137888 700272 137894 700284
rect 178678 700272 178684 700284
rect 178736 700272 178742 700324
rect 184842 700272 184848 700324
rect 184900 700312 184906 700324
rect 429838 700312 429844 700324
rect 184900 700284 429844 700312
rect 184900 700272 184906 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 504358 700272 504364 700324
rect 504416 700312 504422 700324
rect 527174 700312 527180 700324
rect 504416 700284 527180 700312
rect 504416 700272 504422 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 547138 700272 547144 700324
rect 547196 700312 547202 700324
rect 559650 700312 559656 700324
rect 547196 700284 559656 700312
rect 547196 700272 547202 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 240778 699700 240784 699712
rect 235224 699672 240784 699700
rect 235224 699660 235230 699672
rect 240778 699660 240784 699672
rect 240836 699660 240842 699712
rect 258718 699660 258724 699712
rect 258776 699700 258782 699712
rect 267642 699700 267648 699712
rect 258776 699672 267648 699700
rect 258776 699660 258782 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 359458 699660 359464 699712
rect 359516 699700 359522 699712
rect 364978 699700 364984 699712
rect 359516 699672 364984 699700
rect 359516 699660 359522 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 154114 698912 154120 698964
rect 154172 698952 154178 698964
rect 195238 698952 195244 698964
rect 154172 698924 195244 698952
rect 154172 698912 154178 698924
rect 195238 698912 195244 698924
rect 195296 698912 195302 698964
rect 260098 698912 260104 698964
rect 260156 698952 260162 698964
rect 283834 698952 283840 698964
rect 260156 698924 283840 698952
rect 260156 698912 260162 698924
rect 283834 698912 283840 698924
rect 283892 698912 283898 698964
rect 180702 697552 180708 697604
rect 180760 697592 180766 697604
rect 397454 697592 397460 697604
rect 180760 697564 397460 697592
rect 180760 697552 180766 697564
rect 397454 697552 397460 697564
rect 397512 697552 397518 697604
rect 367738 696940 367744 696992
rect 367796 696980 367802 696992
rect 580166 696980 580172 696992
rect 367796 696952 580172 696980
rect 367796 696940 367802 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 264238 696192 264244 696244
rect 264296 696232 264302 696244
rect 462314 696232 462320 696244
rect 264296 696204 462320 696232
rect 264296 696192 264302 696204
rect 462314 696192 462320 696204
rect 462372 696192 462378 696244
rect 237558 694764 237564 694816
rect 237616 694804 237622 694816
rect 477494 694804 477500 694816
rect 237616 694776 477500 694804
rect 237616 694764 237622 694776
rect 477494 694764 477500 694776
rect 477552 694764 477558 694816
rect 215662 693404 215668 693456
rect 215720 693444 215726 693456
rect 347774 693444 347780 693456
rect 215720 693416 347780 693444
rect 215720 693404 215726 693416
rect 347774 693404 347780 693416
rect 347832 693404 347838 693456
rect 411898 683136 411904 683188
rect 411956 683176 411962 683188
rect 580166 683176 580172 683188
rect 411956 683148 580172 683176
rect 411956 683136 411962 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 71038 670732 71044 670744
rect 3568 670704 71044 670732
rect 3568 670692 3574 670704
rect 71038 670692 71044 670704
rect 71096 670692 71102 670744
rect 222838 670692 222844 670744
rect 222896 670732 222902 670744
rect 580166 670732 580172 670744
rect 222896 670704 580172 670732
rect 222896 670692 222902 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 249058 656928 249064 656940
rect 3568 656900 249064 656928
rect 3568 656888 3574 656900
rect 249058 656888 249064 656900
rect 249116 656888 249122 656940
rect 262858 643084 262864 643136
rect 262916 643124 262922 643136
rect 580166 643124 580172 643136
rect 262916 643096 580172 643124
rect 262916 643084 262922 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 6914 632680 6920 632732
rect 6972 632720 6978 632732
rect 188338 632720 188344 632732
rect 6972 632692 188344 632720
rect 6972 632680 6978 632692
rect 188338 632680 188344 632692
rect 188396 632680 188402 632732
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 7558 632108 7564 632120
rect 3568 632080 7564 632108
rect 3568 632068 3574 632080
rect 7558 632068 7564 632080
rect 7616 632068 7622 632120
rect 269758 630640 269764 630692
rect 269816 630680 269822 630692
rect 580166 630680 580172 630692
rect 269816 630652 580172 630680
rect 269816 630640 269822 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 116578 618304 116584 618316
rect 3568 618276 116584 618304
rect 3568 618264 3574 618276
rect 116578 618264 116584 618276
rect 116636 618264 116642 618316
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 97258 605860 97264 605872
rect 3568 605832 97264 605860
rect 3568 605820 3574 605832
rect 97258 605820 97264 605832
rect 97316 605820 97322 605872
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 253198 579680 253204 579692
rect 3384 579652 253204 579680
rect 3384 579640 3390 579652
rect 253198 579640 253204 579652
rect 253256 579640 253262 579692
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 108298 565876 108304 565888
rect 3292 565848 108304 565876
rect 3292 565836 3298 565848
rect 108298 565836 108304 565848
rect 108356 565836 108362 565888
rect 232498 563048 232504 563100
rect 232556 563088 232562 563100
rect 579798 563088 579804 563100
rect 232556 563060 579804 563088
rect 232556 563048 232562 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 14458 553432 14464 553444
rect 3384 553404 14464 553432
rect 3384 553392 3390 553404
rect 14458 553392 14464 553404
rect 14516 553392 14522 553444
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 94498 527184 94504 527196
rect 3016 527156 94504 527184
rect 3016 527144 3022 527156
rect 94498 527144 94504 527156
rect 94556 527144 94562 527196
rect 266998 524424 267004 524476
rect 267056 524464 267062 524476
rect 580166 524464 580172 524476
rect 267056 524436 580172 524464
rect 267056 524424 267062 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 270494 514808 270500 514820
rect 3568 514780 270500 514808
rect 3568 514768 3574 514780
rect 270494 514768 270500 514780
rect 270552 514768 270558 514820
rect 200022 510620 200028 510672
rect 200080 510660 200086 510672
rect 580166 510660 580172 510672
rect 200080 510632 580172 510660
rect 200080 510620 200086 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 251818 501004 251824 501016
rect 3108 500976 251824 501004
rect 3108 500964 3114 500976
rect 251818 500964 251824 500976
rect 251876 500964 251882 501016
rect 428458 484372 428464 484424
rect 428516 484412 428522 484424
rect 580166 484412 580172 484424
rect 428516 484384 580172 484412
rect 428516 484372 428522 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 251910 474756 251916 474768
rect 3108 474728 251916 474756
rect 3108 474716 3114 474728
rect 251910 474716 251916 474728
rect 251968 474716 251974 474768
rect 410518 470568 410524 470620
rect 410576 470608 410582 470620
rect 579982 470608 579988 470620
rect 410576 470580 579988 470608
rect 410576 470568 410582 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 166258 462380 166264 462392
rect 3568 462352 166264 462380
rect 3568 462340 3574 462352
rect 166258 462340 166264 462352
rect 166316 462340 166322 462392
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 11698 448576 11704 448588
rect 3200 448548 11704 448576
rect 3200 448536 3206 448548
rect 11698 448536 11704 448548
rect 11756 448536 11762 448588
rect 425698 430584 425704 430636
rect 425756 430624 425762 430636
rect 580166 430624 580172 430636
rect 425756 430596 580172 430624
rect 425756 430584 425762 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 2774 423512 2780 423564
rect 2832 423552 2838 423564
rect 4798 423552 4804 423564
rect 2832 423524 4804 423552
rect 2832 423512 2838 423524
rect 4798 423512 4804 423524
rect 4856 423512 4862 423564
rect 226978 418140 226984 418192
rect 227036 418180 227042 418192
rect 580166 418180 580172 418192
rect 227036 418152 580172 418180
rect 227036 418140 227042 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 15838 409884 15844 409896
rect 2924 409856 15844 409884
rect 2924 409844 2930 409856
rect 15838 409844 15844 409856
rect 15896 409844 15902 409896
rect 206278 404336 206284 404388
rect 206336 404376 206342 404388
rect 580166 404376 580172 404388
rect 206336 404348 580172 404376
rect 206336 404336 206342 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 407758 378156 407764 378208
rect 407816 378196 407822 378208
rect 580166 378196 580172 378208
rect 407816 378168 580172 378196
rect 407816 378156 407822 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3510 371220 3516 371272
rect 3568 371260 3574 371272
rect 173158 371260 173164 371272
rect 3568 371232 173164 371260
rect 3568 371220 3574 371232
rect 173158 371220 173164 371232
rect 173216 371220 173222 371272
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 213178 357456 213184 357468
rect 3200 357428 213184 357456
rect 3200 357416 3206 357428
rect 213178 357416 213184 357428
rect 213236 357416 213242 357468
rect 204898 351908 204904 351960
rect 204956 351948 204962 351960
rect 580166 351948 580172 351960
rect 204956 351920 580172 351948
rect 204956 351908 204962 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 224218 345080 224224 345092
rect 3384 345052 224224 345080
rect 3384 345040 3390 345052
rect 224218 345040 224224 345052
rect 224276 345040 224282 345092
rect 257430 324300 257436 324352
rect 257488 324340 257494 324352
rect 580166 324340 580172 324352
rect 257488 324312 580172 324340
rect 257488 324300 257494 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 54478 320832 54484 320884
rect 54536 320872 54542 320884
rect 215018 320872 215024 320884
rect 54536 320844 215024 320872
rect 54536 320832 54542 320844
rect 215018 320832 215024 320844
rect 215076 320832 215082 320884
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 162118 318832 162124 318844
rect 3384 318804 162124 318832
rect 3384 318792 3390 318804
rect 162118 318792 162124 318804
rect 162176 318792 162182 318844
rect 88334 318044 88340 318096
rect 88392 318084 88398 318096
rect 234982 318084 234988 318096
rect 88392 318056 234988 318084
rect 88392 318044 88398 318056
rect 234982 318044 234988 318056
rect 235040 318044 235046 318096
rect 71774 316684 71780 316736
rect 71832 316724 71838 316736
rect 245286 316724 245292 316736
rect 71832 316696 245292 316724
rect 71832 316684 71838 316696
rect 245286 316684 245292 316696
rect 245344 316684 245350 316736
rect 198642 315256 198648 315308
rect 198700 315296 198706 315308
rect 331214 315296 331220 315308
rect 198700 315268 331220 315296
rect 198700 315256 198706 315268
rect 331214 315256 331220 315268
rect 331272 315256 331278 315308
rect 201494 312536 201500 312588
rect 201552 312576 201558 312588
rect 249978 312576 249984 312588
rect 201552 312548 249984 312576
rect 201552 312536 201558 312548
rect 249978 312536 249984 312548
rect 250036 312536 250042 312588
rect 254578 311856 254584 311908
rect 254636 311896 254642 311908
rect 580166 311896 580172 311908
rect 254636 311868 580172 311896
rect 254636 311856 254642 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 225322 309748 225328 309800
rect 225380 309788 225386 309800
rect 232498 309788 232504 309800
rect 225380 309760 232504 309788
rect 225380 309748 225386 309760
rect 232498 309748 232504 309760
rect 232556 309748 232562 309800
rect 238846 309748 238852 309800
rect 238904 309788 238910 309800
rect 412634 309788 412640 309800
rect 238904 309760 412640 309788
rect 238904 309748 238910 309760
rect 412634 309748 412640 309760
rect 412692 309748 412698 309800
rect 208578 307028 208584 307080
rect 208636 307068 208642 307080
rect 226978 307068 226984 307080
rect 208636 307040 226984 307068
rect 208636 307028 208642 307040
rect 226978 307028 226984 307040
rect 227036 307028 227042 307080
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 251266 305028 251272 305040
rect 3292 305000 251272 305028
rect 3292 304988 3298 305000
rect 251266 304988 251272 305000
rect 251324 304988 251330 305040
rect 97258 304308 97264 304360
rect 97316 304348 97322 304360
rect 224678 304348 224684 304360
rect 97316 304320 224684 304348
rect 97316 304308 97322 304320
rect 224678 304308 224684 304320
rect 224736 304308 224742 304360
rect 224218 304240 224224 304292
rect 224276 304280 224282 304292
rect 249886 304280 249892 304292
rect 224276 304252 249892 304280
rect 224276 304240 224282 304252
rect 249886 304240 249892 304252
rect 249944 304240 249950 304292
rect 206002 303628 206008 303680
rect 206060 303668 206066 303680
rect 299474 303668 299480 303680
rect 206060 303640 299480 303668
rect 206060 303628 206066 303640
rect 299474 303628 299480 303640
rect 299532 303628 299538 303680
rect 162118 302880 162124 302932
rect 162176 302920 162182 302932
rect 246574 302920 246580 302932
rect 162176 302892 246580 302920
rect 162176 302880 162182 302892
rect 246574 302880 246580 302892
rect 246632 302880 246638 302932
rect 249058 302608 249064 302660
rect 249116 302648 249122 302660
rect 252554 302648 252560 302660
rect 249116 302620 252560 302648
rect 249116 302608 249122 302620
rect 252554 302608 252560 302620
rect 252612 302608 252618 302660
rect 236914 302268 236920 302320
rect 236972 302308 236978 302320
rect 276658 302308 276664 302320
rect 236972 302280 276664 302308
rect 236972 302268 236978 302280
rect 276658 302268 276664 302280
rect 276716 302268 276722 302320
rect 218882 302200 218888 302252
rect 218940 302240 218946 302252
rect 316034 302240 316040 302252
rect 218940 302212 316040 302240
rect 218940 302200 218946 302212
rect 316034 302200 316040 302212
rect 316092 302200 316098 302252
rect 198550 301452 198556 301504
rect 198608 301492 198614 301504
rect 206278 301492 206284 301504
rect 198608 301464 206284 301492
rect 198608 301452 198614 301464
rect 206278 301452 206284 301464
rect 206336 301452 206342 301504
rect 207934 301452 207940 301504
rect 207992 301492 207998 301504
rect 367738 301492 367744 301504
rect 207992 301464 367744 301492
rect 207992 301452 207998 301464
rect 367738 301452 367744 301464
rect 367796 301452 367802 301504
rect 233694 300976 233700 301028
rect 233752 301016 233758 301028
rect 273898 301016 273904 301028
rect 233752 300988 273904 301016
rect 233752 300976 233758 300988
rect 273898 300976 273904 300988
rect 273956 300976 273962 301028
rect 203426 300908 203432 300960
rect 203484 300948 203490 300960
rect 280798 300948 280804 300960
rect 203484 300920 280804 300948
rect 203484 300908 203490 300920
rect 280798 300908 280804 300920
rect 280856 300908 280862 300960
rect 204990 300840 204996 300892
rect 205048 300880 205054 300892
rect 582834 300880 582840 300892
rect 205048 300852 582840 300880
rect 205048 300840 205054 300852
rect 582834 300840 582840 300852
rect 582892 300840 582898 300892
rect 3418 300092 3424 300144
rect 3476 300132 3482 300144
rect 251174 300132 251180 300144
rect 3476 300104 251180 300132
rect 3476 300092 3482 300104
rect 251174 300092 251180 300104
rect 251232 300092 251238 300144
rect 253290 300092 253296 300144
rect 253348 300132 253354 300144
rect 504358 300132 504364 300144
rect 253348 300104 504364 300132
rect 253348 300092 253354 300104
rect 504358 300092 504364 300104
rect 504416 300092 504422 300144
rect 239490 299616 239496 299668
rect 239548 299656 239554 299668
rect 298094 299656 298100 299668
rect 239548 299628 298100 299656
rect 239548 299616 239554 299628
rect 298094 299616 298100 299628
rect 298152 299616 298158 299668
rect 202138 299548 202144 299600
rect 202196 299588 202202 299600
rect 268470 299588 268476 299600
rect 202196 299560 268476 299588
rect 202196 299548 202202 299560
rect 268470 299548 268476 299560
rect 268528 299548 268534 299600
rect 219526 299480 219532 299532
rect 219584 299520 219590 299532
rect 302234 299520 302240 299532
rect 219584 299492 302240 299520
rect 219584 299480 219590 299492
rect 302234 299480 302240 299492
rect 302292 299480 302298 299532
rect 221458 299412 221464 299464
rect 221516 299452 221522 299464
rect 222838 299452 222844 299464
rect 221516 299424 222844 299452
rect 221516 299412 221522 299424
rect 222838 299412 222844 299424
rect 222896 299412 222902 299464
rect 4798 298732 4804 298784
rect 4856 298772 4862 298784
rect 202782 298772 202788 298784
rect 4856 298744 202788 298772
rect 4856 298732 4862 298744
rect 202782 298732 202788 298744
rect 202840 298732 202846 298784
rect 231118 298460 231124 298512
rect 231176 298500 231182 298512
rect 259546 298500 259552 298512
rect 231176 298472 259552 298500
rect 231176 298460 231182 298472
rect 259546 298460 259552 298472
rect 259604 298460 259610 298512
rect 223390 298392 223396 298444
rect 223448 298432 223454 298444
rect 260834 298432 260840 298444
rect 223448 298404 260840 298432
rect 223448 298392 223454 298404
rect 260834 298392 260840 298404
rect 260892 298392 260898 298444
rect 216306 298324 216312 298376
rect 216364 298364 216370 298376
rect 263686 298364 263692 298376
rect 216364 298336 263692 298364
rect 216364 298324 216370 298336
rect 263686 298324 263692 298336
rect 263744 298324 263750 298376
rect 227898 298256 227904 298308
rect 227956 298296 227962 298308
rect 278038 298296 278044 298308
rect 227956 298268 278044 298296
rect 227956 298256 227962 298268
rect 278038 298256 278044 298268
rect 278096 298256 278102 298308
rect 206646 298188 206652 298240
rect 206704 298228 206710 298240
rect 299566 298228 299572 298240
rect 206704 298200 299572 298228
rect 206704 298188 206710 298200
rect 299566 298188 299572 298200
rect 299624 298188 299630 298240
rect 197262 298120 197268 298172
rect 197320 298160 197326 298172
rect 303614 298160 303620 298172
rect 197320 298132 303620 298160
rect 197320 298120 197326 298132
rect 303614 298120 303620 298132
rect 303672 298120 303678 298172
rect 247862 296964 247868 297016
rect 247920 297004 247926 297016
rect 267090 297004 267096 297016
rect 247920 296976 267096 297004
rect 247920 296964 247926 296976
rect 267090 296964 267096 296976
rect 267148 296964 267154 297016
rect 240134 296896 240140 296948
rect 240192 296936 240198 296948
rect 269850 296936 269856 296948
rect 240192 296908 269856 296936
rect 240192 296896 240198 296908
rect 269850 296896 269856 296908
rect 269908 296896 269914 296948
rect 232406 296828 232412 296880
rect 232464 296868 232470 296880
rect 265066 296868 265072 296880
rect 232464 296840 265072 296868
rect 232464 296828 232470 296840
rect 265066 296828 265072 296840
rect 265124 296828 265130 296880
rect 213730 296760 213736 296812
rect 213788 296800 213794 296812
rect 262306 296800 262312 296812
rect 213788 296772 262312 296800
rect 213788 296760 213794 296772
rect 262306 296760 262312 296772
rect 262364 296760 262370 296812
rect 210510 296692 210516 296744
rect 210568 296732 210574 296744
rect 583018 296732 583024 296744
rect 210568 296704 583024 296732
rect 210568 296692 210574 296704
rect 583018 296692 583024 296704
rect 583076 296692 583082 296744
rect 11698 295944 11704 295996
rect 11756 295984 11762 295996
rect 201494 295984 201500 295996
rect 11756 295956 201500 295984
rect 11756 295944 11762 295956
rect 201494 295944 201500 295956
rect 201552 295944 201558 295996
rect 213178 295944 213184 295996
rect 213236 295984 213242 295996
rect 228542 295984 228548 295996
rect 213236 295956 228548 295984
rect 213236 295944 213242 295956
rect 228542 295944 228548 295956
rect 228600 295944 228606 295996
rect 233050 295672 233056 295724
rect 233108 295712 233114 295724
rect 258166 295712 258172 295724
rect 233108 295684 258172 295712
rect 233108 295672 233114 295684
rect 258166 295672 258172 295684
rect 258224 295672 258230 295724
rect 224034 295604 224040 295656
rect 224092 295644 224098 295656
rect 264974 295644 264980 295656
rect 224092 295616 264980 295644
rect 224092 295604 224098 295616
rect 264974 295604 264980 295616
rect 265032 295604 265038 295656
rect 213086 295536 213092 295588
rect 213144 295576 213150 295588
rect 260926 295576 260932 295588
rect 213144 295548 260932 295576
rect 213144 295536 213150 295548
rect 260926 295536 260932 295548
rect 260984 295536 260990 295588
rect 204070 295468 204076 295520
rect 204128 295508 204134 295520
rect 204898 295508 204904 295520
rect 204128 295480 204904 295508
rect 204128 295468 204134 295480
rect 204898 295468 204904 295480
rect 204956 295468 204962 295520
rect 247218 295468 247224 295520
rect 247276 295508 247282 295520
rect 296714 295508 296720 295520
rect 247276 295480 296720 295508
rect 247276 295468 247282 295480
rect 296714 295468 296720 295480
rect 296772 295468 296778 295520
rect 193122 295400 193128 295452
rect 193180 295440 193186 295452
rect 226610 295440 226616 295452
rect 193180 295412 226616 295440
rect 193180 295400 193186 295412
rect 226610 295400 226616 295412
rect 226668 295400 226674 295452
rect 241422 295400 241428 295452
rect 241480 295440 241486 295452
rect 291194 295440 291200 295452
rect 241480 295412 291200 295440
rect 241480 295400 241486 295412
rect 291194 295400 291200 295412
rect 291252 295400 291258 295452
rect 180518 295332 180524 295384
rect 180576 295372 180582 295384
rect 214374 295372 214380 295384
rect 180576 295344 214380 295372
rect 180576 295332 180582 295344
rect 214374 295332 214380 295344
rect 214432 295332 214438 295384
rect 229186 295332 229192 295384
rect 229244 295372 229250 295384
rect 309134 295372 309140 295384
rect 229244 295344 309140 295372
rect 229244 295332 229250 295344
rect 309134 295332 309140 295344
rect 309192 295332 309198 295384
rect 240778 294652 240784 294704
rect 240836 294692 240842 294704
rect 255498 294692 255504 294704
rect 240836 294664 255504 294692
rect 240836 294652 240842 294664
rect 255498 294652 255504 294664
rect 255556 294652 255562 294704
rect 211798 294584 211804 294636
rect 211856 294624 211862 294636
rect 240134 294624 240140 294636
rect 211856 294596 240140 294624
rect 211856 294584 211862 294596
rect 240134 294584 240140 294596
rect 240192 294584 240198 294636
rect 43438 294312 43444 294364
rect 43496 294352 43502 294364
rect 227254 294352 227260 294364
rect 43496 294324 227260 294352
rect 43496 294312 43502 294324
rect 227254 294312 227260 294324
rect 227312 294312 227318 294364
rect 234338 294312 234344 294364
rect 234396 294352 234402 294364
rect 273990 294352 273996 294364
rect 234396 294324 273996 294352
rect 234396 294312 234402 294324
rect 273990 294312 273996 294324
rect 274048 294312 274054 294364
rect 196618 294244 196624 294296
rect 196676 294284 196682 294296
rect 222746 294284 222752 294296
rect 196676 294256 222752 294284
rect 196676 294244 196682 294256
rect 222746 294244 222752 294256
rect 222804 294244 222810 294296
rect 225966 294244 225972 294296
rect 226024 294284 226030 294296
rect 267182 294284 267188 294296
rect 226024 294256 267188 294284
rect 226024 294244 226030 294256
rect 267182 294244 267188 294256
rect 267240 294244 267246 294296
rect 218238 294176 218244 294228
rect 218296 294216 218302 294228
rect 244274 294216 244280 294228
rect 218296 294188 244280 294216
rect 218296 294176 218302 294188
rect 244274 294176 244280 294188
rect 244332 294176 244338 294228
rect 222102 294108 222108 294160
rect 222160 294148 222166 294160
rect 254026 294148 254032 294160
rect 222160 294120 254032 294148
rect 222160 294108 222166 294120
rect 254026 294108 254032 294120
rect 254084 294108 254090 294160
rect 193858 294040 193864 294092
rect 193916 294080 193922 294092
rect 231762 294080 231768 294092
rect 193916 294052 231768 294080
rect 193916 294040 193922 294052
rect 231762 294040 231768 294052
rect 231820 294040 231826 294092
rect 240134 294040 240140 294092
rect 240192 294080 240198 294092
rect 250530 294080 250536 294092
rect 240192 294052 250536 294080
rect 240192 294040 240198 294052
rect 250530 294040 250536 294052
rect 250588 294040 250594 294092
rect 197078 293972 197084 294024
rect 197136 294012 197142 294024
rect 204714 294012 204720 294024
rect 197136 293984 204720 294012
rect 197136 293972 197142 293984
rect 204714 293972 204720 293984
rect 204772 293972 204778 294024
rect 245930 293972 245936 294024
rect 245988 294012 245994 294024
rect 250438 294012 250444 294024
rect 245988 293984 250444 294012
rect 245988 293972 245994 293984
rect 250438 293972 250444 293984
rect 250496 293972 250502 294024
rect 244274 293224 244280 293276
rect 244332 293264 244338 293276
rect 258074 293264 258080 293276
rect 244332 293236 258080 293264
rect 244332 293224 244338 293236
rect 258074 293224 258080 293236
rect 258132 293224 258138 293276
rect 242710 292816 242716 292868
rect 242768 292856 242774 292868
rect 262214 292856 262220 292868
rect 242768 292828 262220 292856
rect 242768 292816 242774 292828
rect 262214 292816 262220 292828
rect 262272 292816 262278 292868
rect 220814 292748 220820 292800
rect 220872 292788 220878 292800
rect 250162 292788 250168 292800
rect 220872 292760 250168 292788
rect 220872 292748 220878 292760
rect 250162 292748 250168 292760
rect 250220 292748 250226 292800
rect 217594 292680 217600 292732
rect 217652 292720 217658 292732
rect 253382 292720 253388 292732
rect 217652 292692 253388 292720
rect 217652 292680 217658 292692
rect 253382 292680 253388 292692
rect 253440 292680 253446 292732
rect 212442 292612 212448 292664
rect 212500 292652 212506 292664
rect 253934 292652 253940 292664
rect 212500 292624 253940 292652
rect 212500 292612 212506 292624
rect 253934 292612 253940 292624
rect 253992 292612 253998 292664
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 21358 292584 21364 292596
rect 3476 292556 21364 292584
rect 3476 292544 3482 292556
rect 21358 292544 21364 292556
rect 21416 292544 21422 292596
rect 195790 292544 195796 292596
rect 195848 292584 195854 292596
rect 205358 292584 205364 292596
rect 195848 292556 205364 292584
rect 195848 292544 195854 292556
rect 205358 292544 205364 292556
rect 205416 292544 205422 292596
rect 207290 292544 207296 292596
rect 207348 292584 207354 292596
rect 271230 292584 271236 292596
rect 207348 292556 271236 292584
rect 207348 292544 207354 292556
rect 271230 292544 271236 292556
rect 271288 292544 271294 292596
rect 201402 292476 201408 292528
rect 201460 292516 201466 292528
rect 204990 292516 204996 292528
rect 201460 292488 204996 292516
rect 201460 292476 201466 292488
rect 204990 292476 204996 292488
rect 205048 292476 205054 292528
rect 210234 292068 210240 292120
rect 210292 292108 210298 292120
rect 210292 292080 219434 292108
rect 210292 292068 210298 292080
rect 11698 291184 11704 291236
rect 11756 291224 11762 291236
rect 197354 291224 197360 291236
rect 11756 291196 197360 291224
rect 11756 291184 11762 291196
rect 197354 291184 197360 291196
rect 197412 291184 197418 291236
rect 219406 291224 219434 292080
rect 241146 292068 241152 292120
rect 241204 292108 241210 292120
rect 241204 292080 248414 292108
rect 241204 292068 241210 292080
rect 248386 291292 248414 292080
rect 253750 291320 253756 291372
rect 253808 291360 253814 291372
rect 259454 291360 259460 291372
rect 253808 291332 259460 291360
rect 253808 291320 253814 291332
rect 259454 291320 259460 291332
rect 259512 291320 259518 291372
rect 255406 291292 255412 291304
rect 248386 291264 255412 291292
rect 255406 291252 255412 291264
rect 255464 291252 255470 291304
rect 256694 291224 256700 291236
rect 219406 291196 256700 291224
rect 256694 291184 256700 291196
rect 256752 291184 256758 291236
rect 253750 291116 253756 291168
rect 253808 291156 253814 291168
rect 407758 291156 407764 291168
rect 253808 291128 407764 291156
rect 253808 291116 253814 291128
rect 407758 291116 407764 291128
rect 407816 291116 407822 291168
rect 188982 289824 188988 289876
rect 189040 289864 189046 289876
rect 197354 289864 197360 289876
rect 189040 289836 197360 289864
rect 189040 289824 189046 289836
rect 197354 289824 197360 289836
rect 197412 289824 197418 289876
rect 195238 289756 195244 289808
rect 195296 289796 195302 289808
rect 197722 289796 197728 289808
rect 195296 289768 197728 289796
rect 195296 289756 195302 289768
rect 197722 289756 197728 289768
rect 197780 289756 197786 289808
rect 253750 288464 253756 288516
rect 253808 288504 253814 288516
rect 272518 288504 272524 288516
rect 253808 288476 272524 288504
rect 253808 288464 253814 288476
rect 272518 288464 272524 288476
rect 272576 288464 272582 288516
rect 186222 288396 186228 288448
rect 186280 288436 186286 288448
rect 197354 288436 197360 288448
rect 186280 288408 197360 288436
rect 186280 288396 186286 288408
rect 197354 288396 197360 288408
rect 197412 288396 197418 288448
rect 252922 288396 252928 288448
rect 252980 288436 252986 288448
rect 296806 288436 296812 288448
rect 252980 288408 296812 288436
rect 252980 288396 252986 288408
rect 296806 288396 296812 288408
rect 296864 288396 296870 288448
rect 190362 287104 190368 287156
rect 190420 287144 190426 287156
rect 197354 287144 197360 287156
rect 190420 287116 197360 287144
rect 190420 287104 190426 287116
rect 197354 287104 197360 287116
rect 197412 287104 197418 287156
rect 182082 287036 182088 287088
rect 182140 287076 182146 287088
rect 197446 287076 197452 287088
rect 182140 287048 197452 287076
rect 182140 287036 182146 287048
rect 197446 287036 197452 287048
rect 197504 287036 197510 287088
rect 253750 287036 253756 287088
rect 253808 287076 253814 287088
rect 305638 287076 305644 287088
rect 253808 287048 305644 287076
rect 253808 287036 253814 287048
rect 305638 287036 305644 287048
rect 305696 287036 305702 287088
rect 71038 286968 71044 287020
rect 71096 287008 71102 287020
rect 197354 287008 197360 287020
rect 71096 286980 197360 287008
rect 71096 286968 71102 286980
rect 197354 286968 197360 286980
rect 197412 286968 197418 287020
rect 253750 285676 253756 285728
rect 253808 285716 253814 285728
rect 381538 285716 381544 285728
rect 253808 285688 381544 285716
rect 253808 285676 253814 285688
rect 381538 285676 381544 285688
rect 381596 285676 381602 285728
rect 253842 285608 253848 285660
rect 253900 285648 253906 285660
rect 410518 285648 410524 285660
rect 253900 285620 410524 285648
rect 253900 285608 253906 285620
rect 410518 285608 410524 285620
rect 410576 285608 410582 285660
rect 3510 284928 3516 284980
rect 3568 284968 3574 284980
rect 196618 284968 196624 284980
rect 3568 284940 196624 284968
rect 3568 284928 3574 284940
rect 196618 284928 196624 284940
rect 196676 284928 196682 284980
rect 188890 284316 188896 284368
rect 188948 284356 188954 284368
rect 197354 284356 197360 284368
rect 188948 284328 197360 284356
rect 188948 284316 188954 284328
rect 197354 284316 197360 284328
rect 197412 284316 197418 284368
rect 253750 282888 253756 282940
rect 253808 282928 253814 282940
rect 278130 282928 278136 282940
rect 253808 282900 278136 282928
rect 253808 282888 253814 282900
rect 278130 282888 278136 282900
rect 278188 282888 278194 282940
rect 250438 282140 250444 282192
rect 250496 282180 250502 282192
rect 580258 282180 580264 282192
rect 250496 282152 580264 282180
rect 250496 282140 250502 282152
rect 580258 282140 580264 282152
rect 580316 282140 580322 282192
rect 252554 280304 252560 280356
rect 252612 280344 252618 280356
rect 255590 280344 255596 280356
rect 252612 280316 255596 280344
rect 252612 280304 252618 280316
rect 255590 280304 255596 280316
rect 255648 280304 255654 280356
rect 183462 280168 183468 280220
rect 183520 280208 183526 280220
rect 197354 280208 197360 280220
rect 183520 280180 197360 280208
rect 183520 280168 183526 280180
rect 197354 280168 197360 280180
rect 197412 280168 197418 280220
rect 253750 280168 253756 280220
rect 253808 280208 253814 280220
rect 295334 280208 295340 280220
rect 253808 280180 295340 280208
rect 253808 280168 253814 280180
rect 295334 280168 295340 280180
rect 295392 280168 295398 280220
rect 35158 278740 35164 278792
rect 35216 278780 35222 278792
rect 197354 278780 197360 278792
rect 35216 278752 197360 278780
rect 35216 278740 35222 278752
rect 197354 278740 197360 278752
rect 197412 278740 197418 278792
rect 253382 277992 253388 278044
rect 253440 278032 253446 278044
rect 263594 278032 263600 278044
rect 253440 278004 263600 278032
rect 253440 277992 253446 278004
rect 263594 277992 263600 278004
rect 263652 277992 263658 278044
rect 190086 277448 190092 277500
rect 190144 277488 190150 277500
rect 197446 277488 197452 277500
rect 190144 277460 197452 277488
rect 190144 277448 190150 277460
rect 197446 277448 197452 277460
rect 197504 277448 197510 277500
rect 187418 277380 187424 277432
rect 187476 277420 187482 277432
rect 197354 277420 197360 277432
rect 187476 277392 197360 277420
rect 187476 277380 187482 277392
rect 197354 277380 197360 277392
rect 197412 277380 197418 277432
rect 253842 277380 253848 277432
rect 253900 277420 253906 277432
rect 283098 277420 283104 277432
rect 253900 277392 283104 277420
rect 253900 277380 253906 277392
rect 283098 277380 283104 277392
rect 283156 277380 283162 277432
rect 251910 276972 251916 277024
rect 251968 277012 251974 277024
rect 252554 277012 252560 277024
rect 251968 276984 252560 277012
rect 251968 276972 251974 276984
rect 252554 276972 252560 276984
rect 252612 276972 252618 277024
rect 195882 276088 195888 276140
rect 195940 276128 195946 276140
rect 197722 276128 197728 276140
rect 195940 276100 197728 276128
rect 195940 276088 195946 276100
rect 197722 276088 197728 276100
rect 197780 276088 197786 276140
rect 190270 276020 190276 276072
rect 190328 276060 190334 276072
rect 197354 276060 197360 276072
rect 190328 276032 197360 276060
rect 190328 276020 190334 276032
rect 197354 276020 197360 276032
rect 197412 276020 197418 276072
rect 253290 276020 253296 276072
rect 253348 276060 253354 276072
rect 566458 276060 566464 276072
rect 253348 276032 566464 276060
rect 253348 276020 253354 276032
rect 566458 276020 566464 276032
rect 566516 276020 566522 276072
rect 187510 274728 187516 274780
rect 187568 274768 187574 274780
rect 197354 274768 197360 274780
rect 187568 274740 197360 274768
rect 187568 274728 187574 274740
rect 197354 274728 197360 274740
rect 197412 274728 197418 274780
rect 184750 274660 184756 274712
rect 184808 274700 184814 274712
rect 197446 274700 197452 274712
rect 184808 274672 197452 274700
rect 184808 274660 184814 274672
rect 197446 274660 197452 274672
rect 197504 274660 197510 274712
rect 253290 274660 253296 274712
rect 253348 274700 253354 274712
rect 385678 274700 385684 274712
rect 253348 274672 385684 274700
rect 253348 274660 253354 274672
rect 385678 274660 385684 274672
rect 385736 274660 385742 274712
rect 116578 274592 116584 274644
rect 116636 274632 116642 274644
rect 197354 274632 197360 274644
rect 116636 274604 197360 274632
rect 116636 274592 116642 274604
rect 197354 274592 197360 274604
rect 197412 274592 197418 274644
rect 252646 274252 252652 274304
rect 252704 274292 252710 274304
rect 254578 274292 254584 274304
rect 252704 274264 254584 274292
rect 252704 274252 252710 274264
rect 254578 274252 254584 274264
rect 254636 274252 254642 274304
rect 253750 273912 253756 273964
rect 253808 273952 253814 273964
rect 283006 273952 283012 273964
rect 253808 273924 283012 273952
rect 253808 273912 253814 273924
rect 283006 273912 283012 273924
rect 283064 273912 283070 273964
rect 253474 272484 253480 272536
rect 253532 272524 253538 272536
rect 287054 272524 287060 272536
rect 253532 272496 287060 272524
rect 253532 272484 253538 272496
rect 287054 272484 287060 272496
rect 287112 272484 287118 272536
rect 252646 272144 252652 272196
rect 252704 272184 252710 272196
rect 254210 272184 254216 272196
rect 252704 272156 254216 272184
rect 252704 272144 252710 272156
rect 254210 272144 254216 272156
rect 254268 272144 254274 272196
rect 251818 271872 251824 271924
rect 251876 271912 251882 271924
rect 252646 271912 252652 271924
rect 251876 271884 252652 271912
rect 251876 271872 251882 271884
rect 252646 271872 252652 271884
rect 252704 271872 252710 271924
rect 574738 271872 574744 271924
rect 574796 271912 574802 271924
rect 580166 271912 580172 271924
rect 574796 271884 580172 271912
rect 574796 271872 574802 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 169754 271804 169760 271856
rect 169812 271844 169818 271856
rect 197354 271844 197360 271856
rect 169812 271816 197360 271844
rect 169812 271804 169818 271816
rect 197354 271804 197360 271816
rect 197412 271804 197418 271856
rect 250530 271124 250536 271176
rect 250588 271164 250594 271176
rect 580350 271164 580356 271176
rect 250588 271136 580356 271164
rect 250588 271124 250594 271136
rect 580350 271124 580356 271136
rect 580408 271124 580414 271176
rect 192846 270512 192852 270564
rect 192904 270552 192910 270564
rect 197446 270552 197452 270564
rect 192904 270524 197452 270552
rect 192904 270512 192910 270524
rect 197446 270512 197452 270524
rect 197504 270512 197510 270564
rect 192938 269152 192944 269204
rect 192996 269192 193002 269204
rect 197446 269192 197452 269204
rect 192996 269164 197452 269192
rect 192996 269152 193002 269164
rect 197446 269152 197452 269164
rect 197504 269152 197510 269204
rect 186130 269084 186136 269136
rect 186188 269124 186194 269136
rect 197354 269124 197360 269136
rect 186188 269096 197360 269124
rect 186188 269084 186194 269096
rect 197354 269084 197360 269096
rect 197412 269084 197418 269136
rect 18598 267724 18604 267776
rect 18656 267764 18662 267776
rect 197354 267764 197360 267776
rect 18656 267736 197360 267764
rect 18656 267724 18662 267736
rect 197354 267724 197360 267736
rect 197412 267724 197418 267776
rect 253198 267724 253204 267776
rect 253256 267764 253262 267776
rect 271138 267764 271144 267776
rect 253256 267736 271144 267764
rect 253256 267724 253262 267736
rect 271138 267724 271144 267736
rect 271196 267724 271202 267776
rect 108298 267656 108304 267708
rect 108356 267696 108362 267708
rect 197446 267696 197452 267708
rect 108356 267668 197452 267696
rect 108356 267656 108362 267668
rect 197446 267656 197452 267668
rect 197504 267656 197510 267708
rect 188338 267588 188344 267640
rect 188396 267628 188402 267640
rect 197354 267628 197360 267640
rect 188396 267600 197360 267628
rect 188396 267588 188402 267600
rect 197354 267588 197360 267600
rect 197412 267588 197418 267640
rect 253750 266432 253756 266484
rect 253808 266472 253814 266484
rect 276750 266472 276756 266484
rect 253808 266444 276756 266472
rect 253808 266432 253814 266444
rect 276750 266432 276756 266444
rect 276808 266432 276814 266484
rect 253290 266364 253296 266416
rect 253348 266404 253354 266416
rect 290090 266404 290096 266416
rect 253348 266376 290096 266404
rect 253348 266364 253354 266376
rect 290090 266364 290096 266376
rect 290148 266364 290154 266416
rect 7558 266296 7564 266348
rect 7616 266336 7622 266348
rect 197354 266336 197360 266348
rect 7616 266308 197360 266336
rect 7616 266296 7622 266308
rect 197354 266296 197360 266308
rect 197412 266296 197418 266348
rect 253750 265004 253756 265056
rect 253808 265044 253814 265056
rect 267274 265044 267280 265056
rect 253808 265016 267280 265044
rect 253808 265004 253814 265016
rect 267274 265004 267280 265016
rect 267332 265004 267338 265056
rect 187602 264936 187608 264988
rect 187660 264976 187666 264988
rect 197446 264976 197452 264988
rect 187660 264948 197452 264976
rect 187660 264936 187666 264948
rect 197446 264936 197452 264948
rect 197504 264936 197510 264988
rect 253842 264936 253848 264988
rect 253900 264976 253906 264988
rect 303706 264976 303712 264988
rect 253900 264948 303712 264976
rect 253900 264936 253906 264948
rect 303706 264936 303712 264948
rect 303764 264936 303770 264988
rect 253750 264868 253756 264920
rect 253808 264908 253814 264920
rect 428458 264908 428464 264920
rect 253808 264880 428464 264908
rect 253808 264868 253814 264880
rect 428458 264868 428464 264880
rect 428516 264868 428522 264920
rect 188706 263644 188712 263696
rect 188764 263684 188770 263696
rect 197354 263684 197360 263696
rect 188764 263656 197360 263684
rect 188764 263644 188770 263656
rect 197354 263644 197360 263656
rect 197412 263644 197418 263696
rect 17218 263576 17224 263628
rect 17276 263616 17282 263628
rect 197446 263616 197452 263628
rect 17276 263588 197452 263616
rect 17276 263576 17282 263588
rect 197446 263576 197452 263588
rect 197504 263576 197510 263628
rect 14458 263508 14464 263560
rect 14516 263548 14522 263560
rect 197354 263548 197360 263560
rect 14516 263520 197360 263548
rect 14516 263508 14522 263520
rect 197354 263508 197360 263520
rect 197412 263508 197418 263560
rect 191650 262216 191656 262268
rect 191708 262256 191714 262268
rect 197354 262256 197360 262268
rect 191708 262228 197360 262256
rect 191708 262216 191714 262228
rect 197354 262216 197360 262228
rect 197412 262216 197418 262268
rect 253750 262216 253756 262268
rect 253808 262256 253814 262268
rect 300854 262256 300860 262268
rect 253808 262228 300860 262256
rect 253808 262216 253814 262228
rect 300854 262216 300860 262228
rect 300912 262216 300918 262268
rect 195698 260924 195704 260976
rect 195756 260964 195762 260976
rect 197538 260964 197544 260976
rect 195756 260936 197544 260964
rect 195756 260924 195762 260936
rect 197538 260924 197544 260936
rect 197596 260924 197602 260976
rect 172422 260856 172428 260908
rect 172480 260896 172486 260908
rect 197446 260896 197452 260908
rect 172480 260868 197452 260896
rect 172480 260856 172486 260868
rect 197446 260856 197452 260868
rect 197504 260856 197510 260908
rect 253382 260856 253388 260908
rect 253440 260896 253446 260908
rect 293954 260896 293960 260908
rect 253440 260868 293960 260896
rect 253440 260856 253446 260868
rect 293954 260856 293960 260868
rect 294012 260856 294018 260908
rect 94498 260788 94504 260840
rect 94556 260828 94562 260840
rect 197354 260828 197360 260840
rect 94556 260800 197360 260828
rect 94556 260788 94562 260800
rect 197354 260788 197360 260800
rect 197412 260788 197418 260840
rect 253198 259496 253204 259548
rect 253256 259536 253262 259548
rect 256786 259536 256792 259548
rect 253256 259508 256792 259536
rect 253256 259496 253262 259508
rect 256786 259496 256792 259508
rect 256844 259496 256850 259548
rect 175182 259428 175188 259480
rect 175240 259468 175246 259480
rect 197354 259468 197360 259480
rect 175240 259440 197360 259468
rect 175240 259428 175246 259440
rect 197354 259428 197360 259440
rect 197412 259428 197418 259480
rect 252830 259428 252836 259480
rect 252888 259468 252894 259480
rect 382918 259468 382924 259480
rect 252888 259440 382924 259468
rect 252888 259428 252894 259440
rect 382918 259428 382924 259440
rect 382976 259428 382982 259480
rect 271230 259360 271236 259412
rect 271288 259400 271294 259412
rect 579614 259400 579620 259412
rect 271288 259372 579620 259400
rect 271288 259360 271294 259372
rect 579614 259360 579620 259372
rect 579672 259360 579678 259412
rect 252554 259020 252560 259072
rect 252612 259060 252618 259072
rect 255498 259060 255504 259072
rect 252612 259032 255504 259060
rect 252612 259020 252618 259032
rect 255498 259020 255504 259032
rect 255556 259020 255562 259072
rect 191742 258272 191748 258324
rect 191800 258312 191806 258324
rect 197446 258312 197452 258324
rect 191800 258284 197452 258312
rect 191800 258272 191806 258284
rect 197446 258272 197452 258284
rect 197504 258272 197510 258324
rect 188798 258068 188804 258120
rect 188856 258108 188862 258120
rect 197354 258108 197360 258120
rect 188856 258080 197360 258108
rect 188856 258068 188862 258080
rect 197354 258068 197360 258080
rect 197412 258068 197418 258120
rect 253842 258068 253848 258120
rect 253900 258108 253906 258120
rect 276842 258108 276848 258120
rect 253900 258080 276848 258108
rect 253900 258068 253906 258080
rect 276842 258068 276848 258080
rect 276900 258068 276906 258120
rect 250346 258000 250352 258052
rect 250404 258040 250410 258052
rect 253750 258040 253756 258052
rect 250404 258012 253756 258040
rect 250404 258000 250410 258012
rect 253750 258000 253756 258012
rect 253808 258000 253814 258052
rect 253014 257524 253020 257576
rect 253072 257564 253078 257576
rect 257430 257564 257436 257576
rect 253072 257536 257436 257564
rect 253072 257524 253078 257536
rect 257430 257524 257436 257536
rect 257488 257524 257494 257576
rect 184658 256776 184664 256828
rect 184716 256816 184722 256828
rect 197354 256816 197360 256828
rect 184716 256788 197360 256816
rect 184716 256776 184722 256788
rect 197354 256776 197360 256788
rect 197412 256776 197418 256828
rect 14458 256708 14464 256760
rect 14516 256748 14522 256760
rect 197446 256748 197452 256760
rect 14516 256720 197452 256748
rect 14516 256708 14522 256720
rect 197446 256708 197452 256720
rect 197504 256708 197510 256760
rect 253106 256640 253112 256692
rect 253164 256680 253170 256692
rect 582374 256680 582380 256692
rect 253164 256652 582380 256680
rect 253164 256640 253170 256652
rect 582374 256640 582380 256652
rect 582432 256640 582438 256692
rect 253750 256572 253756 256624
rect 253808 256612 253814 256624
rect 425698 256612 425704 256624
rect 253808 256584 425704 256612
rect 253808 256572 253814 256584
rect 425698 256572 425704 256584
rect 425756 256572 425762 256624
rect 177850 255280 177856 255332
rect 177908 255320 177914 255332
rect 197446 255320 197452 255332
rect 177908 255292 197452 255320
rect 177908 255280 177914 255292
rect 197446 255280 197452 255292
rect 197504 255280 197510 255332
rect 184842 255212 184848 255264
rect 184900 255252 184906 255264
rect 197354 255252 197360 255264
rect 184900 255224 197360 255252
rect 184900 255212 184906 255224
rect 197354 255212 197360 255224
rect 197412 255212 197418 255264
rect 253014 253988 253020 254040
rect 253072 254028 253078 254040
rect 256878 254028 256884 254040
rect 253072 254000 256884 254028
rect 253072 253988 253078 254000
rect 256878 253988 256884 254000
rect 256936 253988 256942 254040
rect 3142 253920 3148 253972
rect 3200 253960 3206 253972
rect 169018 253960 169024 253972
rect 3200 253932 169024 253960
rect 3200 253920 3206 253932
rect 169018 253920 169024 253932
rect 169076 253920 169082 253972
rect 193030 253920 193036 253972
rect 193088 253960 193094 253972
rect 197354 253960 197360 253972
rect 193088 253932 197360 253960
rect 193088 253920 193094 253932
rect 197354 253920 197360 253932
rect 197412 253920 197418 253972
rect 253750 253920 253756 253972
rect 253808 253960 253814 253972
rect 271230 253960 271236 253972
rect 253808 253932 271236 253960
rect 253808 253920 253814 253932
rect 271230 253920 271236 253932
rect 271288 253920 271294 253972
rect 25498 252560 25504 252612
rect 25556 252600 25562 252612
rect 197354 252600 197360 252612
rect 25556 252572 197360 252600
rect 25556 252560 25562 252572
rect 197354 252560 197360 252572
rect 197412 252560 197418 252612
rect 253842 252560 253848 252612
rect 253900 252600 253906 252612
rect 304994 252600 305000 252612
rect 253900 252572 305000 252600
rect 253900 252560 253906 252572
rect 304994 252560 305000 252572
rect 305052 252560 305058 252612
rect 253750 252492 253756 252544
rect 253808 252532 253814 252544
rect 411898 252532 411904 252544
rect 253808 252504 411904 252532
rect 253808 252492 253814 252504
rect 411898 252492 411904 252504
rect 411956 252492 411962 252544
rect 181990 251268 181996 251320
rect 182048 251308 182054 251320
rect 197446 251308 197452 251320
rect 182048 251280 197452 251308
rect 182048 251268 182054 251280
rect 197446 251268 197452 251280
rect 197504 251268 197510 251320
rect 180610 251200 180616 251252
rect 180668 251240 180674 251252
rect 197354 251240 197360 251252
rect 180668 251212 197360 251240
rect 180668 251200 180674 251212
rect 197354 251200 197360 251212
rect 197412 251200 197418 251252
rect 187326 250452 187332 250504
rect 187384 250492 187390 250504
rect 198090 250492 198096 250504
rect 187384 250464 198096 250492
rect 187384 250452 187390 250464
rect 198090 250452 198096 250464
rect 198148 250452 198154 250504
rect 253474 250452 253480 250504
rect 253532 250492 253538 250504
rect 284294 250492 284300 250504
rect 253532 250464 284300 250492
rect 253532 250452 253538 250464
rect 284294 250452 284300 250464
rect 284352 250452 284358 250504
rect 253382 249976 253388 250028
rect 253440 250016 253446 250028
rect 259638 250016 259644 250028
rect 253440 249988 259644 250016
rect 253440 249976 253446 249988
rect 259638 249976 259644 249988
rect 259696 249976 259702 250028
rect 191558 249772 191564 249824
rect 191616 249812 191622 249824
rect 197446 249812 197452 249824
rect 191616 249784 197452 249812
rect 191616 249772 191622 249784
rect 197446 249772 197452 249784
rect 197504 249772 197510 249824
rect 178678 249704 178684 249756
rect 178736 249744 178742 249756
rect 197354 249744 197360 249756
rect 178736 249716 197360 249744
rect 178736 249704 178742 249716
rect 197354 249704 197360 249716
rect 197412 249704 197418 249756
rect 253750 249704 253756 249756
rect 253808 249744 253814 249756
rect 266998 249744 267004 249756
rect 253808 249716 267004 249744
rect 253808 249704 253814 249716
rect 266998 249704 267004 249716
rect 267056 249704 267062 249756
rect 194502 248684 194508 248736
rect 194560 248724 194566 248736
rect 197354 248724 197360 248736
rect 194560 248696 197360 248724
rect 194560 248684 194566 248696
rect 197354 248684 197360 248696
rect 197412 248684 197418 248736
rect 253750 248412 253756 248464
rect 253808 248452 253814 248464
rect 306374 248452 306380 248464
rect 253808 248424 306380 248452
rect 253808 248412 253814 248424
rect 306374 248412 306380 248424
rect 306432 248412 306438 248464
rect 180702 248344 180708 248396
rect 180760 248384 180766 248396
rect 197446 248384 197452 248396
rect 180760 248356 197452 248384
rect 180760 248344 180766 248356
rect 197446 248344 197452 248356
rect 197504 248344 197510 248396
rect 253842 248344 253848 248396
rect 253900 248384 253906 248396
rect 270494 248384 270500 248396
rect 253900 248356 270500 248384
rect 253900 248344 253906 248356
rect 270494 248344 270500 248356
rect 270552 248344 270558 248396
rect 194410 247052 194416 247104
rect 194468 247092 194474 247104
rect 197538 247092 197544 247104
rect 194468 247064 197544 247092
rect 194468 247052 194474 247064
rect 197538 247052 197544 247064
rect 197596 247052 197602 247104
rect 253750 247052 253756 247104
rect 253808 247092 253814 247104
rect 263778 247092 263784 247104
rect 253808 247064 263784 247092
rect 253808 247052 253814 247064
rect 263778 247052 263784 247064
rect 263836 247052 263842 247104
rect 15838 246984 15844 247036
rect 15896 247024 15902 247036
rect 197354 247024 197360 247036
rect 15896 246996 197360 247024
rect 15896 246984 15902 246996
rect 197354 246984 197360 246996
rect 197412 246984 197418 247036
rect 253750 245624 253756 245676
rect 253808 245664 253814 245676
rect 298186 245664 298192 245676
rect 253808 245636 298192 245664
rect 253808 245624 253814 245636
rect 298186 245624 298192 245636
rect 298244 245624 298250 245676
rect 253842 245556 253848 245608
rect 253900 245596 253906 245608
rect 264238 245596 264244 245608
rect 253900 245568 264244 245596
rect 253900 245556 253906 245568
rect 264238 245556 264244 245568
rect 264296 245556 264302 245608
rect 3602 244876 3608 244928
rect 3660 244916 3666 244928
rect 191098 244916 191104 244928
rect 3660 244888 191104 244916
rect 3660 244876 3666 244888
rect 191098 244876 191104 244888
rect 191156 244876 191162 244928
rect 195606 244264 195612 244316
rect 195664 244304 195670 244316
rect 197446 244304 197452 244316
rect 195664 244276 197452 244304
rect 195664 244264 195670 244276
rect 197446 244264 197452 244276
rect 197504 244264 197510 244316
rect 253750 244264 253756 244316
rect 253808 244304 253814 244316
rect 292850 244304 292856 244316
rect 253808 244276 292856 244304
rect 253808 244264 253814 244276
rect 292850 244264 292856 244276
rect 292908 244264 292914 244316
rect 579890 244304 579896 244316
rect 296686 244276 579896 244304
rect 21358 244196 21364 244248
rect 21416 244236 21422 244248
rect 197354 244236 197360 244248
rect 21416 244208 197360 244236
rect 21416 244196 21422 244208
rect 197354 244196 197360 244208
rect 197412 244196 197418 244248
rect 253382 244196 253388 244248
rect 253440 244236 253446 244248
rect 296686 244236 296714 244276
rect 579890 244264 579896 244276
rect 579948 244264 579954 244316
rect 253440 244208 296714 244236
rect 253440 244196 253446 244208
rect 253750 242972 253756 243024
rect 253808 243012 253814 243024
rect 260098 243012 260104 243024
rect 253808 242984 260104 243012
rect 253808 242972 253814 242984
rect 260098 242972 260104 242984
rect 260156 242972 260162 243024
rect 192846 242836 192852 242888
rect 192904 242876 192910 242888
rect 198734 242876 198740 242888
rect 192904 242848 198740 242876
rect 192904 242836 192910 242848
rect 198734 242836 198740 242848
rect 198792 242836 198798 242888
rect 253750 242836 253756 242888
rect 253808 242876 253814 242888
rect 547138 242876 547144 242888
rect 253808 242848 547144 242876
rect 253808 242836 253814 242848
rect 547138 242836 547144 242848
rect 547196 242836 547202 242888
rect 252554 241544 252560 241596
rect 252612 241584 252618 241596
rect 255498 241584 255504 241596
rect 252612 241556 255504 241584
rect 252612 241544 252618 241556
rect 255498 241544 255504 241556
rect 255556 241544 255562 241596
rect 190178 241476 190184 241528
rect 190236 241516 190242 241528
rect 197354 241516 197360 241528
rect 190236 241488 197360 241516
rect 190236 241476 190242 241488
rect 197354 241476 197360 241488
rect 197412 241476 197418 241528
rect 3050 240116 3056 240168
rect 3108 240156 3114 240168
rect 191834 240156 191840 240168
rect 3108 240128 191840 240156
rect 3108 240116 3114 240128
rect 191834 240116 191840 240128
rect 191892 240116 191898 240168
rect 249058 240116 249064 240168
rect 249116 240156 249122 240168
rect 250254 240156 250260 240168
rect 249116 240128 250260 240156
rect 249116 240116 249122 240128
rect 250254 240116 250260 240128
rect 250312 240116 250318 240168
rect 253750 240116 253756 240168
rect 253808 240156 253814 240168
rect 311894 240156 311900 240168
rect 253808 240128 311900 240156
rect 253808 240116 253814 240128
rect 311894 240116 311900 240128
rect 311952 240116 311958 240168
rect 206010 240048 206016 240100
rect 206068 240088 206074 240100
rect 582466 240088 582472 240100
rect 206068 240060 582472 240088
rect 206068 240048 206074 240060
rect 582466 240048 582472 240060
rect 582524 240048 582530 240100
rect 169018 239980 169024 240032
rect 169076 240020 169082 240032
rect 242710 240020 242716 240032
rect 169076 239992 242716 240020
rect 169076 239980 169082 239992
rect 242710 239980 242716 239992
rect 242768 239980 242774 240032
rect 244006 239980 244012 240032
rect 244064 240020 244070 240032
rect 268378 240020 268384 240032
rect 244064 239992 268384 240020
rect 244064 239980 244070 239992
rect 268378 239980 268384 239992
rect 268436 239980 268442 240032
rect 200758 239912 200764 239964
rect 200816 239952 200822 239964
rect 206370 239952 206376 239964
rect 200816 239924 206376 239952
rect 200816 239912 200822 239924
rect 206370 239912 206376 239924
rect 206428 239912 206434 239964
rect 236914 239912 236920 239964
rect 236972 239952 236978 239964
rect 258718 239952 258724 239964
rect 236972 239924 258724 239952
rect 236972 239912 236978 239924
rect 258718 239912 258724 239924
rect 258776 239912 258782 239964
rect 190546 239844 190552 239896
rect 190604 239884 190610 239896
rect 212442 239884 212448 239896
rect 190604 239856 212448 239884
rect 190604 239844 190610 239856
rect 212442 239844 212448 239856
rect 212500 239844 212506 239896
rect 195790 239776 195796 239828
rect 195848 239816 195854 239828
rect 238754 239816 238760 239828
rect 195848 239788 238760 239816
rect 195848 239776 195854 239788
rect 238754 239776 238760 239788
rect 238812 239776 238818 239828
rect 249242 239776 249248 239828
rect 249300 239816 249306 239828
rect 254118 239816 254124 239828
rect 249300 239788 254124 239816
rect 249300 239776 249306 239788
rect 254118 239776 254124 239788
rect 254176 239776 254182 239828
rect 198734 239368 198740 239420
rect 198792 239408 198798 239420
rect 215938 239408 215944 239420
rect 198792 239380 215944 239408
rect 198792 239368 198798 239380
rect 215938 239368 215944 239380
rect 215996 239368 216002 239420
rect 245010 239368 245016 239420
rect 245068 239408 245074 239420
rect 252738 239408 252744 239420
rect 245068 239380 252744 239408
rect 245068 239368 245074 239380
rect 252738 239368 252744 239380
rect 252796 239368 252802 239420
rect 246298 238756 246304 238808
rect 246356 238796 246362 238808
rect 250162 238796 250168 238808
rect 246356 238768 250168 238796
rect 246356 238756 246362 238768
rect 250162 238756 250168 238768
rect 250220 238756 250226 238808
rect 177942 238688 177948 238740
rect 178000 238728 178006 238740
rect 211798 238728 211804 238740
rect 178000 238700 211804 238728
rect 178000 238688 178006 238700
rect 211798 238688 211804 238700
rect 211856 238688 211862 238740
rect 222102 238688 222108 238740
rect 222160 238728 222166 238740
rect 583110 238728 583116 238740
rect 222160 238700 583116 238728
rect 222160 238688 222166 238700
rect 583110 238688 583116 238700
rect 583168 238688 583174 238740
rect 191098 238620 191104 238672
rect 191156 238660 191162 238672
rect 216950 238660 216956 238672
rect 191156 238632 216956 238660
rect 191156 238620 191162 238632
rect 216950 238620 216956 238632
rect 217008 238620 217014 238672
rect 221458 238620 221464 238672
rect 221516 238660 221522 238672
rect 574738 238660 574744 238672
rect 221516 238632 574744 238660
rect 221516 238620 221522 238632
rect 574738 238620 574744 238632
rect 574796 238620 574802 238672
rect 228542 238552 228548 238604
rect 228600 238592 228606 238604
rect 359458 238592 359464 238604
rect 228600 238564 359464 238592
rect 228600 238552 228606 238564
rect 359458 238552 359464 238564
rect 359516 238552 359522 238604
rect 191834 238484 191840 238536
rect 191892 238524 191898 238536
rect 233694 238524 233700 238536
rect 191892 238496 233700 238524
rect 191892 238484 191898 238496
rect 233694 238484 233700 238496
rect 233752 238484 233758 238536
rect 247218 238484 247224 238536
rect 247276 238524 247282 238536
rect 269758 238524 269764 238536
rect 247276 238496 269764 238524
rect 247276 238484 247282 238496
rect 269758 238484 269764 238496
rect 269816 238484 269822 238536
rect 173158 238416 173164 238468
rect 173216 238456 173222 238468
rect 229186 238456 229192 238468
rect 173216 238428 229192 238456
rect 173216 238416 173222 238428
rect 229186 238416 229192 238428
rect 229244 238416 229250 238468
rect 235626 238076 235632 238128
rect 235684 238116 235690 238128
rect 266998 238116 267004 238128
rect 235684 238088 267004 238116
rect 235684 238076 235690 238088
rect 266998 238076 267004 238088
rect 267056 238076 267062 238128
rect 218882 238008 218888 238060
rect 218940 238048 218946 238060
rect 300946 238048 300952 238060
rect 218940 238020 300952 238048
rect 218940 238008 218946 238020
rect 300946 238008 300952 238020
rect 301004 238008 301010 238060
rect 202782 237804 202788 237856
rect 202840 237844 202846 237856
rect 205542 237844 205548 237856
rect 202840 237816 205548 237844
rect 202840 237804 202846 237816
rect 205542 237804 205548 237816
rect 205600 237804 205606 237856
rect 200206 237396 200212 237448
rect 200264 237436 200270 237448
rect 206278 237436 206284 237448
rect 200264 237408 206284 237436
rect 200264 237396 200270 237408
rect 206278 237396 206284 237408
rect 206336 237396 206342 237448
rect 233050 237396 233056 237448
rect 233108 237436 233114 237448
rect 237374 237436 237380 237448
rect 233108 237408 237380 237436
rect 233108 237396 233114 237408
rect 237374 237396 237380 237408
rect 237432 237396 237438 237448
rect 245286 237328 245292 237380
rect 245344 237368 245350 237380
rect 582558 237368 582564 237380
rect 245344 237340 582564 237368
rect 245344 237328 245350 237340
rect 582558 237328 582564 237340
rect 582616 237328 582622 237380
rect 244918 236716 244924 236768
rect 244976 236756 244982 236768
rect 251082 236756 251088 236768
rect 244976 236728 251088 236756
rect 244976 236716 244982 236728
rect 251082 236716 251088 236728
rect 251140 236716 251146 236768
rect 199838 236648 199844 236700
rect 199896 236688 199902 236700
rect 281626 236688 281632 236700
rect 199896 236660 281632 236688
rect 199896 236648 199902 236660
rect 281626 236648 281632 236660
rect 281684 236648 281690 236700
rect 205542 235900 205548 235952
rect 205600 235940 205606 235952
rect 582926 235940 582932 235952
rect 205600 235912 582932 235940
rect 205600 235900 205606 235912
rect 582926 235900 582932 235912
rect 582984 235900 582990 235952
rect 166258 235832 166264 235884
rect 166316 235872 166322 235884
rect 244642 235872 244648 235884
rect 166316 235844 244648 235872
rect 166316 235832 166322 235844
rect 244642 235832 244648 235844
rect 244700 235832 244706 235884
rect 242158 235356 242164 235408
rect 242216 235396 242222 235408
rect 252830 235396 252836 235408
rect 242216 235368 252836 235396
rect 242216 235356 242222 235368
rect 252830 235356 252836 235368
rect 252888 235356 252894 235408
rect 243538 235288 243544 235340
rect 243596 235328 243602 235340
rect 265066 235328 265072 235340
rect 243596 235300 265072 235328
rect 243596 235288 243602 235300
rect 265066 235288 265072 235300
rect 265124 235288 265130 235340
rect 247862 235220 247868 235272
rect 247920 235260 247926 235272
rect 322198 235260 322204 235272
rect 247920 235232 322204 235260
rect 247920 235220 247926 235232
rect 322198 235220 322204 235232
rect 322256 235220 322262 235272
rect 237558 234540 237564 234592
rect 237616 234580 237622 234592
rect 542354 234580 542360 234592
rect 237616 234552 542360 234580
rect 237616 234540 237622 234552
rect 542354 234540 542360 234552
rect 542412 234540 542418 234592
rect 253842 233928 253848 233980
rect 253900 233968 253906 233980
rect 255498 233968 255504 233980
rect 253900 233940 255504 233968
rect 253900 233928 253906 233940
rect 255498 233928 255504 233940
rect 255556 233928 255562 233980
rect 188706 233860 188712 233912
rect 188764 233900 188770 233912
rect 306466 233900 306472 233912
rect 188764 233872 306472 233900
rect 188764 233860 188770 233872
rect 306466 233860 306472 233872
rect 306524 233860 306530 233912
rect 231118 233180 231124 233232
rect 231176 233220 231182 233232
rect 233234 233220 233240 233232
rect 231176 233192 233240 233220
rect 231176 233180 231182 233192
rect 233234 233180 233240 233192
rect 233292 233180 233298 233232
rect 566458 233180 566464 233232
rect 566516 233220 566522 233232
rect 580166 233220 580172 233232
rect 566516 233192 580172 233220
rect 566516 233180 566522 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 249794 232636 249800 232688
rect 249852 232676 249858 232688
rect 287146 232676 287152 232688
rect 249852 232648 287152 232676
rect 249852 232636 249858 232648
rect 287146 232636 287152 232648
rect 287204 232636 287210 232688
rect 191098 232568 191104 232620
rect 191156 232608 191162 232620
rect 254210 232608 254216 232620
rect 191156 232580 254216 232608
rect 191156 232568 191162 232580
rect 254210 232568 254216 232580
rect 254268 232568 254274 232620
rect 206646 232500 206652 232552
rect 206704 232540 206710 232552
rect 302878 232540 302884 232552
rect 206704 232512 302884 232540
rect 206704 232500 206710 232512
rect 302878 232500 302884 232512
rect 302936 232500 302942 232552
rect 200850 231072 200856 231124
rect 200908 231112 200914 231124
rect 284478 231112 284484 231124
rect 200908 231084 284484 231112
rect 200908 231072 200914 231084
rect 284478 231072 284484 231084
rect 284536 231072 284542 231124
rect 190086 228420 190092 228472
rect 190144 228460 190150 228472
rect 269758 228460 269764 228472
rect 190144 228432 269764 228460
rect 190144 228420 190150 228432
rect 269758 228420 269764 228432
rect 269816 228420 269822 228472
rect 21358 228352 21364 228404
rect 21416 228392 21422 228404
rect 213730 228392 213736 228404
rect 21416 228364 213736 228392
rect 21416 228352 21422 228364
rect 213730 228352 213736 228364
rect 213788 228352 213794 228404
rect 230474 225700 230480 225752
rect 230532 225740 230538 225752
rect 231854 225740 231860 225752
rect 230532 225712 231860 225740
rect 230532 225700 230538 225712
rect 231854 225700 231860 225712
rect 231912 225700 231918 225752
rect 196986 225564 196992 225616
rect 197044 225604 197050 225616
rect 230474 225604 230480 225616
rect 197044 225576 230480 225604
rect 197044 225564 197050 225576
rect 230474 225564 230480 225576
rect 230532 225564 230538 225616
rect 235258 225564 235264 225616
rect 235316 225604 235322 225616
rect 252646 225604 252652 225616
rect 235316 225576 252652 225604
rect 235316 225564 235322 225576
rect 252646 225564 252652 225576
rect 252704 225564 252710 225616
rect 200022 224204 200028 224256
rect 200080 224244 200086 224256
rect 230566 224244 230572 224256
rect 200080 224216 230572 224244
rect 200080 224204 200086 224216
rect 230566 224204 230572 224216
rect 230624 224204 230630 224256
rect 231762 223524 231768 223576
rect 231820 223564 231826 223576
rect 233326 223564 233332 223576
rect 231820 223536 233332 223564
rect 231820 223524 231826 223536
rect 233326 223524 233332 223536
rect 233384 223524 233390 223576
rect 199930 222844 199936 222896
rect 199988 222884 199994 222896
rect 230658 222884 230664 222896
rect 199988 222856 230664 222884
rect 199988 222844 199994 222856
rect 230658 222844 230664 222856
rect 230716 222844 230722 222896
rect 7558 220056 7564 220108
rect 7616 220096 7622 220108
rect 240778 220096 240784 220108
rect 7616 220068 240784 220096
rect 7616 220056 7622 220068
rect 240778 220056 240784 220068
rect 240836 220056 240842 220108
rect 4798 218696 4804 218748
rect 4856 218736 4862 218748
rect 240134 218736 240140 218748
rect 4856 218708 240140 218736
rect 4856 218696 4862 218708
rect 240134 218696 240140 218708
rect 240192 218696 240198 218748
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 17218 215268 17224 215280
rect 3384 215240 17224 215268
rect 3384 215228 3390 215240
rect 17218 215228 17224 215240
rect 17276 215228 17282 215280
rect 211154 211760 211160 211812
rect 211212 211800 211218 211812
rect 287238 211800 287244 211812
rect 211212 211772 287244 211800
rect 211212 211760 211218 211772
rect 287238 211760 287244 211772
rect 287296 211760 287302 211812
rect 257338 206932 257344 206984
rect 257396 206972 257402 206984
rect 579890 206972 579896 206984
rect 257396 206944 579896 206972
rect 257396 206932 257402 206944
rect 579890 206932 579896 206944
rect 579948 206932 579954 206984
rect 198550 206252 198556 206304
rect 198608 206292 198614 206304
rect 285766 206292 285772 206304
rect 198608 206264 285772 206292
rect 198608 206252 198614 206264
rect 285766 206252 285772 206264
rect 285824 206252 285830 206304
rect 195698 204892 195704 204944
rect 195756 204932 195762 204944
rect 281718 204932 281724 204944
rect 195756 204904 281724 204932
rect 195756 204892 195762 204904
rect 281718 204892 281724 204904
rect 281776 204892 281782 204944
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 259638 202824 259644 202836
rect 3108 202796 259644 202824
rect 3108 202784 3114 202796
rect 259638 202784 259644 202796
rect 259696 202784 259702 202836
rect 229830 202104 229836 202156
rect 229888 202144 229894 202156
rect 284570 202144 284576 202156
rect 229888 202116 284576 202144
rect 229888 202104 229894 202116
rect 284570 202104 284576 202116
rect 284628 202104 284634 202156
rect 215018 200744 215024 200796
rect 215076 200784 215082 200796
rect 287330 200784 287336 200796
rect 215076 200756 287336 200784
rect 215076 200744 215082 200756
rect 287330 200744 287336 200756
rect 287388 200744 287394 200796
rect 202138 196596 202144 196648
rect 202196 196636 202202 196648
rect 280154 196636 280160 196648
rect 202196 196608 280160 196636
rect 202196 196596 202202 196608
rect 280154 196596 280160 196608
rect 280212 196596 280218 196648
rect 181990 195236 181996 195288
rect 182048 195276 182054 195288
rect 292758 195276 292764 195288
rect 182048 195248 292764 195276
rect 182048 195236 182054 195248
rect 292758 195236 292764 195248
rect 292816 195236 292822 195288
rect 234338 193808 234344 193860
rect 234396 193848 234402 193860
rect 305086 193848 305092 193860
rect 234396 193820 305092 193848
rect 234396 193808 234402 193820
rect 305086 193808 305092 193820
rect 305144 193808 305150 193860
rect 188890 193128 188896 193180
rect 188948 193168 188954 193180
rect 580166 193168 580172 193180
rect 188948 193140 580172 193168
rect 188948 193128 188954 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 224034 191156 224040 191208
rect 224092 191196 224098 191208
rect 233418 191196 233424 191208
rect 224092 191168 233424 191196
rect 224092 191156 224098 191168
rect 233418 191156 233424 191168
rect 233476 191156 233482 191208
rect 217594 191088 217600 191140
rect 217652 191128 217658 191140
rect 299658 191128 299664 191140
rect 217652 191100 299664 191128
rect 217652 191088 217658 191100
rect 299658 191088 299664 191100
rect 299716 191088 299722 191140
rect 172422 189864 172428 189916
rect 172480 189904 172486 189916
rect 288618 189904 288624 189916
rect 172480 189876 288624 189904
rect 172480 189864 172486 189876
rect 288618 189864 288624 189876
rect 288676 189864 288682 189916
rect 175182 189796 175188 189848
rect 175240 189836 175246 189848
rect 295518 189836 295524 189848
rect 175240 189808 295524 189836
rect 175240 189796 175246 189808
rect 295518 189796 295524 189808
rect 295576 189796 295582 189848
rect 177850 189728 177856 189780
rect 177908 189768 177914 189780
rect 299750 189768 299756 189780
rect 177908 189740 299756 189768
rect 177908 189728 177914 189740
rect 299750 189728 299756 189740
rect 299808 189728 299814 189780
rect 245930 188436 245936 188488
rect 245988 188476 245994 188488
rect 284386 188476 284392 188488
rect 245988 188448 284392 188476
rect 245988 188436 245994 188448
rect 284386 188436 284392 188448
rect 284444 188436 284450 188488
rect 210510 188368 210516 188420
rect 210568 188408 210574 188420
rect 276934 188408 276940 188420
rect 210568 188380 276940 188408
rect 210568 188368 210574 188380
rect 276934 188368 276940 188380
rect 276992 188368 276998 188420
rect 184658 188300 184664 188352
rect 184716 188340 184722 188352
rect 296898 188340 296904 188352
rect 184716 188312 296904 188340
rect 184716 188300 184722 188312
rect 296898 188300 296904 188312
rect 296956 188300 296962 188352
rect 236270 187008 236276 187060
rect 236328 187048 236334 187060
rect 292666 187048 292672 187060
rect 236328 187020 292672 187048
rect 236328 187008 236334 187020
rect 292666 187008 292672 187020
rect 292724 187008 292730 187060
rect 238846 186940 238852 186992
rect 238904 186980 238910 186992
rect 303798 186980 303804 186992
rect 238904 186952 303804 186980
rect 238904 186940 238910 186952
rect 303798 186940 303804 186952
rect 303856 186940 303862 186992
rect 190270 185852 190276 185904
rect 190328 185892 190334 185904
rect 235994 185892 236000 185904
rect 190328 185864 236000 185892
rect 190328 185852 190334 185864
rect 235994 185852 236000 185864
rect 236052 185852 236058 185904
rect 186222 185784 186228 185836
rect 186280 185824 186286 185836
rect 240226 185824 240232 185836
rect 186280 185796 240232 185824
rect 186280 185784 186286 185796
rect 240226 185784 240232 185796
rect 240284 185784 240290 185836
rect 201494 185716 201500 185768
rect 201552 185756 201558 185768
rect 231946 185756 231952 185768
rect 201552 185728 231952 185756
rect 201552 185716 201558 185728
rect 231946 185716 231952 185728
rect 232004 185716 232010 185768
rect 232406 185716 232412 185768
rect 232464 185756 232470 185768
rect 294138 185756 294144 185768
rect 232464 185728 294144 185756
rect 232464 185716 232470 185728
rect 294138 185716 294144 185728
rect 294196 185716 294202 185768
rect 184750 185648 184756 185700
rect 184808 185688 184814 185700
rect 291378 185688 291384 185700
rect 184808 185660 291384 185688
rect 184808 185648 184814 185660
rect 291378 185648 291384 185660
rect 291436 185648 291442 185700
rect 3510 185580 3516 185632
rect 3568 185620 3574 185632
rect 193858 185620 193864 185632
rect 3568 185592 193864 185620
rect 3568 185580 3574 185592
rect 193858 185580 193864 185592
rect 193916 185580 193922 185632
rect 223390 185580 223396 185632
rect 223448 185620 223454 185632
rect 285858 185620 285864 185632
rect 223448 185592 285864 185620
rect 223448 185580 223454 185592
rect 285858 185580 285864 185592
rect 285916 185580 285922 185632
rect 197262 184288 197268 184340
rect 197320 184328 197326 184340
rect 230750 184328 230756 184340
rect 197320 184300 230756 184328
rect 197320 184288 197326 184300
rect 230750 184288 230756 184300
rect 230808 184288 230814 184340
rect 278130 184288 278136 184340
rect 278188 184328 278194 184340
rect 307754 184328 307760 184340
rect 278188 184300 307760 184328
rect 278188 184288 278194 184300
rect 307754 184288 307760 184300
rect 307812 184288 307818 184340
rect 227898 184220 227904 184272
rect 227956 184260 227962 184272
rect 288434 184260 288440 184272
rect 227956 184232 288440 184260
rect 227956 184220 227962 184232
rect 288434 184220 288440 184232
rect 288492 184220 288498 184272
rect 225322 184152 225328 184204
rect 225380 184192 225386 184204
rect 289906 184192 289912 184204
rect 225380 184164 289912 184192
rect 225380 184152 225386 184164
rect 289906 184152 289912 184164
rect 289964 184152 289970 184204
rect 100662 183540 100668 183592
rect 100720 183580 100726 183592
rect 209038 183580 209044 183592
rect 100720 183552 209044 183580
rect 100720 183540 100726 183552
rect 209038 183540 209044 183552
rect 209096 183540 209102 183592
rect 220170 183132 220176 183184
rect 220228 183172 220234 183184
rect 232130 183172 232136 183184
rect 220228 183144 232136 183172
rect 220228 183132 220234 183144
rect 232130 183132 232136 183144
rect 232188 183132 232194 183184
rect 191650 183064 191656 183116
rect 191708 183104 191714 183116
rect 234614 183104 234620 183116
rect 191708 183076 234620 183104
rect 191708 183064 191714 183076
rect 234614 183064 234620 183076
rect 234672 183064 234678 183116
rect 188982 182996 188988 183048
rect 189040 183036 189046 183048
rect 244366 183036 244372 183048
rect 189040 183008 244372 183036
rect 189040 182996 189046 183008
rect 244366 182996 244372 183008
rect 244424 182996 244430 183048
rect 187326 182928 187332 182980
rect 187384 182968 187390 182980
rect 247034 182968 247040 182980
rect 187384 182940 247040 182968
rect 187384 182928 187390 182940
rect 247034 182928 247040 182940
rect 247092 182928 247098 182980
rect 214374 182860 214380 182912
rect 214432 182900 214438 182912
rect 298278 182900 298284 182912
rect 214432 182872 298284 182900
rect 214432 182860 214438 182872
rect 298278 182860 298284 182872
rect 298336 182860 298342 182912
rect 203426 182792 203432 182844
rect 203484 182832 203490 182844
rect 296990 182832 296996 182844
rect 203484 182804 296996 182832
rect 203484 182792 203490 182804
rect 296990 182792 296996 182804
rect 297048 182792 297054 182844
rect 127066 182384 127072 182436
rect 127124 182424 127130 182436
rect 170582 182424 170588 182436
rect 127124 182396 170588 182424
rect 127124 182384 127130 182396
rect 170582 182384 170588 182396
rect 170640 182384 170646 182436
rect 108114 182316 108120 182368
rect 108172 182356 108178 182368
rect 169018 182356 169024 182368
rect 108172 182328 169024 182356
rect 108172 182316 108178 182328
rect 169018 182316 169024 182328
rect 169076 182316 169082 182368
rect 105906 182248 105912 182300
rect 105964 182288 105970 182300
rect 167638 182288 167644 182300
rect 105964 182260 167644 182288
rect 105964 182248 105970 182260
rect 167638 182248 167644 182260
rect 167696 182248 167702 182300
rect 130746 182180 130752 182232
rect 130804 182220 130810 182232
rect 204898 182220 204904 182232
rect 130804 182192 204904 182220
rect 130804 182180 130810 182192
rect 204898 182180 204904 182192
rect 204956 182180 204962 182232
rect 215662 181432 215668 181484
rect 215720 181472 215726 181484
rect 232038 181472 232044 181484
rect 215720 181444 232044 181472
rect 215720 181432 215726 181444
rect 232038 181432 232044 181444
rect 232096 181432 232102 181484
rect 243354 181432 243360 181484
rect 243412 181472 243418 181484
rect 295426 181472 295432 181484
rect 243412 181444 295432 181472
rect 243412 181432 243418 181444
rect 295426 181432 295432 181444
rect 295484 181432 295490 181484
rect 132402 181092 132408 181144
rect 132460 181132 132466 181144
rect 166534 181132 166540 181144
rect 132460 181104 166540 181132
rect 132460 181092 132466 181104
rect 166534 181092 166540 181104
rect 166592 181092 166598 181144
rect 124950 181024 124956 181076
rect 125008 181064 125014 181076
rect 167822 181064 167828 181076
rect 125008 181036 167828 181064
rect 125008 181024 125014 181036
rect 167822 181024 167828 181036
rect 167880 181024 167886 181076
rect 103330 180956 103336 181008
rect 103388 180996 103394 181008
rect 166258 180996 166264 181008
rect 103388 180968 166264 180996
rect 103388 180956 103394 180968
rect 166258 180956 166264 180968
rect 166316 180956 166322 181008
rect 114462 180888 114468 180940
rect 114520 180928 114526 180940
rect 178678 180928 178684 180940
rect 114520 180900 178684 180928
rect 114520 180888 114526 180900
rect 178678 180888 178684 180900
rect 178736 180888 178742 180940
rect 119522 180820 119528 180872
rect 119580 180860 119586 180872
rect 213270 180860 213276 180872
rect 119580 180832 213276 180860
rect 119580 180820 119586 180832
rect 213270 180820 213276 180832
rect 213328 180820 213334 180872
rect 180518 180412 180524 180464
rect 180576 180452 180582 180464
rect 227622 180452 227628 180464
rect 180576 180424 227628 180452
rect 180576 180412 180582 180424
rect 227622 180412 227628 180424
rect 227680 180412 227686 180464
rect 190178 180344 190184 180396
rect 190236 180384 190242 180396
rect 237466 180384 237472 180396
rect 190236 180356 237472 180384
rect 190236 180344 190242 180356
rect 237466 180344 237472 180356
rect 237524 180344 237530 180396
rect 187418 180276 187424 180328
rect 187476 180316 187482 180328
rect 234706 180316 234712 180328
rect 187476 180288 234712 180316
rect 187476 180276 187482 180288
rect 234706 180276 234712 180288
rect 234764 180276 234770 180328
rect 276750 180276 276756 180328
rect 276808 180316 276814 180328
rect 288710 180316 288716 180328
rect 276808 180288 288716 180316
rect 276808 180276 276814 180288
rect 288710 180276 288716 180288
rect 288768 180276 288774 180328
rect 226610 180208 226616 180260
rect 226668 180248 226674 180260
rect 280338 180248 280344 180260
rect 226668 180220 280344 180248
rect 226668 180208 226674 180220
rect 280338 180208 280344 180220
rect 280396 180208 280402 180260
rect 188798 180140 188804 180192
rect 188856 180180 188862 180192
rect 242986 180180 242992 180192
rect 188856 180152 242992 180180
rect 188856 180140 188862 180152
rect 242986 180140 242992 180152
rect 243044 180140 243050 180192
rect 272518 180140 272524 180192
rect 272576 180180 272582 180192
rect 301038 180180 301044 180192
rect 272576 180152 301044 180180
rect 272576 180140 272582 180152
rect 301038 180140 301044 180152
rect 301096 180140 301102 180192
rect 224678 180072 224684 180124
rect 224736 180112 224742 180124
rect 291286 180112 291292 180124
rect 224736 180084 291292 180112
rect 224736 180072 224742 180084
rect 291286 180072 291292 180084
rect 291344 180072 291350 180124
rect 123754 179596 123760 179648
rect 123812 179636 123818 179648
rect 169202 179636 169208 179648
rect 123812 179608 169208 179636
rect 123812 179596 123818 179608
rect 169202 179596 169208 179608
rect 169260 179596 169266 179648
rect 97534 179528 97540 179580
rect 97592 179568 97598 179580
rect 173158 179568 173164 179580
rect 97592 179540 173164 179568
rect 97592 179528 97598 179540
rect 173158 179528 173164 179540
rect 173216 179528 173222 179580
rect 129458 179460 129464 179512
rect 129516 179500 129522 179512
rect 214190 179500 214196 179512
rect 129516 179472 214196 179500
rect 129516 179460 129522 179472
rect 214190 179460 214196 179472
rect 214248 179460 214254 179512
rect 114370 179392 114376 179444
rect 114428 179432 114434 179444
rect 211798 179432 211804 179444
rect 114428 179404 211804 179432
rect 114428 179392 114434 179404
rect 211798 179392 211804 179404
rect 211856 179392 211862 179444
rect 218238 178916 218244 178968
rect 218296 178956 218302 178968
rect 229094 178956 229100 178968
rect 218296 178928 229100 178956
rect 218296 178916 218302 178928
rect 229094 178916 229100 178928
rect 229152 178916 229158 178968
rect 208578 178848 208584 178900
rect 208636 178888 208642 178900
rect 238846 178888 238852 178900
rect 208636 178860 238852 178888
rect 208636 178848 208642 178860
rect 238846 178848 238852 178860
rect 238904 178848 238910 178900
rect 273898 178848 273904 178900
rect 273956 178888 273962 178900
rect 295610 178888 295616 178900
rect 273956 178860 295616 178888
rect 273956 178848 273962 178860
rect 295610 178848 295616 178860
rect 295668 178848 295674 178900
rect 191558 178780 191564 178832
rect 191616 178820 191622 178832
rect 244274 178820 244280 178832
rect 191616 178792 244280 178820
rect 191616 178780 191622 178792
rect 244274 178780 244280 178792
rect 244332 178780 244338 178832
rect 271138 178780 271144 178832
rect 271196 178820 271202 178832
rect 294046 178820 294052 178832
rect 271196 178792 294052 178820
rect 271196 178780 271202 178792
rect 294046 178780 294052 178792
rect 294104 178780 294110 178832
rect 206278 178712 206284 178764
rect 206336 178752 206342 178764
rect 291470 178752 291476 178764
rect 206336 178724 291476 178752
rect 206336 178712 206342 178724
rect 291470 178712 291476 178724
rect 291528 178712 291534 178764
rect 204070 178644 204076 178696
rect 204128 178684 204134 178696
rect 301130 178684 301136 178696
rect 204128 178656 301136 178684
rect 204128 178644 204134 178656
rect 301130 178644 301136 178656
rect 301188 178644 301194 178696
rect 118418 178304 118424 178356
rect 118476 178344 118482 178356
rect 166350 178344 166356 178356
rect 118476 178316 166356 178344
rect 118476 178304 118482 178316
rect 166350 178304 166356 178316
rect 166408 178304 166414 178356
rect 110690 178236 110696 178288
rect 110748 178276 110754 178288
rect 169110 178276 169116 178288
rect 110748 178248 169116 178276
rect 110748 178236 110754 178248
rect 169110 178236 169116 178248
rect 169168 178236 169174 178288
rect 112254 178168 112260 178220
rect 112312 178208 112318 178220
rect 177298 178208 177304 178220
rect 112312 178180 177304 178208
rect 112312 178168 112318 178180
rect 177298 178168 177304 178180
rect 177356 178168 177362 178220
rect 133138 178100 133144 178152
rect 133196 178140 133202 178152
rect 214006 178140 214012 178152
rect 133196 178112 214012 178140
rect 133196 178100 133202 178112
rect 214006 178100 214012 178112
rect 214064 178100 214070 178152
rect 109586 178032 109592 178084
rect 109644 178072 109650 178084
rect 213178 178072 213184 178084
rect 109644 178044 213184 178072
rect 109644 178032 109650 178044
rect 213178 178032 213184 178044
rect 213236 178032 213242 178084
rect 227254 177964 227260 178016
rect 227312 178004 227318 178016
rect 229186 178004 229192 178016
rect 227312 177976 229192 178004
rect 227312 177964 227318 177976
rect 229186 177964 229192 177976
rect 229244 177964 229250 178016
rect 268470 177964 268476 178016
rect 268528 178004 268534 178016
rect 296622 178004 296628 178016
rect 268528 177976 296628 178004
rect 268528 177964 268534 177976
rect 296622 177964 296628 177976
rect 296680 177964 296686 178016
rect 222746 177488 222752 177540
rect 222804 177528 222810 177540
rect 236086 177528 236092 177540
rect 222804 177500 236092 177528
rect 222804 177488 222810 177500
rect 236086 177488 236092 177500
rect 236144 177488 236150 177540
rect 220814 177420 220820 177472
rect 220872 177460 220878 177472
rect 238754 177460 238760 177472
rect 220872 177432 238760 177460
rect 220872 177420 220878 177432
rect 238754 177420 238760 177432
rect 238812 177420 238818 177472
rect 271230 177420 271236 177472
rect 271288 177460 271294 177472
rect 288526 177460 288532 177472
rect 271288 177432 288532 177460
rect 271288 177420 271294 177432
rect 288526 177420 288532 177432
rect 288584 177420 288590 177472
rect 194410 177352 194416 177404
rect 194468 177392 194474 177404
rect 236270 177392 236276 177404
rect 194468 177364 236276 177392
rect 194468 177352 194474 177364
rect 236270 177352 236276 177364
rect 236328 177352 236334 177404
rect 276842 177352 276848 177404
rect 276900 177392 276906 177404
rect 302326 177392 302332 177404
rect 276900 177364 302332 177392
rect 276900 177352 276906 177364
rect 302326 177352 302332 177364
rect 302384 177352 302390 177404
rect 195606 177284 195612 177336
rect 195664 177324 195670 177336
rect 292574 177324 292580 177336
rect 195664 177296 292580 177324
rect 195664 177284 195670 177296
rect 292574 177284 292580 177296
rect 292632 177284 292638 177336
rect 128170 177012 128176 177064
rect 128228 177052 128234 177064
rect 214098 177052 214104 177064
rect 128228 177024 214104 177052
rect 128228 177012 128234 177024
rect 214098 177012 214104 177024
rect 214156 177012 214162 177064
rect 107010 176944 107016 176996
rect 107068 176984 107074 176996
rect 165338 176984 165344 176996
rect 107068 176956 165344 176984
rect 107068 176944 107074 176956
rect 165338 176944 165344 176956
rect 165396 176944 165402 176996
rect 148226 176876 148232 176928
rect 148284 176916 148290 176928
rect 214558 176916 214564 176928
rect 148284 176888 214564 176916
rect 148284 176876 148290 176888
rect 214558 176876 214564 176888
rect 214616 176876 214622 176928
rect 104618 176808 104624 176860
rect 104676 176848 104682 176860
rect 170490 176848 170496 176860
rect 104676 176820 170496 176848
rect 104676 176808 104682 176820
rect 170490 176808 170496 176820
rect 170548 176808 170554 176860
rect 125870 176740 125876 176792
rect 125928 176780 125934 176792
rect 197998 176780 198004 176792
rect 125928 176752 198004 176780
rect 125928 176740 125934 176752
rect 197998 176740 198004 176752
rect 198056 176740 198062 176792
rect 136082 176672 136088 176724
rect 136140 176712 136146 176724
rect 136140 176684 136772 176712
rect 136140 176672 136146 176684
rect 136744 176644 136772 176684
rect 158990 176672 158996 176724
rect 159048 176712 159054 176724
rect 165430 176712 165436 176724
rect 159048 176684 165436 176712
rect 159048 176672 159054 176684
rect 165430 176672 165436 176684
rect 165488 176672 165494 176724
rect 213914 176644 213920 176656
rect 136744 176616 213920 176644
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 134426 176196 134432 176248
rect 134484 176236 134490 176248
rect 165522 176236 165528 176248
rect 134484 176208 165528 176236
rect 134484 176196 134490 176208
rect 165522 176196 165528 176208
rect 165580 176196 165586 176248
rect 121914 176128 121920 176180
rect 121972 176168 121978 176180
rect 166442 176168 166448 176180
rect 121972 176140 166448 176168
rect 121972 176128 121978 176140
rect 166442 176128 166448 176140
rect 166500 176128 166506 176180
rect 194502 176128 194508 176180
rect 194560 176168 194566 176180
rect 242894 176168 242900 176180
rect 194560 176140 242900 176168
rect 194560 176128 194566 176140
rect 242894 176128 242900 176140
rect 242952 176128 242958 176180
rect 276658 176128 276664 176180
rect 276716 176168 276722 176180
rect 279326 176168 279332 176180
rect 276716 176140 279332 176168
rect 276716 176128 276722 176140
rect 279326 176128 279332 176140
rect 279384 176128 279390 176180
rect 116946 176060 116952 176112
rect 117004 176100 117010 176112
rect 169294 176100 169300 176112
rect 117004 176072 169300 176100
rect 117004 176060 117010 176072
rect 169294 176060 169300 176072
rect 169352 176060 169358 176112
rect 187510 176060 187516 176112
rect 187568 176100 187574 176112
rect 236178 176100 236184 176112
rect 187568 176072 236184 176100
rect 187568 176060 187574 176072
rect 236178 176060 236184 176072
rect 236236 176060 236242 176112
rect 278038 176060 278044 176112
rect 278096 176100 278102 176112
rect 289998 176100 290004 176112
rect 278096 176072 290004 176100
rect 278096 176060 278102 176072
rect 289998 176060 290004 176072
rect 290056 176060 290062 176112
rect 120810 175992 120816 176044
rect 120868 176032 120874 176044
rect 180058 176032 180064 176044
rect 120868 176004 180064 176032
rect 120868 175992 120874 176004
rect 180058 175992 180064 176004
rect 180116 175992 180122 176044
rect 183462 175992 183468 176044
rect 183520 176032 183526 176044
rect 237558 176032 237564 176044
rect 183520 176004 237564 176032
rect 183520 175992 183526 176004
rect 237558 175992 237564 176004
rect 237616 175992 237622 176044
rect 276934 175992 276940 176044
rect 276992 176032 276998 176044
rect 289814 176032 289820 176044
rect 276992 176004 289820 176032
rect 276992 175992 276998 176004
rect 289814 175992 289820 176004
rect 289872 175992 289878 176044
rect 115750 175924 115756 175976
rect 115808 175964 115814 175976
rect 211890 175964 211896 175976
rect 115808 175936 211896 175964
rect 115808 175924 115814 175936
rect 211890 175924 211896 175936
rect 211948 175924 211954 175976
rect 238202 175924 238208 175976
rect 238260 175964 238266 175976
rect 280246 175964 280252 175976
rect 238260 175936 280252 175964
rect 238260 175924 238266 175936
rect 280246 175924 280252 175936
rect 280304 175924 280310 175976
rect 235350 175244 235356 175296
rect 235408 175284 235414 175296
rect 265802 175284 265808 175296
rect 235408 175256 265808 175284
rect 235408 175244 235414 175256
rect 265802 175244 265808 175256
rect 265860 175244 265866 175296
rect 165522 175176 165528 175228
rect 165580 175216 165586 175228
rect 213914 175216 213920 175228
rect 165580 175188 213920 175216
rect 165580 175176 165586 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 231118 175176 231124 175228
rect 231176 175216 231182 175228
rect 250438 175216 250444 175228
rect 231176 175188 250444 175216
rect 231176 175176 231182 175188
rect 250438 175176 250444 175188
rect 250496 175176 250502 175228
rect 231762 175108 231768 175160
rect 231820 175148 231826 175160
rect 245010 175148 245016 175160
rect 231820 175120 245016 175148
rect 231820 175108 231826 175120
rect 245010 175108 245016 175120
rect 245068 175108 245074 175160
rect 165430 174496 165436 174548
rect 165488 174536 165494 174548
rect 214650 174536 214656 174548
rect 165488 174508 214656 174536
rect 165488 174496 165494 174508
rect 214650 174496 214656 174508
rect 214708 174496 214714 174548
rect 256050 174020 256056 174072
rect 256108 174060 256114 174072
rect 265342 174060 265348 174072
rect 256108 174032 265348 174060
rect 256108 174020 256114 174032
rect 265342 174020 265348 174032
rect 265400 174020 265406 174072
rect 247862 173952 247868 174004
rect 247920 173992 247926 174004
rect 265802 173992 265808 174004
rect 247920 173964 265808 173992
rect 247920 173952 247926 173964
rect 265802 173952 265808 173964
rect 265860 173952 265866 174004
rect 238018 173884 238024 173936
rect 238076 173924 238082 173936
rect 265618 173924 265624 173936
rect 238076 173896 265624 173924
rect 238076 173884 238082 173896
rect 265618 173884 265624 173896
rect 265676 173884 265682 173936
rect 166534 173816 166540 173868
rect 166592 173856 166598 173868
rect 213914 173856 213920 173868
rect 166592 173828 213920 173856
rect 166592 173816 166598 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 231210 173816 231216 173868
rect 231268 173856 231274 173868
rect 265250 173856 265256 173868
rect 231268 173828 265256 173856
rect 231268 173816 231274 173828
rect 265250 173816 265256 173828
rect 265308 173816 265314 173868
rect 204898 173748 204904 173800
rect 204956 173788 204962 173800
rect 214006 173788 214012 173800
rect 204956 173760 214012 173788
rect 204956 173748 204962 173760
rect 214006 173748 214012 173760
rect 214064 173748 214070 173800
rect 231762 173748 231768 173800
rect 231820 173788 231826 173800
rect 252002 173788 252008 173800
rect 231820 173760 252008 173788
rect 231820 173748 231826 173760
rect 252002 173748 252008 173760
rect 252060 173748 252066 173800
rect 231670 173680 231676 173732
rect 231728 173720 231734 173732
rect 235994 173720 236000 173732
rect 231728 173692 236000 173720
rect 231728 173680 231734 173692
rect 235994 173680 236000 173692
rect 236052 173680 236058 173732
rect 254670 173136 254676 173188
rect 254728 173176 254734 173188
rect 265894 173176 265900 173188
rect 254728 173148 265900 173176
rect 254728 173136 254734 173148
rect 265894 173136 265900 173148
rect 265952 173136 265958 173188
rect 243630 172592 243636 172644
rect 243688 172632 243694 172644
rect 265894 172632 265900 172644
rect 243688 172604 265900 172632
rect 243688 172592 243694 172604
rect 265894 172592 265900 172604
rect 265952 172592 265958 172644
rect 236822 172524 236828 172576
rect 236880 172564 236886 172576
rect 265802 172564 265808 172576
rect 236880 172536 265808 172564
rect 236880 172524 236886 172536
rect 265802 172524 265808 172536
rect 265860 172524 265866 172576
rect 231762 172456 231768 172508
rect 231820 172496 231826 172508
rect 251266 172496 251272 172508
rect 231820 172468 251272 172496
rect 231820 172456 231826 172468
rect 251266 172456 251272 172468
rect 251324 172456 251330 172508
rect 231670 172388 231676 172440
rect 231728 172428 231734 172440
rect 251358 172428 251364 172440
rect 231728 172400 251364 172428
rect 231728 172388 231734 172400
rect 251358 172388 251364 172400
rect 251416 172388 251422 172440
rect 231670 171708 231676 171760
rect 231728 171748 231734 171760
rect 235258 171748 235264 171760
rect 231728 171720 235264 171748
rect 231728 171708 231734 171720
rect 235258 171708 235264 171720
rect 235316 171708 235322 171760
rect 258810 171504 258816 171556
rect 258868 171544 258874 171556
rect 265342 171544 265348 171556
rect 258868 171516 265348 171544
rect 258868 171504 258874 171516
rect 265342 171504 265348 171516
rect 265400 171504 265406 171556
rect 251818 171164 251824 171216
rect 251876 171204 251882 171216
rect 265894 171204 265900 171216
rect 251876 171176 265900 171204
rect 251876 171164 251882 171176
rect 265894 171164 265900 171176
rect 265952 171164 265958 171216
rect 247678 171096 247684 171148
rect 247736 171136 247742 171148
rect 265802 171136 265808 171148
rect 247736 171108 265808 171136
rect 247736 171096 247742 171108
rect 265802 171096 265808 171108
rect 265860 171096 265866 171148
rect 170582 171028 170588 171080
rect 170640 171068 170646 171080
rect 213914 171068 213920 171080
rect 170640 171040 213920 171068
rect 170640 171028 170646 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 231762 171028 231768 171080
rect 231820 171068 231826 171080
rect 263686 171068 263692 171080
rect 231820 171040 263692 171068
rect 231820 171028 231826 171040
rect 263686 171028 263692 171040
rect 263744 171028 263750 171080
rect 282730 171028 282736 171080
rect 282788 171068 282794 171080
rect 296990 171068 296996 171080
rect 282788 171040 296996 171068
rect 282788 171028 282794 171040
rect 296990 171028 296996 171040
rect 297048 171028 297054 171080
rect 197998 170960 198004 171012
rect 198056 171000 198062 171012
rect 214006 171000 214012 171012
rect 198056 170972 214012 171000
rect 198056 170960 198062 170972
rect 214006 170960 214012 170972
rect 214064 170960 214070 171012
rect 282822 170960 282828 171012
rect 282880 171000 282886 171012
rect 289998 171000 290004 171012
rect 282880 170972 290004 171000
rect 282880 170960 282886 170972
rect 289998 170960 290004 170972
rect 290056 170960 290062 171012
rect 231302 170552 231308 170604
rect 231360 170592 231366 170604
rect 236178 170592 236184 170604
rect 231360 170564 236184 170592
rect 231360 170552 231366 170564
rect 236178 170552 236184 170564
rect 236236 170552 236242 170604
rect 231762 170484 231768 170536
rect 231820 170524 231826 170536
rect 236270 170524 236276 170536
rect 231820 170496 236276 170524
rect 231820 170484 231826 170496
rect 236270 170484 236276 170496
rect 236328 170484 236334 170536
rect 236638 170348 236644 170400
rect 236696 170388 236702 170400
rect 265710 170388 265716 170400
rect 236696 170360 265716 170388
rect 236696 170348 236702 170360
rect 265710 170348 265716 170360
rect 265768 170348 265774 170400
rect 168006 169736 168012 169788
rect 168064 169776 168070 169788
rect 170398 169776 170404 169788
rect 168064 169748 170404 169776
rect 168064 169736 168070 169748
rect 170398 169736 170404 169748
rect 170456 169736 170462 169788
rect 246390 169736 246396 169788
rect 246448 169776 246454 169788
rect 265342 169776 265348 169788
rect 246448 169748 265348 169776
rect 246448 169736 246454 169748
rect 265342 169736 265348 169748
rect 265400 169736 265406 169788
rect 167822 169668 167828 169720
rect 167880 169708 167886 169720
rect 213914 169708 213920 169720
rect 167880 169680 213920 169708
rect 167880 169668 167886 169680
rect 213914 169668 213920 169680
rect 213972 169668 213978 169720
rect 231762 169668 231768 169720
rect 231820 169708 231826 169720
rect 258074 169708 258080 169720
rect 231820 169680 258080 169708
rect 231820 169668 231826 169680
rect 258074 169668 258080 169680
rect 258132 169668 258138 169720
rect 282822 169668 282828 169720
rect 282880 169708 282886 169720
rect 289814 169708 289820 169720
rect 282880 169680 289820 169708
rect 282880 169668 282886 169680
rect 289814 169668 289820 169680
rect 289872 169668 289878 169720
rect 169202 169600 169208 169652
rect 169260 169640 169266 169652
rect 214006 169640 214012 169652
rect 169260 169612 214012 169640
rect 169260 169600 169266 169612
rect 214006 169600 214012 169612
rect 214064 169600 214070 169652
rect 231670 169532 231676 169584
rect 231728 169572 231734 169584
rect 237374 169572 237380 169584
rect 231728 169544 237380 169572
rect 231728 169532 231734 169544
rect 237374 169532 237380 169544
rect 237432 169532 237438 169584
rect 240870 168512 240876 168564
rect 240928 168552 240934 168564
rect 240928 168524 248414 168552
rect 240928 168512 240934 168524
rect 245010 168444 245016 168496
rect 245068 168484 245074 168496
rect 246574 168484 246580 168496
rect 245068 168456 246580 168484
rect 245068 168444 245074 168456
rect 246574 168444 246580 168456
rect 246632 168444 246638 168496
rect 248386 168484 248414 168524
rect 260282 168512 260288 168564
rect 260340 168552 260346 168564
rect 265618 168552 265624 168564
rect 260340 168524 265624 168552
rect 260340 168512 260346 168524
rect 265618 168512 265624 168524
rect 265676 168512 265682 168564
rect 265802 168484 265808 168496
rect 248386 168456 265808 168484
rect 265802 168444 265808 168456
rect 265860 168444 265866 168496
rect 235534 168376 235540 168428
rect 235592 168416 235598 168428
rect 264422 168416 264428 168428
rect 235592 168388 264428 168416
rect 235592 168376 235598 168388
rect 264422 168376 264428 168388
rect 264480 168376 264486 168428
rect 166442 168308 166448 168360
rect 166500 168348 166506 168360
rect 213914 168348 213920 168360
rect 166500 168320 213920 168348
rect 166500 168308 166506 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 231762 168308 231768 168360
rect 231820 168348 231826 168360
rect 260926 168348 260932 168360
rect 231820 168320 260932 168348
rect 231820 168308 231826 168320
rect 260926 168308 260932 168320
rect 260984 168308 260990 168360
rect 282454 168308 282460 168360
rect 282512 168348 282518 168360
rect 292574 168348 292580 168360
rect 282512 168320 292580 168348
rect 282512 168308 282518 168320
rect 292574 168308 292580 168320
rect 292632 168308 292638 168360
rect 180058 168240 180064 168292
rect 180116 168280 180122 168292
rect 214006 168280 214012 168292
rect 180116 168252 214012 168280
rect 180116 168240 180122 168252
rect 214006 168240 214012 168252
rect 214064 168240 214070 168292
rect 231670 168240 231676 168292
rect 231728 168280 231734 168292
rect 254026 168280 254032 168292
rect 231728 168252 254032 168280
rect 231728 168240 231734 168252
rect 254026 168240 254032 168252
rect 254084 168240 254090 168292
rect 231578 168172 231584 168224
rect 231636 168212 231642 168224
rect 250070 168212 250076 168224
rect 231636 168184 250076 168212
rect 231636 168172 231642 168184
rect 250070 168172 250076 168184
rect 250128 168172 250134 168224
rect 246482 167628 246488 167680
rect 246540 167668 246546 167680
rect 265434 167668 265440 167680
rect 246540 167640 265440 167668
rect 246540 167628 246546 167640
rect 265434 167628 265440 167640
rect 265492 167628 265498 167680
rect 262950 167084 262956 167136
rect 263008 167124 263014 167136
rect 265158 167124 265164 167136
rect 263008 167096 265164 167124
rect 263008 167084 263014 167096
rect 265158 167084 265164 167096
rect 265216 167084 265222 167136
rect 239674 167016 239680 167068
rect 239732 167056 239738 167068
rect 265802 167056 265808 167068
rect 239732 167028 265808 167056
rect 239732 167016 239738 167028
rect 265802 167016 265808 167028
rect 265860 167016 265866 167068
rect 231762 166948 231768 167000
rect 231820 166988 231826 167000
rect 244918 166988 244924 167000
rect 231820 166960 244924 166988
rect 231820 166948 231826 166960
rect 244918 166948 244924 166960
rect 244976 166948 244982 167000
rect 282086 166948 282092 167000
rect 282144 166988 282150 167000
rect 294230 166988 294236 167000
rect 282144 166960 294236 166988
rect 282144 166948 282150 166960
rect 294230 166948 294236 166960
rect 294288 166948 294294 167000
rect 382918 166948 382924 167000
rect 382976 166988 382982 167000
rect 580166 166988 580172 167000
rect 382976 166960 580172 166988
rect 382976 166948 382982 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 169294 166880 169300 166932
rect 169352 166920 169358 166932
rect 214006 166920 214012 166932
rect 169352 166892 214012 166920
rect 169352 166880 169358 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 231118 166880 231124 166932
rect 231176 166920 231182 166932
rect 234614 166920 234620 166932
rect 231176 166892 234620 166920
rect 231176 166880 231182 166892
rect 234614 166880 234620 166892
rect 234672 166880 234678 166932
rect 166350 166812 166356 166864
rect 166408 166852 166414 166864
rect 213914 166852 213920 166864
rect 166408 166824 213920 166852
rect 166408 166812 166414 166824
rect 213914 166812 213920 166824
rect 213972 166812 213978 166864
rect 240778 166268 240784 166320
rect 240836 166308 240842 166320
rect 265342 166308 265348 166320
rect 240836 166280 265348 166308
rect 240836 166268 240842 166280
rect 265342 166268 265348 166280
rect 265400 166268 265406 166320
rect 231486 166064 231492 166116
rect 231544 166104 231550 166116
rect 236086 166104 236092 166116
rect 231544 166076 236092 166104
rect 231544 166064 231550 166076
rect 236086 166064 236092 166076
rect 236144 166064 236150 166116
rect 261478 165656 261484 165708
rect 261536 165696 261542 165708
rect 265802 165696 265808 165708
rect 261536 165668 265808 165696
rect 261536 165656 261542 165668
rect 265802 165656 265808 165668
rect 265860 165656 265866 165708
rect 245102 165588 245108 165640
rect 245160 165628 245166 165640
rect 265710 165628 265716 165640
rect 245160 165600 265716 165628
rect 245160 165588 245166 165600
rect 265710 165588 265716 165600
rect 265768 165588 265774 165640
rect 178678 165520 178684 165572
rect 178736 165560 178742 165572
rect 213914 165560 213920 165572
rect 178736 165532 213920 165560
rect 178736 165520 178742 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 231762 165520 231768 165572
rect 231820 165560 231826 165572
rect 255406 165560 255412 165572
rect 231820 165532 255412 165560
rect 231820 165520 231826 165532
rect 255406 165520 255412 165532
rect 255464 165520 255470 165572
rect 281994 165520 282000 165572
rect 282052 165560 282058 165572
rect 294138 165560 294144 165572
rect 282052 165532 294144 165560
rect 282052 165520 282058 165532
rect 294138 165520 294144 165532
rect 294196 165520 294202 165572
rect 211890 165452 211896 165504
rect 211948 165492 211954 165504
rect 214650 165492 214656 165504
rect 211948 165464 214656 165492
rect 211948 165452 211954 165464
rect 214650 165452 214656 165464
rect 214708 165452 214714 165504
rect 231302 165452 231308 165504
rect 231360 165492 231366 165504
rect 234706 165492 234712 165504
rect 231360 165464 234712 165492
rect 231360 165452 231366 165464
rect 234706 165452 234712 165464
rect 234764 165452 234770 165504
rect 282822 165452 282828 165504
rect 282880 165492 282886 165504
rect 291470 165492 291476 165504
rect 282880 165464 291476 165492
rect 282880 165452 282886 165464
rect 291470 165452 291476 165464
rect 291528 165452 291534 165504
rect 236914 164840 236920 164892
rect 236972 164880 236978 164892
rect 261386 164880 261392 164892
rect 236972 164852 261392 164880
rect 236972 164840 236978 164852
rect 261386 164840 261392 164852
rect 261444 164840 261450 164892
rect 230658 164568 230664 164620
rect 230716 164608 230722 164620
rect 232130 164608 232136 164620
rect 230716 164580 232136 164608
rect 230716 164568 230722 164580
rect 232130 164568 232136 164580
rect 232188 164568 232194 164620
rect 257430 164296 257436 164348
rect 257488 164336 257494 164348
rect 265802 164336 265808 164348
rect 257488 164308 265808 164336
rect 257488 164296 257494 164308
rect 265802 164296 265808 164308
rect 265860 164296 265866 164348
rect 242250 164228 242256 164280
rect 242308 164268 242314 164280
rect 265434 164268 265440 164280
rect 242308 164240 265440 164268
rect 242308 164228 242314 164240
rect 265434 164228 265440 164240
rect 265492 164228 265498 164280
rect 177298 164160 177304 164212
rect 177356 164200 177362 164212
rect 213914 164200 213920 164212
rect 177356 164172 213920 164200
rect 177356 164160 177362 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 231670 164160 231676 164212
rect 231728 164200 231734 164212
rect 242158 164200 242164 164212
rect 231728 164172 242164 164200
rect 231728 164160 231734 164172
rect 242158 164160 242164 164172
rect 242216 164160 242222 164212
rect 282822 164160 282828 164212
rect 282880 164200 282886 164212
rect 295518 164200 295524 164212
rect 282880 164172 295524 164200
rect 282880 164160 282886 164172
rect 295518 164160 295524 164172
rect 295576 164160 295582 164212
rect 211798 164092 211804 164144
rect 211856 164132 211862 164144
rect 214466 164132 214472 164144
rect 211856 164104 214472 164132
rect 211856 164092 211862 164104
rect 214466 164092 214472 164104
rect 214524 164092 214530 164144
rect 282086 163208 282092 163260
rect 282144 163248 282150 163260
rect 288618 163248 288624 163260
rect 282144 163220 288624 163248
rect 282144 163208 282150 163220
rect 288618 163208 288624 163220
rect 288676 163208 288682 163260
rect 250622 163004 250628 163056
rect 250680 163044 250686 163056
rect 265526 163044 265532 163056
rect 250680 163016 265532 163044
rect 250680 163004 250686 163016
rect 265526 163004 265532 163016
rect 265584 163004 265590 163056
rect 242342 162936 242348 162988
rect 242400 162976 242406 162988
rect 265342 162976 265348 162988
rect 242400 162948 265348 162976
rect 242400 162936 242406 162948
rect 265342 162936 265348 162948
rect 265400 162936 265406 162988
rect 235258 162868 235264 162920
rect 235316 162908 235322 162920
rect 265894 162908 265900 162920
rect 235316 162880 265900 162908
rect 235316 162868 235322 162880
rect 265894 162868 265900 162880
rect 265952 162868 265958 162920
rect 169110 162800 169116 162852
rect 169168 162840 169174 162852
rect 213914 162840 213920 162852
rect 169168 162812 213920 162840
rect 169168 162800 169174 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 231762 162800 231768 162852
rect 231820 162840 231826 162852
rect 249978 162840 249984 162852
rect 231820 162812 249984 162840
rect 231820 162800 231826 162812
rect 249978 162800 249984 162812
rect 250036 162800 250042 162852
rect 282086 162800 282092 162852
rect 282144 162840 282150 162852
rect 298094 162840 298100 162852
rect 282144 162812 298100 162840
rect 282144 162800 282150 162812
rect 298094 162800 298100 162812
rect 298152 162800 298158 162852
rect 231670 162732 231676 162784
rect 231728 162772 231734 162784
rect 238846 162772 238852 162784
rect 231728 162744 238852 162772
rect 231728 162732 231734 162744
rect 238846 162732 238852 162744
rect 238904 162732 238910 162784
rect 282822 162732 282828 162784
rect 282880 162772 282886 162784
rect 292850 162772 292856 162784
rect 282880 162744 292856 162772
rect 282880 162732 282886 162744
rect 292850 162732 292856 162744
rect 292908 162732 292914 162784
rect 260190 162120 260196 162172
rect 260248 162160 260254 162172
rect 265802 162160 265808 162172
rect 260248 162132 265808 162160
rect 260248 162120 260254 162132
rect 265802 162120 265808 162132
rect 265860 162120 265866 162172
rect 231762 161984 231768 162036
rect 231820 162024 231826 162036
rect 237558 162024 237564 162036
rect 231820 161996 237564 162024
rect 231820 161984 231826 161996
rect 237558 161984 237564 161996
rect 237616 161984 237622 162036
rect 249518 161508 249524 161560
rect 249576 161548 249582 161560
rect 265342 161548 265348 161560
rect 249576 161520 265348 161548
rect 249576 161508 249582 161520
rect 265342 161508 265348 161520
rect 265400 161508 265406 161560
rect 238294 161440 238300 161492
rect 238352 161480 238358 161492
rect 265802 161480 265808 161492
rect 238352 161452 265808 161480
rect 238352 161440 238358 161452
rect 265802 161440 265808 161452
rect 265860 161440 265866 161492
rect 169018 161372 169024 161424
rect 169076 161412 169082 161424
rect 213914 161412 213920 161424
rect 169076 161384 213920 161412
rect 169076 161372 169082 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 231762 161372 231768 161424
rect 231820 161412 231826 161424
rect 262306 161412 262312 161424
rect 231820 161384 262312 161412
rect 231820 161372 231826 161384
rect 262306 161372 262312 161384
rect 262364 161372 262370 161424
rect 282822 161372 282828 161424
rect 282880 161412 282886 161424
rect 291194 161412 291200 161424
rect 282880 161384 291200 161412
rect 282880 161372 282886 161384
rect 291194 161372 291200 161384
rect 291252 161372 291258 161424
rect 231394 161304 231400 161356
rect 231452 161344 231458 161356
rect 245010 161344 245016 161356
rect 231452 161316 245016 161344
rect 231452 161304 231458 161316
rect 245010 161304 245016 161316
rect 245068 161304 245074 161356
rect 167730 160692 167736 160744
rect 167788 160732 167794 160744
rect 214098 160732 214104 160744
rect 167788 160704 214104 160732
rect 167788 160692 167794 160704
rect 214098 160692 214104 160704
rect 214156 160692 214162 160744
rect 281534 160624 281540 160676
rect 281592 160664 281598 160676
rect 283190 160664 283196 160676
rect 281592 160636 283196 160664
rect 281592 160624 281598 160636
rect 283190 160624 283196 160636
rect 283248 160624 283254 160676
rect 255958 160216 255964 160268
rect 256016 160256 256022 160268
rect 265618 160256 265624 160268
rect 256016 160228 265624 160256
rect 256016 160216 256022 160228
rect 265618 160216 265624 160228
rect 265676 160216 265682 160268
rect 244918 160148 244924 160200
rect 244976 160188 244982 160200
rect 265342 160188 265348 160200
rect 244976 160160 265348 160188
rect 244976 160148 244982 160160
rect 265342 160148 265348 160160
rect 265400 160148 265406 160200
rect 239490 160080 239496 160132
rect 239548 160120 239554 160132
rect 265802 160120 265808 160132
rect 239548 160092 265808 160120
rect 239548 160080 239554 160092
rect 265802 160080 265808 160092
rect 265860 160080 265866 160132
rect 167638 160012 167644 160064
rect 167696 160052 167702 160064
rect 213914 160052 213920 160064
rect 167696 160024 213920 160052
rect 167696 160012 167702 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 231486 160012 231492 160064
rect 231544 160052 231550 160064
rect 249242 160052 249248 160064
rect 231544 160024 249248 160052
rect 231544 160012 231550 160024
rect 249242 160012 249248 160024
rect 249300 160012 249306 160064
rect 281534 160012 281540 160064
rect 281592 160052 281598 160064
rect 284478 160052 284484 160064
rect 281592 160024 284484 160052
rect 281592 160012 281598 160024
rect 284478 160012 284484 160024
rect 284536 160012 284542 160064
rect 170490 159944 170496 159996
rect 170548 159984 170554 159996
rect 214006 159984 214012 159996
rect 170548 159956 214012 159984
rect 170548 159944 170554 159956
rect 214006 159944 214012 159956
rect 214064 159944 214070 159996
rect 231762 159944 231768 159996
rect 231820 159984 231826 159996
rect 240226 159984 240232 159996
rect 231820 159956 240232 159984
rect 231820 159944 231826 159956
rect 240226 159944 240232 159956
rect 240284 159944 240290 159996
rect 263042 158856 263048 158908
rect 263100 158896 263106 158908
rect 265618 158896 265624 158908
rect 263100 158868 265624 158896
rect 263100 158856 263106 158868
rect 265618 158856 265624 158868
rect 265676 158856 265682 158908
rect 249426 158788 249432 158840
rect 249484 158828 249490 158840
rect 265342 158828 265348 158840
rect 249484 158800 265348 158828
rect 249484 158788 249490 158800
rect 265342 158788 265348 158800
rect 265400 158788 265406 158840
rect 242158 158720 242164 158772
rect 242216 158760 242222 158772
rect 265802 158760 265808 158772
rect 242216 158732 265808 158760
rect 242216 158720 242222 158732
rect 265802 158720 265808 158732
rect 265860 158720 265866 158772
rect 166258 158652 166264 158704
rect 166316 158692 166322 158704
rect 213914 158692 213920 158704
rect 166316 158664 213920 158692
rect 166316 158652 166322 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 231762 158652 231768 158704
rect 231820 158692 231826 158704
rect 260834 158692 260840 158704
rect 231820 158664 260840 158692
rect 231820 158652 231826 158664
rect 260834 158652 260840 158664
rect 260892 158652 260898 158704
rect 282730 158652 282736 158704
rect 282788 158692 282794 158704
rect 295610 158692 295616 158704
rect 282788 158664 295616 158692
rect 282788 158652 282794 158664
rect 295610 158652 295616 158664
rect 295668 158652 295674 158704
rect 282822 158584 282828 158636
rect 282880 158624 282886 158636
rect 288710 158624 288716 158636
rect 282880 158596 288716 158624
rect 282880 158584 282886 158596
rect 288710 158584 288716 158596
rect 288768 158584 288774 158636
rect 254762 157972 254768 158024
rect 254820 158012 254826 158024
rect 265986 158012 265992 158024
rect 254820 157984 265992 158012
rect 254820 157972 254826 157984
rect 265986 157972 265992 157984
rect 266044 157972 266050 158024
rect 236730 157428 236736 157480
rect 236788 157468 236794 157480
rect 265618 157468 265624 157480
rect 236788 157440 265624 157468
rect 236788 157428 236794 157440
rect 265618 157428 265624 157440
rect 265676 157428 265682 157480
rect 232498 157360 232504 157412
rect 232556 157400 232562 157412
rect 265526 157400 265532 157412
rect 232556 157372 265532 157400
rect 232556 157360 232562 157372
rect 265526 157360 265532 157372
rect 265584 157360 265590 157412
rect 209038 157292 209044 157344
rect 209096 157332 209102 157344
rect 213914 157332 213920 157344
rect 209096 157304 213920 157332
rect 209096 157292 209102 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 231762 157292 231768 157344
rect 231820 157332 231826 157344
rect 259546 157332 259552 157344
rect 231820 157304 259552 157332
rect 231820 157292 231826 157304
rect 259546 157292 259552 157304
rect 259604 157292 259610 157344
rect 231670 157224 231676 157276
rect 231728 157264 231734 157276
rect 256786 157264 256792 157276
rect 231728 157236 256792 157264
rect 231728 157224 231734 157236
rect 256786 157224 256792 157236
rect 256844 157224 256850 157276
rect 281718 156544 281724 156596
rect 281776 156584 281782 156596
rect 284570 156584 284576 156596
rect 281776 156556 284576 156584
rect 281776 156544 281782 156556
rect 284570 156544 284576 156556
rect 284628 156544 284634 156596
rect 253198 156068 253204 156120
rect 253256 156108 253262 156120
rect 265894 156108 265900 156120
rect 253256 156080 265900 156108
rect 253256 156068 253262 156080
rect 265894 156068 265900 156080
rect 265952 156068 265958 156120
rect 246666 156000 246672 156052
rect 246724 156040 246730 156052
rect 265526 156040 265532 156052
rect 246724 156012 265532 156040
rect 246724 156000 246730 156012
rect 265526 156000 265532 156012
rect 265584 156000 265590 156052
rect 238202 155932 238208 155984
rect 238260 155972 238266 155984
rect 265802 155972 265808 155984
rect 238260 155944 265808 155972
rect 238260 155932 238266 155944
rect 265802 155932 265808 155944
rect 265860 155932 265866 155984
rect 173158 155864 173164 155916
rect 173216 155904 173222 155916
rect 213914 155904 213920 155916
rect 173216 155876 213920 155904
rect 173216 155864 173222 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 231118 155796 231124 155848
rect 231176 155836 231182 155848
rect 233234 155836 233240 155848
rect 231176 155808 233240 155836
rect 231176 155796 231182 155808
rect 233234 155796 233240 155808
rect 233292 155796 233298 155848
rect 231762 155728 231768 155780
rect 231820 155768 231826 155780
rect 246298 155768 246304 155780
rect 231820 155740 246304 155768
rect 231820 155728 231826 155740
rect 246298 155728 246304 155740
rect 246356 155728 246362 155780
rect 258902 155524 258908 155576
rect 258960 155564 258966 155576
rect 261662 155564 261668 155576
rect 258960 155536 261668 155564
rect 258960 155524 258966 155536
rect 261662 155524 261668 155536
rect 261720 155524 261726 155576
rect 230566 155388 230572 155440
rect 230624 155428 230630 155440
rect 232038 155428 232044 155440
rect 230624 155400 232044 155428
rect 230624 155388 230630 155400
rect 232038 155388 232044 155400
rect 232096 155388 232102 155440
rect 250714 154640 250720 154692
rect 250772 154680 250778 154692
rect 265802 154680 265808 154692
rect 250772 154652 265808 154680
rect 250772 154640 250778 154652
rect 265802 154640 265808 154652
rect 265860 154640 265866 154692
rect 239582 154572 239588 154624
rect 239640 154612 239646 154624
rect 265710 154612 265716 154624
rect 239640 154584 265716 154612
rect 239640 154572 239646 154584
rect 265710 154572 265716 154584
rect 265768 154572 265774 154624
rect 281718 154504 281724 154556
rect 281776 154544 281782 154556
rect 300946 154544 300952 154556
rect 281776 154516 300952 154544
rect 281776 154504 281782 154516
rect 300946 154504 300952 154516
rect 301004 154504 301010 154556
rect 252186 153824 252192 153876
rect 252244 153864 252250 153876
rect 265250 153864 265256 153876
rect 252244 153836 265256 153864
rect 252244 153824 252250 153836
rect 265250 153824 265256 153836
rect 265308 153824 265314 153876
rect 282822 153416 282828 153468
rect 282880 153456 282886 153468
rect 287238 153456 287244 153468
rect 282880 153428 287244 153456
rect 282880 153416 282886 153428
rect 287238 153416 287244 153428
rect 287296 153416 287302 153468
rect 180058 153280 180064 153332
rect 180116 153320 180122 153332
rect 213914 153320 213920 153332
rect 180116 153292 213920 153320
rect 180116 153280 180122 153292
rect 213914 153280 213920 153292
rect 213972 153280 213978 153332
rect 241146 153280 241152 153332
rect 241204 153320 241210 153332
rect 265894 153320 265900 153332
rect 241204 153292 265900 153320
rect 241204 153280 241210 153292
rect 265894 153280 265900 153292
rect 265952 153280 265958 153332
rect 169018 153212 169024 153264
rect 169076 153252 169082 153264
rect 214006 153252 214012 153264
rect 169076 153224 214012 153252
rect 169076 153212 169082 153224
rect 214006 153212 214012 153224
rect 214064 153212 214070 153264
rect 234154 153212 234160 153264
rect 234212 153252 234218 153264
rect 265802 153252 265808 153264
rect 234212 153224 265808 153252
rect 234212 153212 234218 153224
rect 265802 153212 265808 153224
rect 265860 153212 265866 153264
rect 231762 153144 231768 153196
rect 231820 153184 231826 153196
rect 262214 153184 262220 153196
rect 231820 153156 262220 153184
rect 231820 153144 231826 153156
rect 262214 153144 262220 153156
rect 262272 153144 262278 153196
rect 282730 153144 282736 153196
rect 282788 153184 282794 153196
rect 304994 153184 305000 153196
rect 282788 153156 305000 153184
rect 282788 153144 282794 153156
rect 304994 153144 305000 153156
rect 305052 153144 305058 153196
rect 381538 153144 381544 153196
rect 381596 153184 381602 153196
rect 579798 153184 579804 153196
rect 381596 153156 579804 153184
rect 381596 153144 381602 153156
rect 579798 153144 579804 153156
rect 579856 153144 579862 153196
rect 231670 153076 231676 153128
rect 231728 153116 231734 153128
rect 244366 153116 244372 153128
rect 231728 153088 244372 153116
rect 231728 153076 231734 153088
rect 244366 153076 244372 153088
rect 244424 153076 244430 153128
rect 234522 152464 234528 152516
rect 234580 152504 234586 152516
rect 242066 152504 242072 152516
rect 234580 152476 242072 152504
rect 234580 152464 234586 152476
rect 242066 152464 242072 152476
rect 242124 152464 242130 152516
rect 245194 152464 245200 152516
rect 245252 152504 245258 152516
rect 265986 152504 265992 152516
rect 245252 152476 265992 152504
rect 245252 152464 245258 152476
rect 265986 152464 265992 152476
rect 266044 152464 266050 152516
rect 241054 151920 241060 151972
rect 241112 151960 241118 151972
rect 265710 151960 265716 151972
rect 241112 151932 265716 151960
rect 241112 151920 241118 151932
rect 265710 151920 265716 151932
rect 265768 151920 265774 151972
rect 196618 151852 196624 151904
rect 196676 151892 196682 151904
rect 213914 151892 213920 151904
rect 196676 151864 213920 151892
rect 196676 151852 196682 151864
rect 213914 151852 213920 151864
rect 213972 151852 213978 151904
rect 177390 151784 177396 151836
rect 177448 151824 177454 151836
rect 214006 151824 214012 151836
rect 177448 151796 214012 151824
rect 177448 151784 177454 151796
rect 214006 151784 214012 151796
rect 214064 151784 214070 151836
rect 261754 151784 261760 151836
rect 261812 151824 261818 151836
rect 265802 151824 265808 151836
rect 261812 151796 265808 151824
rect 261812 151784 261818 151796
rect 265802 151784 265808 151796
rect 265860 151784 265866 151836
rect 282822 151716 282828 151768
rect 282880 151756 282886 151768
rect 301130 151756 301136 151768
rect 282880 151728 301136 151756
rect 282880 151716 282886 151728
rect 301130 151716 301136 151728
rect 301188 151716 301194 151768
rect 231670 151648 231676 151700
rect 231728 151688 231734 151700
rect 234522 151688 234528 151700
rect 231728 151660 234528 151688
rect 231728 151648 231734 151660
rect 234522 151648 234528 151660
rect 234580 151648 234586 151700
rect 231762 151580 231768 151632
rect 231820 151620 231826 151632
rect 238754 151620 238760 151632
rect 231820 151592 238760 151620
rect 231820 151580 231826 151592
rect 238754 151580 238760 151592
rect 238812 151580 238818 151632
rect 258718 150560 258724 150612
rect 258776 150600 258782 150612
rect 265894 150600 265900 150612
rect 258776 150572 265900 150600
rect 258776 150560 258782 150572
rect 265894 150560 265900 150572
rect 265952 150560 265958 150612
rect 198090 150492 198096 150544
rect 198148 150532 198154 150544
rect 213914 150532 213920 150544
rect 198148 150504 213920 150532
rect 198148 150492 198154 150504
rect 213914 150492 213920 150504
rect 213972 150492 213978 150544
rect 254854 150492 254860 150544
rect 254912 150532 254918 150544
rect 265986 150532 265992 150544
rect 254912 150504 265992 150532
rect 254912 150492 254918 150504
rect 265986 150492 265992 150504
rect 266044 150492 266050 150544
rect 170490 150424 170496 150476
rect 170548 150464 170554 150476
rect 214006 150464 214012 150476
rect 170548 150436 214012 150464
rect 170548 150424 170554 150436
rect 214006 150424 214012 150436
rect 214064 150424 214070 150476
rect 246574 150424 246580 150476
rect 246632 150464 246638 150476
rect 265802 150464 265808 150476
rect 246632 150436 265808 150464
rect 246632 150424 246638 150436
rect 265802 150424 265808 150436
rect 265860 150424 265866 150476
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 11698 150396 11704 150408
rect 3476 150368 11704 150396
rect 3476 150356 3482 150368
rect 11698 150356 11704 150368
rect 11756 150356 11762 150408
rect 170398 150356 170404 150408
rect 170456 150396 170462 150408
rect 213914 150396 213920 150408
rect 170456 150368 213920 150396
rect 170456 150356 170462 150368
rect 213914 150356 213920 150368
rect 213972 150356 213978 150408
rect 282822 150356 282828 150408
rect 282880 150396 282886 150408
rect 291378 150396 291384 150408
rect 282880 150368 291384 150396
rect 282880 150356 282886 150368
rect 291378 150356 291384 150368
rect 291436 150356 291442 150408
rect 231670 150288 231676 150340
rect 231728 150328 231734 150340
rect 249058 150328 249064 150340
rect 231728 150300 249064 150328
rect 231728 150288 231734 150300
rect 249058 150288 249064 150300
rect 249116 150288 249122 150340
rect 231762 150220 231768 150272
rect 231820 150260 231826 150272
rect 253934 150260 253940 150272
rect 231820 150232 253940 150260
rect 231820 150220 231826 150232
rect 253934 150220 253940 150232
rect 253992 150220 253998 150272
rect 230934 150016 230940 150068
rect 230992 150056 230998 150068
rect 233418 150056 233424 150068
rect 230992 150028 233424 150056
rect 230992 150016 230998 150028
rect 233418 150016 233424 150028
rect 233476 150016 233482 150068
rect 231210 149676 231216 149728
rect 231268 149716 231274 149728
rect 245102 149716 245108 149728
rect 231268 149688 245108 149716
rect 231268 149676 231274 149688
rect 245102 149676 245108 149688
rect 245160 149676 245166 149728
rect 281534 149608 281540 149660
rect 281592 149648 281598 149660
rect 284294 149648 284300 149660
rect 281592 149620 284300 149648
rect 281592 149608 281598 149620
rect 284294 149608 284300 149620
rect 284352 149608 284358 149660
rect 263134 149200 263140 149252
rect 263192 149240 263198 149252
rect 265342 149240 265348 149252
rect 263192 149212 265348 149240
rect 263192 149200 263198 149212
rect 265342 149200 265348 149212
rect 265400 149200 265406 149252
rect 249334 149132 249340 149184
rect 249392 149172 249398 149184
rect 265802 149172 265808 149184
rect 249392 149144 265808 149172
rect 249392 149132 249398 149144
rect 265802 149132 265808 149144
rect 265860 149132 265866 149184
rect 245010 149064 245016 149116
rect 245068 149104 245074 149116
rect 265894 149104 265900 149116
rect 245068 149076 265900 149104
rect 245068 149064 245074 149076
rect 265894 149064 265900 149076
rect 265952 149064 265958 149116
rect 231762 148996 231768 149048
rect 231820 149036 231826 149048
rect 243538 149036 243544 149048
rect 231820 149008 243544 149036
rect 231820 148996 231826 149008
rect 243538 148996 243544 149008
rect 243596 148996 243602 149048
rect 282822 148996 282828 149048
rect 282880 149036 282886 149048
rect 290090 149036 290096 149048
rect 282880 149008 290096 149036
rect 282880 148996 282886 149008
rect 290090 148996 290096 149008
rect 290148 148996 290154 149048
rect 282270 148588 282276 148640
rect 282328 148628 282334 148640
rect 287330 148628 287336 148640
rect 282328 148600 287336 148628
rect 282328 148588 282334 148600
rect 287330 148588 287336 148600
rect 287388 148588 287394 148640
rect 232774 148316 232780 148368
rect 232832 148356 232838 148368
rect 266078 148356 266084 148368
rect 232832 148328 266084 148356
rect 232832 148316 232838 148328
rect 266078 148316 266084 148328
rect 266136 148316 266142 148368
rect 258994 147704 259000 147756
rect 259052 147744 259058 147756
rect 265802 147744 265808 147756
rect 259052 147716 265808 147744
rect 259052 147704 259058 147716
rect 265802 147704 265808 147716
rect 265860 147704 265866 147756
rect 166258 147636 166264 147688
rect 166316 147676 166322 147688
rect 213914 147676 213920 147688
rect 166316 147648 213920 147676
rect 166316 147636 166322 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 235442 147636 235448 147688
rect 235500 147676 235506 147688
rect 265434 147676 265440 147688
rect 235500 147648 265440 147676
rect 235500 147636 235506 147648
rect 265434 147636 265440 147648
rect 265492 147636 265498 147688
rect 231762 147568 231768 147620
rect 231820 147608 231826 147620
rect 263594 147608 263600 147620
rect 231820 147580 263600 147608
rect 231820 147568 231826 147580
rect 263594 147568 263600 147580
rect 263652 147568 263658 147620
rect 281718 147568 281724 147620
rect 281776 147608 281782 147620
rect 316034 147608 316040 147620
rect 281776 147580 316040 147608
rect 281776 147568 281782 147580
rect 316034 147568 316040 147580
rect 316092 147568 316098 147620
rect 230934 147024 230940 147076
rect 230992 147064 230998 147076
rect 233326 147064 233332 147076
rect 230992 147036 233332 147064
rect 230992 147024 230998 147036
rect 233326 147024 233332 147036
rect 233384 147024 233390 147076
rect 232590 146888 232596 146940
rect 232648 146928 232654 146940
rect 265158 146928 265164 146940
rect 232648 146900 265164 146928
rect 232648 146888 232654 146900
rect 265158 146888 265164 146900
rect 265216 146888 265222 146940
rect 234062 146344 234068 146396
rect 234120 146384 234126 146396
rect 265802 146384 265808 146396
rect 234120 146356 265808 146384
rect 234120 146344 234126 146356
rect 265802 146344 265808 146356
rect 265860 146344 265866 146396
rect 174538 146276 174544 146328
rect 174596 146316 174602 146328
rect 213914 146316 213920 146328
rect 174596 146288 213920 146316
rect 174596 146276 174602 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 232682 146276 232688 146328
rect 232740 146316 232746 146328
rect 265526 146316 265532 146328
rect 232740 146288 265532 146316
rect 232740 146276 232746 146288
rect 265526 146276 265532 146288
rect 265584 146276 265590 146328
rect 231762 146208 231768 146260
rect 231820 146248 231826 146260
rect 244274 146248 244280 146260
rect 231820 146220 244280 146248
rect 231820 146208 231826 146220
rect 244274 146208 244280 146220
rect 244332 146208 244338 146260
rect 281994 146208 282000 146260
rect 282052 146248 282058 146260
rect 299750 146248 299756 146260
rect 282052 146220 299756 146248
rect 282052 146208 282058 146220
rect 299750 146208 299756 146220
rect 299808 146208 299814 146260
rect 231670 146140 231676 146192
rect 231728 146180 231734 146192
rect 242986 146180 242992 146192
rect 231728 146152 242992 146180
rect 231728 146140 231734 146152
rect 242986 146140 242992 146152
rect 243044 146140 243050 146192
rect 282822 146140 282828 146192
rect 282880 146180 282886 146192
rect 296714 146180 296720 146192
rect 282880 146152 296720 146180
rect 282880 146140 282886 146152
rect 296714 146140 296720 146152
rect 296772 146140 296778 146192
rect 231026 146072 231032 146124
rect 231084 146112 231090 146124
rect 237466 146112 237472 146124
rect 231084 146084 237472 146112
rect 231084 146072 231090 146084
rect 237466 146072 237472 146084
rect 237524 146072 237530 146124
rect 238386 145528 238392 145580
rect 238444 145568 238450 145580
rect 261570 145568 261576 145580
rect 238444 145540 261576 145568
rect 238444 145528 238450 145540
rect 261570 145528 261576 145540
rect 261628 145528 261634 145580
rect 233970 145052 233976 145104
rect 234028 145092 234034 145104
rect 265802 145092 265808 145104
rect 234028 145064 265808 145092
rect 234028 145052 234034 145064
rect 265802 145052 265808 145064
rect 265860 145052 265866 145104
rect 252094 144984 252100 145036
rect 252152 145024 252158 145036
rect 265526 145024 265532 145036
rect 252152 144996 265532 145024
rect 252152 144984 252158 144996
rect 265526 144984 265532 144996
rect 265584 144984 265590 145036
rect 178678 144916 178684 144968
rect 178736 144956 178742 144968
rect 213914 144956 213920 144968
rect 178736 144928 213920 144956
rect 178736 144916 178742 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 231578 144848 231584 144900
rect 231636 144888 231642 144900
rect 231636 144860 258074 144888
rect 231636 144848 231642 144860
rect 258046 144820 258074 144860
rect 261846 144848 261852 144900
rect 261904 144888 261910 144900
rect 265710 144888 265716 144900
rect 261904 144860 265716 144888
rect 261904 144848 261910 144860
rect 265710 144848 265716 144860
rect 265768 144848 265774 144900
rect 263778 144820 263784 144832
rect 258046 144792 263784 144820
rect 263778 144780 263784 144792
rect 263836 144780 263842 144832
rect 282546 144780 282552 144832
rect 282604 144820 282610 144832
rect 285766 144820 285772 144832
rect 282604 144792 285772 144820
rect 282604 144780 282610 144792
rect 285766 144780 285772 144792
rect 285824 144780 285830 144832
rect 282822 143692 282828 143744
rect 282880 143732 282886 143744
rect 287054 143732 287060 143744
rect 282880 143704 287060 143732
rect 282880 143692 282886 143704
rect 287054 143692 287060 143704
rect 287112 143692 287118 143744
rect 177298 143624 177304 143676
rect 177356 143664 177362 143676
rect 214006 143664 214012 143676
rect 177356 143636 214012 143664
rect 177356 143624 177362 143636
rect 214006 143624 214012 143636
rect 214064 143624 214070 143676
rect 250806 143624 250812 143676
rect 250864 143664 250870 143676
rect 265434 143664 265440 143676
rect 250864 143636 265440 143664
rect 250864 143624 250870 143636
rect 265434 143624 265440 143636
rect 265492 143624 265498 143676
rect 171870 143556 171876 143608
rect 171928 143596 171934 143608
rect 213914 143596 213920 143608
rect 171928 143568 213920 143596
rect 171928 143556 171934 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 229922 143556 229928 143608
rect 229980 143596 229986 143608
rect 265802 143596 265808 143608
rect 229980 143568 265808 143596
rect 229980 143556 229986 143568
rect 265802 143556 265808 143568
rect 265860 143556 265866 143608
rect 231670 143488 231676 143540
rect 231728 143528 231734 143540
rect 259454 143528 259460 143540
rect 231728 143500 259460 143528
rect 231728 143488 231734 143500
rect 259454 143488 259460 143500
rect 259512 143488 259518 143540
rect 281626 143488 281632 143540
rect 281684 143528 281690 143540
rect 301038 143528 301044 143540
rect 281684 143500 301044 143528
rect 281684 143488 281690 143500
rect 301038 143488 301044 143500
rect 301096 143488 301102 143540
rect 231762 143420 231768 143472
rect 231820 143460 231826 143472
rect 251174 143460 251180 143472
rect 231820 143432 251180 143460
rect 231820 143420 231826 143432
rect 251174 143420 251180 143432
rect 251232 143420 251238 143472
rect 231118 143352 231124 143404
rect 231176 143392 231182 143404
rect 233786 143392 233792 143404
rect 231176 143364 233792 143392
rect 231176 143352 231182 143364
rect 233786 143352 233792 143364
rect 233844 143352 233850 143404
rect 233878 142808 233884 142860
rect 233936 142848 233942 142860
rect 265618 142848 265624 142860
rect 233936 142820 265624 142848
rect 233936 142808 233942 142820
rect 265618 142808 265624 142820
rect 265676 142808 265682 142860
rect 260374 142332 260380 142384
rect 260432 142372 260438 142384
rect 264330 142372 264336 142384
rect 260432 142344 264336 142372
rect 260432 142332 260438 142344
rect 264330 142332 264336 142344
rect 264388 142332 264394 142384
rect 243722 142264 243728 142316
rect 243780 142304 243786 142316
rect 265342 142304 265348 142316
rect 243780 142276 265348 142304
rect 243780 142264 243786 142276
rect 265342 142264 265348 142276
rect 265400 142264 265406 142316
rect 188338 142128 188344 142180
rect 188396 142168 188402 142180
rect 213914 142168 213920 142180
rect 188396 142140 213920 142168
rect 188396 142128 188402 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 231762 142060 231768 142112
rect 231820 142100 231826 142112
rect 255590 142100 255596 142112
rect 231820 142072 255596 142100
rect 231820 142060 231826 142072
rect 255590 142060 255596 142072
rect 255648 142060 255654 142112
rect 282822 142060 282828 142112
rect 282880 142100 282886 142112
rect 303706 142100 303712 142112
rect 282880 142072 303712 142100
rect 282880 142060 282886 142072
rect 303706 142060 303712 142072
rect 303764 142060 303770 142112
rect 231302 141448 231308 141500
rect 231360 141488 231366 141500
rect 251818 141488 251824 141500
rect 231360 141460 251824 141488
rect 231360 141448 231366 141460
rect 251818 141448 251824 141460
rect 251876 141448 251882 141500
rect 245286 141380 245292 141432
rect 245344 141420 245350 141432
rect 266078 141420 266084 141432
rect 245344 141392 266084 141420
rect 245344 141380 245350 141392
rect 266078 141380 266084 141392
rect 266136 141380 266142 141432
rect 175918 140836 175924 140888
rect 175976 140876 175982 140888
rect 213914 140876 213920 140888
rect 175976 140848 213920 140876
rect 175976 140836 175982 140848
rect 213914 140836 213920 140848
rect 213972 140836 213978 140888
rect 170398 140768 170404 140820
rect 170456 140808 170462 140820
rect 214006 140808 214012 140820
rect 170456 140780 214012 140808
rect 170456 140768 170462 140780
rect 214006 140768 214012 140780
rect 214064 140768 214070 140820
rect 256326 140768 256332 140820
rect 256384 140808 256390 140820
rect 265802 140808 265808 140820
rect 256384 140780 265808 140808
rect 256384 140768 256390 140780
rect 265802 140768 265808 140780
rect 265860 140768 265866 140820
rect 231670 140700 231676 140752
rect 231728 140740 231734 140752
rect 256694 140740 256700 140752
rect 231728 140712 256700 140740
rect 231728 140700 231734 140712
rect 256694 140700 256700 140712
rect 256752 140700 256758 140752
rect 281902 140700 281908 140752
rect 281960 140740 281966 140752
rect 296806 140740 296812 140752
rect 281960 140712 296812 140740
rect 281960 140700 281966 140712
rect 296806 140700 296812 140712
rect 296864 140700 296870 140752
rect 231762 140632 231768 140684
rect 231820 140672 231826 140684
rect 247034 140672 247040 140684
rect 231820 140644 247040 140672
rect 231820 140632 231826 140644
rect 247034 140632 247040 140644
rect 247092 140632 247098 140684
rect 210418 139408 210424 139460
rect 210476 139448 210482 139460
rect 213914 139448 213920 139460
rect 210476 139420 213920 139448
rect 210476 139408 210482 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 257338 139408 257344 139460
rect 257396 139448 257402 139460
rect 265434 139448 265440 139460
rect 257396 139420 265440 139448
rect 257396 139408 257402 139420
rect 265434 139408 265440 139420
rect 265492 139408 265498 139460
rect 282822 139340 282828 139392
rect 282880 139380 282886 139392
rect 313274 139380 313280 139392
rect 282880 139352 313280 139380
rect 282880 139340 282886 139352
rect 313274 139340 313280 139352
rect 313332 139340 313338 139392
rect 282730 139272 282736 139324
rect 282788 139312 282794 139324
rect 292758 139312 292764 139324
rect 282788 139284 292764 139312
rect 282788 139272 282794 139284
rect 292758 139272 292764 139284
rect 292816 139272 292822 139324
rect 231210 138660 231216 138712
rect 231268 138700 231274 138712
rect 244918 138700 244924 138712
rect 231268 138672 244924 138700
rect 231268 138660 231274 138672
rect 244918 138660 244924 138672
rect 244976 138660 244982 138712
rect 247770 138116 247776 138168
rect 247828 138156 247834 138168
rect 265618 138156 265624 138168
rect 247828 138128 265624 138156
rect 247828 138116 247834 138128
rect 265618 138116 265624 138128
rect 265676 138116 265682 138168
rect 202138 138048 202144 138100
rect 202196 138088 202202 138100
rect 213914 138088 213920 138100
rect 202196 138060 213920 138088
rect 202196 138048 202202 138060
rect 213914 138048 213920 138060
rect 213972 138048 213978 138100
rect 243538 138048 243544 138100
rect 243596 138088 243602 138100
rect 265158 138088 265164 138100
rect 243596 138060 265164 138088
rect 243596 138048 243602 138060
rect 265158 138048 265164 138060
rect 265216 138048 265222 138100
rect 171962 137980 171968 138032
rect 172020 138020 172026 138032
rect 214006 138020 214012 138032
rect 172020 137992 214012 138020
rect 172020 137980 172026 137992
rect 214006 137980 214012 137992
rect 214064 137980 214070 138032
rect 229738 137980 229744 138032
rect 229796 138020 229802 138032
rect 265434 138020 265440 138032
rect 229796 137992 265440 138020
rect 229796 137980 229802 137992
rect 265434 137980 265440 137992
rect 265492 137980 265498 138032
rect 3418 137912 3424 137964
rect 3476 137952 3482 137964
rect 14458 137952 14464 137964
rect 3476 137924 14464 137952
rect 3476 137912 3482 137924
rect 14458 137912 14464 137924
rect 14516 137912 14522 137964
rect 231394 137912 231400 137964
rect 231452 137952 231458 137964
rect 262398 137952 262404 137964
rect 231452 137924 262404 137952
rect 231452 137912 231458 137924
rect 262398 137912 262404 137924
rect 262456 137912 262462 137964
rect 282178 137912 282184 137964
rect 282236 137952 282242 137964
rect 298370 137952 298376 137964
rect 282236 137924 298376 137952
rect 282236 137912 282242 137924
rect 298370 137912 298376 137924
rect 298428 137912 298434 137964
rect 231762 137844 231768 137896
rect 231820 137884 231826 137896
rect 242894 137884 242900 137896
rect 231820 137856 242900 137884
rect 231820 137844 231826 137856
rect 242894 137844 242900 137856
rect 242952 137844 242958 137896
rect 282822 137844 282828 137896
rect 282880 137884 282886 137896
rect 293954 137884 293960 137896
rect 282880 137856 293960 137884
rect 282880 137844 282886 137856
rect 293954 137844 293960 137856
rect 294012 137844 294018 137896
rect 231578 137232 231584 137284
rect 231636 137272 231642 137284
rect 243630 137272 243636 137284
rect 231636 137244 243636 137272
rect 231636 137232 231642 137244
rect 243630 137232 243636 137244
rect 243688 137232 243694 137284
rect 249242 136688 249248 136740
rect 249300 136728 249306 136740
rect 265526 136728 265532 136740
rect 249300 136700 265532 136728
rect 249300 136688 249306 136700
rect 265526 136688 265532 136700
rect 265584 136688 265590 136740
rect 206370 136620 206376 136672
rect 206428 136660 206434 136672
rect 213914 136660 213920 136672
rect 206428 136632 213920 136660
rect 206428 136620 206434 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 239398 136620 239404 136672
rect 239456 136660 239462 136672
rect 265618 136660 265624 136672
rect 239456 136632 265624 136660
rect 239456 136620 239462 136632
rect 265618 136620 265624 136632
rect 265676 136620 265682 136672
rect 231394 136552 231400 136604
rect 231452 136592 231458 136604
rect 256050 136592 256056 136604
rect 231452 136564 256056 136592
rect 231452 136552 231458 136564
rect 256050 136552 256056 136564
rect 256108 136552 256114 136604
rect 231762 136484 231768 136536
rect 231820 136524 231826 136536
rect 247862 136524 247868 136536
rect 231820 136496 247868 136524
rect 231820 136484 231826 136496
rect 247862 136484 247868 136496
rect 247920 136484 247926 136536
rect 260098 135464 260104 135516
rect 260156 135504 260162 135516
rect 265342 135504 265348 135516
rect 260156 135476 265348 135504
rect 260156 135464 260162 135476
rect 265342 135464 265348 135476
rect 265400 135464 265406 135516
rect 261478 135396 261484 135448
rect 261536 135436 261542 135448
rect 266078 135436 266084 135448
rect 261536 135408 266084 135436
rect 261536 135396 261542 135408
rect 266078 135396 266084 135408
rect 266136 135396 266142 135448
rect 253382 135328 253388 135380
rect 253440 135368 253446 135380
rect 265618 135368 265624 135380
rect 253440 135340 265624 135368
rect 253440 135328 253446 135340
rect 265618 135328 265624 135340
rect 265676 135328 265682 135380
rect 238110 135260 238116 135312
rect 238168 135300 238174 135312
rect 265894 135300 265900 135312
rect 238168 135272 265900 135300
rect 238168 135260 238174 135272
rect 265894 135260 265900 135272
rect 265952 135260 265958 135312
rect 231486 135192 231492 135244
rect 231544 135232 231550 135244
rect 254670 135232 254676 135244
rect 231544 135204 254676 135232
rect 231544 135192 231550 135204
rect 254670 135192 254676 135204
rect 254728 135192 254734 135244
rect 231026 135056 231032 135108
rect 231084 135096 231090 135108
rect 236638 135096 236644 135108
rect 231084 135068 236644 135096
rect 231084 135056 231090 135068
rect 236638 135056 236644 135068
rect 236696 135056 236702 135108
rect 173342 134512 173348 134564
rect 173400 134552 173406 134564
rect 214834 134552 214840 134564
rect 173400 134524 214840 134552
rect 173400 134512 173406 134524
rect 214834 134512 214840 134524
rect 214892 134512 214898 134564
rect 254578 134036 254584 134088
rect 254636 134076 254642 134088
rect 265894 134076 265900 134088
rect 254636 134048 265900 134076
rect 254636 134036 254642 134048
rect 265894 134036 265900 134048
rect 265952 134036 265958 134088
rect 253290 133968 253296 134020
rect 253348 134008 253354 134020
rect 265526 134008 265532 134020
rect 253348 133980 265532 134008
rect 253348 133968 253354 133980
rect 265526 133968 265532 133980
rect 265584 133968 265590 134020
rect 204898 133900 204904 133952
rect 204956 133940 204962 133952
rect 213914 133940 213920 133952
rect 204956 133912 213920 133940
rect 204956 133900 204962 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 229830 133900 229836 133952
rect 229888 133940 229894 133952
rect 265894 133940 265900 133952
rect 229888 133912 265900 133940
rect 229888 133900 229894 133912
rect 265894 133900 265900 133912
rect 265952 133900 265958 133952
rect 231670 133832 231676 133884
rect 231728 133872 231734 133884
rect 258810 133872 258816 133884
rect 231728 133844 258816 133872
rect 231728 133832 231734 133844
rect 258810 133832 258816 133844
rect 258868 133832 258874 133884
rect 282822 133832 282828 133884
rect 282880 133872 282886 133884
rect 311894 133872 311900 133884
rect 282880 133844 311900 133872
rect 282880 133832 282886 133844
rect 311894 133832 311900 133844
rect 311952 133832 311958 133884
rect 230934 133764 230940 133816
rect 230992 133804 230998 133816
rect 236822 133804 236828 133816
rect 230992 133776 236828 133804
rect 230992 133764 230998 133776
rect 236822 133764 236828 133776
rect 236880 133764 236886 133816
rect 262858 132608 262864 132660
rect 262916 132648 262922 132660
rect 265618 132648 265624 132660
rect 262916 132620 265624 132648
rect 262916 132608 262922 132620
rect 265618 132608 265624 132620
rect 265676 132608 265682 132660
rect 184198 132540 184204 132592
rect 184256 132580 184262 132592
rect 213914 132580 213920 132592
rect 184256 132552 213920 132580
rect 184256 132540 184262 132552
rect 213914 132540 213920 132552
rect 213972 132540 213978 132592
rect 171778 132472 171784 132524
rect 171836 132512 171842 132524
rect 214006 132512 214012 132524
rect 171836 132484 214012 132512
rect 171836 132472 171842 132484
rect 214006 132472 214012 132484
rect 214064 132472 214070 132524
rect 236638 132472 236644 132524
rect 236696 132512 236702 132524
rect 265894 132512 265900 132524
rect 236696 132484 265900 132512
rect 236696 132472 236702 132484
rect 265894 132472 265900 132484
rect 265952 132472 265958 132524
rect 231762 132404 231768 132456
rect 231820 132444 231826 132456
rect 247678 132444 247684 132456
rect 231820 132416 247684 132444
rect 231820 132404 231826 132416
rect 247678 132404 247684 132416
rect 247736 132404 247742 132456
rect 282822 132404 282828 132456
rect 282880 132444 282886 132456
rect 307754 132444 307760 132456
rect 282880 132416 307760 132444
rect 282880 132404 282886 132416
rect 307754 132404 307760 132416
rect 307812 132404 307818 132456
rect 231670 132336 231676 132388
rect 231728 132376 231734 132388
rect 246390 132376 246396 132388
rect 231728 132348 246396 132376
rect 231728 132336 231734 132348
rect 246390 132336 246396 132348
rect 246448 132336 246454 132388
rect 250438 131248 250444 131300
rect 250496 131288 250502 131300
rect 265158 131288 265164 131300
rect 250496 131260 265164 131288
rect 250496 131248 250502 131260
rect 265158 131248 265164 131260
rect 265216 131248 265222 131300
rect 206278 131180 206284 131232
rect 206336 131220 206342 131232
rect 213914 131220 213920 131232
rect 206336 131192 213920 131220
rect 206336 131180 206342 131192
rect 213914 131180 213920 131192
rect 213972 131180 213978 131232
rect 247862 131180 247868 131232
rect 247920 131220 247926 131232
rect 265618 131220 265624 131232
rect 247920 131192 265624 131220
rect 247920 131180 247926 131192
rect 265618 131180 265624 131192
rect 265676 131180 265682 131232
rect 186958 131112 186964 131164
rect 187016 131152 187022 131164
rect 214006 131152 214012 131164
rect 187016 131124 214012 131152
rect 187016 131112 187022 131124
rect 214006 131112 214012 131124
rect 214064 131112 214070 131164
rect 231486 131112 231492 131164
rect 231544 131152 231550 131164
rect 235534 131152 235540 131164
rect 231544 131124 235540 131152
rect 231544 131112 231550 131124
rect 235534 131112 235540 131124
rect 235592 131112 235598 131164
rect 246298 131112 246304 131164
rect 246356 131152 246362 131164
rect 265894 131152 265900 131164
rect 246356 131124 265900 131152
rect 246356 131112 246362 131124
rect 265894 131112 265900 131124
rect 265952 131112 265958 131164
rect 231762 131044 231768 131096
rect 231820 131084 231826 131096
rect 264238 131084 264244 131096
rect 231820 131056 264244 131084
rect 231820 131044 231826 131056
rect 264238 131044 264244 131056
rect 264296 131044 264302 131096
rect 282822 131044 282828 131096
rect 282880 131084 282886 131096
rect 302326 131084 302332 131096
rect 282880 131056 302332 131084
rect 282880 131044 282886 131056
rect 302326 131044 302332 131056
rect 302384 131044 302390 131096
rect 231394 130976 231400 131028
rect 231452 131016 231458 131028
rect 260282 131016 260288 131028
rect 231452 130988 260288 131016
rect 231452 130976 231458 130988
rect 260282 130976 260288 130988
rect 260340 130976 260346 131028
rect 231670 130908 231676 130960
rect 231728 130948 231734 130960
rect 246482 130948 246488 130960
rect 231728 130920 246488 130948
rect 231728 130908 231734 130920
rect 246482 130908 246488 130920
rect 246540 130908 246546 130960
rect 282270 130568 282276 130620
rect 282328 130608 282334 130620
rect 285858 130608 285864 130620
rect 282328 130580 285864 130608
rect 282328 130568 282334 130580
rect 285858 130568 285864 130580
rect 285916 130568 285922 130620
rect 176010 129820 176016 129872
rect 176068 129860 176074 129872
rect 214006 129860 214012 129872
rect 176068 129832 214012 129860
rect 176068 129820 176074 129832
rect 214006 129820 214012 129832
rect 214064 129820 214070 129872
rect 174630 129752 174636 129804
rect 174688 129792 174694 129804
rect 213914 129792 213920 129804
rect 174688 129764 213920 129792
rect 174688 129752 174694 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 231302 129684 231308 129736
rect 231360 129724 231366 129736
rect 240778 129724 240784 129736
rect 231360 129696 240784 129724
rect 231360 129684 231366 129696
rect 240778 129684 240784 129696
rect 240836 129684 240842 129736
rect 231578 129004 231584 129056
rect 231636 129044 231642 129056
rect 257430 129044 257436 129056
rect 231636 129016 257436 129044
rect 231636 129004 231642 129016
rect 257430 129004 257436 129016
rect 257488 129004 257494 129056
rect 282822 128460 282828 128512
rect 282880 128500 282886 128512
rect 287146 128500 287152 128512
rect 282880 128472 287152 128500
rect 282880 128460 282886 128472
rect 287146 128460 287152 128472
rect 287204 128460 287210 128512
rect 257522 128392 257528 128444
rect 257580 128432 257586 128444
rect 265618 128432 265624 128444
rect 257580 128404 265624 128432
rect 257580 128392 257586 128404
rect 265618 128392 265624 128404
rect 265676 128392 265682 128444
rect 177482 128324 177488 128376
rect 177540 128364 177546 128376
rect 213914 128364 213920 128376
rect 177540 128336 213920 128364
rect 177540 128324 177546 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 244918 128324 244924 128376
rect 244976 128364 244982 128376
rect 265894 128364 265900 128376
rect 244976 128336 265900 128364
rect 244976 128324 244982 128336
rect 265894 128324 265900 128336
rect 265952 128324 265958 128376
rect 231670 128256 231676 128308
rect 231728 128296 231734 128308
rect 262950 128296 262956 128308
rect 231728 128268 262956 128296
rect 231728 128256 231734 128268
rect 262950 128256 262956 128268
rect 263008 128256 263014 128308
rect 281718 128256 281724 128308
rect 281776 128296 281782 128308
rect 303798 128296 303804 128308
rect 281776 128268 303804 128296
rect 281776 128256 281782 128268
rect 303798 128256 303804 128268
rect 303856 128256 303862 128308
rect 231762 128188 231768 128240
rect 231820 128228 231826 128240
rect 240870 128228 240876 128240
rect 231820 128200 240876 128228
rect 231820 128188 231826 128200
rect 240870 128188 240876 128200
rect 240928 128188 240934 128240
rect 231670 127780 231676 127832
rect 231728 127820 231734 127832
rect 236914 127820 236920 127832
rect 231728 127792 236920 127820
rect 231728 127780 231734 127792
rect 236914 127780 236920 127792
rect 236972 127780 236978 127832
rect 252002 127032 252008 127084
rect 252060 127072 252066 127084
rect 265894 127072 265900 127084
rect 252060 127044 265900 127072
rect 252060 127032 252066 127044
rect 265894 127032 265900 127044
rect 265952 127032 265958 127084
rect 174722 126964 174728 127016
rect 174780 127004 174786 127016
rect 213914 127004 213920 127016
rect 174780 126976 213920 127004
rect 174780 126964 174786 126976
rect 213914 126964 213920 126976
rect 213972 126964 213978 127016
rect 240778 126964 240784 127016
rect 240836 127004 240842 127016
rect 265342 127004 265348 127016
rect 240836 126976 265348 127004
rect 240836 126964 240842 126976
rect 265342 126964 265348 126976
rect 265400 126964 265406 127016
rect 231118 126896 231124 126948
rect 231176 126936 231182 126948
rect 254762 126936 254768 126948
rect 231176 126908 254768 126936
rect 231176 126896 231182 126908
rect 254762 126896 254768 126908
rect 254820 126896 254826 126948
rect 305638 126896 305644 126948
rect 305696 126936 305702 126948
rect 580166 126936 580172 126948
rect 305696 126908 580172 126936
rect 305696 126896 305702 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 231762 126828 231768 126880
rect 231820 126868 231826 126880
rect 239674 126868 239680 126880
rect 231820 126840 239680 126868
rect 231820 126828 231826 126840
rect 239674 126828 239680 126840
rect 239732 126828 239738 126880
rect 231486 126216 231492 126268
rect 231544 126256 231550 126268
rect 242342 126256 242348 126268
rect 231544 126228 242348 126256
rect 231544 126216 231550 126228
rect 242342 126216 242348 126228
rect 242400 126216 242406 126268
rect 242526 126216 242532 126268
rect 242584 126256 242590 126268
rect 265986 126256 265992 126268
rect 242584 126228 265992 126256
rect 242584 126216 242590 126228
rect 265986 126216 265992 126228
rect 266044 126216 266050 126268
rect 188430 125672 188436 125724
rect 188488 125712 188494 125724
rect 214006 125712 214012 125724
rect 188488 125684 214012 125712
rect 188488 125672 188494 125684
rect 214006 125672 214012 125684
rect 214064 125672 214070 125724
rect 257614 125672 257620 125724
rect 257672 125712 257678 125724
rect 265250 125712 265256 125724
rect 257672 125684 265256 125712
rect 257672 125672 257678 125684
rect 265250 125672 265256 125684
rect 265308 125672 265314 125724
rect 63402 125604 63408 125656
rect 63460 125644 63466 125656
rect 65150 125644 65156 125656
rect 63460 125616 65156 125644
rect 63460 125604 63466 125616
rect 65150 125604 65156 125616
rect 65208 125604 65214 125656
rect 167638 125604 167644 125656
rect 167696 125644 167702 125656
rect 213914 125644 213920 125656
rect 167696 125616 213920 125644
rect 167696 125604 167702 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 247678 125604 247684 125656
rect 247736 125644 247742 125656
rect 265894 125644 265900 125656
rect 247736 125616 265900 125644
rect 247736 125604 247742 125616
rect 265894 125604 265900 125616
rect 265952 125604 265958 125656
rect 231762 125536 231768 125588
rect 231820 125576 231826 125588
rect 242250 125576 242256 125588
rect 231820 125548 242256 125576
rect 231820 125536 231826 125548
rect 242250 125536 242256 125548
rect 242308 125536 242314 125588
rect 282086 125536 282092 125588
rect 282144 125576 282150 125588
rect 285674 125576 285680 125588
rect 282144 125548 285680 125576
rect 282144 125536 282150 125548
rect 285674 125536 285680 125548
rect 285732 125536 285738 125588
rect 231302 124924 231308 124976
rect 231360 124964 231366 124976
rect 233878 124964 233884 124976
rect 231360 124936 233884 124964
rect 231360 124924 231366 124936
rect 233878 124924 233884 124936
rect 233936 124924 233942 124976
rect 230842 124856 230848 124908
rect 230900 124896 230906 124908
rect 249518 124896 249524 124908
rect 230900 124868 249524 124896
rect 230900 124856 230906 124868
rect 249518 124856 249524 124868
rect 249576 124856 249582 124908
rect 282822 124652 282828 124704
rect 282880 124692 282886 124704
rect 288526 124692 288532 124704
rect 282880 124664 288532 124692
rect 282880 124652 282886 124664
rect 288526 124652 288532 124664
rect 288584 124652 288590 124704
rect 251910 124312 251916 124364
rect 251968 124352 251974 124364
rect 265986 124352 265992 124364
rect 251968 124324 265992 124352
rect 251968 124312 251974 124324
rect 265986 124312 265992 124324
rect 266044 124312 266050 124364
rect 199378 124244 199384 124296
rect 199436 124284 199442 124296
rect 213914 124284 213920 124296
rect 199436 124256 213920 124284
rect 199436 124244 199442 124256
rect 213914 124244 213920 124256
rect 213972 124244 213978 124296
rect 249150 124244 249156 124296
rect 249208 124284 249214 124296
rect 265526 124284 265532 124296
rect 249208 124256 265532 124284
rect 249208 124244 249214 124256
rect 265526 124244 265532 124256
rect 265584 124244 265590 124296
rect 167730 124176 167736 124228
rect 167788 124216 167794 124228
rect 214006 124216 214012 124228
rect 167788 124188 214012 124216
rect 167788 124176 167794 124188
rect 214006 124176 214012 124188
rect 214064 124176 214070 124228
rect 240870 124176 240876 124228
rect 240928 124216 240934 124228
rect 265894 124216 265900 124228
rect 240928 124188 265900 124216
rect 240928 124176 240934 124188
rect 265894 124176 265900 124188
rect 265952 124176 265958 124228
rect 231762 124108 231768 124160
rect 231820 124148 231826 124160
rect 250622 124148 250628 124160
rect 231820 124120 250628 124148
rect 231820 124108 231826 124120
rect 250622 124108 250628 124120
rect 250680 124108 250686 124160
rect 282730 124108 282736 124160
rect 282788 124148 282794 124160
rect 300854 124148 300860 124160
rect 282788 124120 300860 124148
rect 282788 124108 282794 124120
rect 300854 124108 300860 124120
rect 300912 124108 300918 124160
rect 282822 124040 282828 124092
rect 282880 124080 282886 124092
rect 295334 124080 295340 124092
rect 282880 124052 295340 124080
rect 282880 124040 282886 124052
rect 295334 124040 295340 124052
rect 295392 124040 295398 124092
rect 231578 123564 231584 123616
rect 231636 123604 231642 123616
rect 235258 123604 235264 123616
rect 231636 123576 235264 123604
rect 231636 123564 231642 123576
rect 235258 123564 235264 123576
rect 235316 123564 235322 123616
rect 230750 123496 230756 123548
rect 230808 123536 230814 123548
rect 253198 123536 253204 123548
rect 230808 123508 253204 123536
rect 230808 123496 230814 123508
rect 253198 123496 253204 123508
rect 253256 123496 253262 123548
rect 242250 123428 242256 123480
rect 242308 123468 242314 123480
rect 265710 123468 265716 123480
rect 242308 123440 265716 123468
rect 242308 123428 242314 123440
rect 265710 123428 265716 123440
rect 265768 123428 265774 123480
rect 250530 122952 250536 123004
rect 250588 122992 250594 123004
rect 265066 122992 265072 123004
rect 250588 122964 265072 122992
rect 250588 122952 250594 122964
rect 265066 122952 265072 122964
rect 265124 122952 265130 123004
rect 170582 122884 170588 122936
rect 170640 122924 170646 122936
rect 213914 122924 213920 122936
rect 170640 122896 213920 122924
rect 170640 122884 170646 122896
rect 213914 122884 213920 122896
rect 213972 122884 213978 122936
rect 254670 122884 254676 122936
rect 254728 122924 254734 122936
rect 265526 122924 265532 122936
rect 254728 122896 265532 122924
rect 254728 122884 254734 122896
rect 265526 122884 265532 122896
rect 265584 122884 265590 122936
rect 166350 122816 166356 122868
rect 166408 122856 166414 122868
rect 214006 122856 214012 122868
rect 166408 122828 214012 122856
rect 166408 122816 166414 122828
rect 214006 122816 214012 122828
rect 214064 122816 214070 122868
rect 231302 122748 231308 122800
rect 231360 122788 231366 122800
rect 260190 122788 260196 122800
rect 231360 122760 260196 122788
rect 231360 122748 231366 122760
rect 260190 122748 260196 122760
rect 260248 122748 260254 122800
rect 282086 122748 282092 122800
rect 282144 122788 282150 122800
rect 309134 122788 309140 122800
rect 282144 122760 309140 122788
rect 282144 122748 282150 122760
rect 309134 122748 309140 122760
rect 309192 122748 309198 122800
rect 167914 122068 167920 122120
rect 167972 122108 167978 122120
rect 198090 122108 198096 122120
rect 167972 122080 198096 122108
rect 167972 122068 167978 122080
rect 198090 122068 198096 122080
rect 198148 122068 198154 122120
rect 231670 122068 231676 122120
rect 231728 122108 231734 122120
rect 250714 122108 250720 122120
rect 231728 122080 250720 122108
rect 231728 122068 231734 122080
rect 250714 122068 250720 122080
rect 250772 122068 250778 122120
rect 211798 121524 211804 121576
rect 211856 121564 211862 121576
rect 214466 121564 214472 121576
rect 211856 121536 214472 121564
rect 211856 121524 211862 121536
rect 214466 121524 214472 121536
rect 214524 121524 214530 121576
rect 253198 121524 253204 121576
rect 253256 121564 253262 121576
rect 265986 121564 265992 121576
rect 253256 121536 265992 121564
rect 253256 121524 253262 121536
rect 265986 121524 265992 121536
rect 266044 121524 266050 121576
rect 197998 121456 198004 121508
rect 198056 121496 198062 121508
rect 213914 121496 213920 121508
rect 198056 121468 213920 121496
rect 198056 121456 198062 121468
rect 213914 121456 213920 121468
rect 213972 121456 213978 121508
rect 233878 121456 233884 121508
rect 233936 121496 233942 121508
rect 265894 121496 265900 121508
rect 233936 121468 265900 121496
rect 233936 121456 233942 121468
rect 265894 121456 265900 121468
rect 265952 121456 265958 121508
rect 231762 121388 231768 121440
rect 231820 121428 231826 121440
rect 258902 121428 258908 121440
rect 231820 121400 258908 121428
rect 231820 121388 231826 121400
rect 258902 121388 258908 121400
rect 258960 121388 258966 121440
rect 282454 121388 282460 121440
rect 282512 121428 282518 121440
rect 302234 121428 302240 121440
rect 282512 121400 302240 121428
rect 282512 121388 282518 121400
rect 302234 121388 302240 121400
rect 302292 121388 302298 121440
rect 230934 121320 230940 121372
rect 230992 121360 230998 121372
rect 238294 121360 238300 121372
rect 230992 121332 238300 121360
rect 230992 121320 230998 121332
rect 238294 121320 238300 121332
rect 238352 121320 238358 121372
rect 281718 121320 281724 121372
rect 281776 121360 281782 121372
rect 291286 121360 291292 121372
rect 281776 121332 291292 121360
rect 281776 121320 281782 121332
rect 291286 121320 291292 121332
rect 291344 121320 291350 121372
rect 231210 120708 231216 120760
rect 231268 120748 231274 120760
rect 264514 120748 264520 120760
rect 231268 120720 264520 120748
rect 231268 120708 231274 120720
rect 264514 120708 264520 120720
rect 264572 120708 264578 120760
rect 178770 120164 178776 120216
rect 178828 120204 178834 120216
rect 213914 120204 213920 120216
rect 178828 120176 213920 120204
rect 178828 120164 178834 120176
rect 213914 120164 213920 120176
rect 213972 120164 213978 120216
rect 258810 120164 258816 120216
rect 258868 120204 258874 120216
rect 265986 120204 265992 120216
rect 258868 120176 265992 120204
rect 258868 120164 258874 120176
rect 265986 120164 265992 120176
rect 266044 120164 266050 120216
rect 170674 120096 170680 120148
rect 170732 120136 170738 120148
rect 214006 120136 214012 120148
rect 170732 120108 214012 120136
rect 170732 120096 170738 120108
rect 214006 120096 214012 120108
rect 214064 120096 214070 120148
rect 238018 120096 238024 120148
rect 238076 120136 238082 120148
rect 265894 120136 265900 120148
rect 238076 120108 265900 120136
rect 238076 120096 238082 120108
rect 265894 120096 265900 120108
rect 265952 120096 265958 120148
rect 230934 120028 230940 120080
rect 230992 120068 230998 120080
rect 255958 120068 255964 120080
rect 230992 120040 255964 120068
rect 230992 120028 230998 120040
rect 255958 120028 255964 120040
rect 256016 120028 256022 120080
rect 282086 120028 282092 120080
rect 282144 120068 282150 120080
rect 298186 120068 298192 120080
rect 282144 120040 298192 120068
rect 282144 120028 282150 120040
rect 298186 120028 298192 120040
rect 298244 120028 298250 120080
rect 231486 119960 231492 120012
rect 231544 120000 231550 120012
rect 249426 120000 249432 120012
rect 231544 119972 249432 120000
rect 231544 119960 231550 119972
rect 249426 119960 249432 119972
rect 249484 119960 249490 120012
rect 231762 119892 231768 119944
rect 231820 119932 231826 119944
rect 239490 119932 239496 119944
rect 231820 119904 239496 119932
rect 231820 119892 231826 119904
rect 239490 119892 239496 119904
rect 239548 119892 239554 119944
rect 169110 118804 169116 118856
rect 169168 118844 169174 118856
rect 214006 118844 214012 118856
rect 169168 118816 214012 118844
rect 169168 118804 169174 118816
rect 214006 118804 214012 118816
rect 214064 118804 214070 118856
rect 173434 118736 173440 118788
rect 173492 118776 173498 118788
rect 213914 118776 213920 118788
rect 173492 118748 213920 118776
rect 173492 118736 173498 118748
rect 213914 118736 213920 118748
rect 213972 118736 213978 118788
rect 256142 118736 256148 118788
rect 256200 118776 256206 118788
rect 265250 118776 265256 118788
rect 256200 118748 265256 118776
rect 256200 118736 256206 118748
rect 265250 118736 265256 118748
rect 265308 118736 265314 118788
rect 254762 118668 254768 118720
rect 254820 118708 254826 118720
rect 265710 118708 265716 118720
rect 254820 118680 265716 118708
rect 254820 118668 254826 118680
rect 265710 118668 265716 118680
rect 265768 118668 265774 118720
rect 230658 118600 230664 118652
rect 230716 118640 230722 118652
rect 263042 118640 263048 118652
rect 230716 118612 263048 118640
rect 230716 118600 230722 118612
rect 263042 118600 263048 118612
rect 263100 118600 263106 118652
rect 282822 118600 282828 118652
rect 282880 118640 282886 118652
rect 292666 118640 292672 118652
rect 282880 118612 292672 118640
rect 282880 118600 282886 118612
rect 292666 118600 292672 118612
rect 292724 118600 292730 118652
rect 231762 118532 231768 118584
rect 231820 118572 231826 118584
rect 242158 118572 242164 118584
rect 231820 118544 242164 118572
rect 231820 118532 231826 118544
rect 242158 118532 242164 118544
rect 242216 118532 242222 118584
rect 282730 118532 282736 118584
rect 282788 118572 282794 118584
rect 289906 118572 289912 118584
rect 282788 118544 289912 118572
rect 282788 118532 282794 118544
rect 289906 118532 289912 118544
rect 289964 118532 289970 118584
rect 230934 117512 230940 117564
rect 230992 117552 230998 117564
rect 236730 117552 236736 117564
rect 230992 117524 236736 117552
rect 230992 117512 230998 117524
rect 236730 117512 236736 117524
rect 236788 117512 236794 117564
rect 262950 117444 262956 117496
rect 263008 117484 263014 117496
rect 265158 117484 265164 117496
rect 263008 117456 265164 117484
rect 263008 117444 263014 117456
rect 265158 117444 265164 117456
rect 265216 117444 265222 117496
rect 191190 117376 191196 117428
rect 191248 117416 191254 117428
rect 214006 117416 214012 117428
rect 191248 117388 214012 117416
rect 191248 117376 191254 117388
rect 214006 117376 214012 117388
rect 214064 117376 214070 117428
rect 257430 117376 257436 117428
rect 257488 117416 257494 117428
rect 265526 117416 265532 117428
rect 257488 117388 265532 117416
rect 257488 117376 257494 117388
rect 265526 117376 265532 117388
rect 265584 117376 265590 117428
rect 169202 117308 169208 117360
rect 169260 117348 169266 117360
rect 213914 117348 213920 117360
rect 169260 117320 213920 117348
rect 169260 117308 169266 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 239490 117308 239496 117360
rect 239548 117348 239554 117360
rect 265710 117348 265716 117360
rect 239548 117320 265716 117348
rect 239548 117308 239554 117320
rect 265710 117308 265716 117320
rect 265768 117308 265774 117360
rect 230658 117240 230664 117292
rect 230716 117280 230722 117292
rect 252186 117280 252192 117292
rect 230716 117252 252192 117280
rect 230716 117240 230722 117252
rect 252186 117240 252192 117252
rect 252244 117240 252250 117292
rect 282822 117240 282828 117292
rect 282880 117280 282886 117292
rect 306466 117280 306472 117292
rect 282880 117252 306472 117280
rect 282880 117240 282886 117252
rect 306466 117240 306472 117252
rect 306524 117240 306530 117292
rect 282730 117172 282736 117224
rect 282788 117212 282794 117224
rect 295426 117212 295432 117224
rect 282788 117184 295432 117212
rect 282788 117172 282794 117184
rect 295426 117172 295432 117184
rect 295484 117172 295490 117224
rect 231210 116560 231216 116612
rect 231268 116600 231274 116612
rect 250806 116600 250812 116612
rect 231268 116572 250812 116600
rect 231268 116560 231274 116572
rect 250806 116560 250812 116572
rect 250864 116560 250870 116612
rect 230566 116492 230572 116544
rect 230624 116532 230630 116544
rect 232498 116532 232504 116544
rect 230624 116504 232504 116532
rect 230624 116492 230630 116504
rect 232498 116492 232504 116504
rect 232556 116492 232562 116544
rect 256234 116084 256240 116136
rect 256292 116124 256298 116136
rect 264514 116124 264520 116136
rect 256292 116096 264520 116124
rect 256292 116084 256298 116096
rect 264514 116084 264520 116096
rect 264572 116084 264578 116136
rect 251818 116016 251824 116068
rect 251876 116056 251882 116068
rect 266078 116056 266084 116068
rect 251876 116028 266084 116056
rect 251876 116016 251882 116028
rect 266078 116016 266084 116028
rect 266136 116016 266142 116068
rect 180150 115948 180156 116000
rect 180208 115988 180214 116000
rect 213914 115988 213920 116000
rect 180208 115960 213920 115988
rect 180208 115948 180214 115960
rect 213914 115948 213920 115960
rect 213972 115948 213978 116000
rect 246390 115948 246396 116000
rect 246448 115988 246454 116000
rect 266170 115988 266176 116000
rect 246448 115960 266176 115988
rect 246448 115948 246454 115960
rect 266170 115948 266176 115960
rect 266228 115948 266234 116000
rect 231762 115880 231768 115932
rect 231820 115920 231826 115932
rect 246666 115920 246672 115932
rect 231820 115892 246672 115920
rect 231820 115880 231826 115892
rect 246666 115880 246672 115892
rect 246724 115880 246730 115932
rect 281718 115880 281724 115932
rect 281776 115920 281782 115932
rect 303614 115920 303620 115932
rect 281776 115892 303620 115920
rect 281776 115880 281782 115892
rect 303614 115880 303620 115892
rect 303672 115880 303678 115932
rect 282086 115812 282092 115864
rect 282144 115852 282150 115864
rect 296898 115852 296904 115864
rect 282144 115824 296904 115852
rect 282144 115812 282150 115824
rect 296898 115812 296904 115824
rect 296956 115812 296962 115864
rect 231578 115200 231584 115252
rect 231636 115240 231642 115252
rect 264422 115240 264428 115252
rect 231636 115212 264428 115240
rect 231636 115200 231642 115212
rect 264422 115200 264428 115212
rect 264480 115200 264486 115252
rect 231762 115132 231768 115184
rect 231820 115172 231826 115184
rect 238202 115172 238208 115184
rect 231820 115144 238208 115172
rect 231820 115132 231826 115144
rect 238202 115132 238208 115144
rect 238260 115132 238266 115184
rect 209130 114588 209136 114640
rect 209188 114628 209194 114640
rect 214006 114628 214012 114640
rect 209188 114600 214012 114628
rect 209188 114588 209194 114600
rect 214006 114588 214012 114600
rect 214064 114588 214070 114640
rect 172054 114520 172060 114572
rect 172112 114560 172118 114572
rect 213914 114560 213920 114572
rect 172112 114532 213920 114560
rect 172112 114520 172118 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 246482 114520 246488 114572
rect 246540 114560 246546 114572
rect 265250 114560 265256 114572
rect 246540 114532 265256 114560
rect 246540 114520 246546 114532
rect 265250 114520 265256 114532
rect 265308 114520 265314 114572
rect 230566 114452 230572 114504
rect 230624 114492 230630 114504
rect 232774 114492 232780 114504
rect 230624 114464 232780 114492
rect 230624 114452 230630 114464
rect 232774 114452 232780 114464
rect 232832 114452 232838 114504
rect 230658 114384 230664 114436
rect 230716 114424 230722 114436
rect 239582 114424 239588 114436
rect 230716 114396 239588 114424
rect 230716 114384 230722 114396
rect 239582 114384 239588 114396
rect 239640 114384 239646 114436
rect 231486 114316 231492 114368
rect 231544 114356 231550 114368
rect 245194 114356 245200 114368
rect 231544 114328 245200 114356
rect 231544 114316 231550 114328
rect 245194 114316 245200 114328
rect 245252 114316 245258 114368
rect 282822 113908 282828 113960
rect 282880 113948 282886 113960
rect 288434 113948 288440 113960
rect 282880 113920 288440 113948
rect 282880 113908 282886 113920
rect 288434 113908 288440 113920
rect 288492 113908 288498 113960
rect 256050 113296 256056 113348
rect 256108 113336 256114 113348
rect 265710 113336 265716 113348
rect 256108 113308 265716 113336
rect 256108 113296 256114 113308
rect 265710 113296 265716 113308
rect 265768 113296 265774 113348
rect 187050 113228 187056 113280
rect 187108 113268 187114 113280
rect 213914 113268 213920 113280
rect 187108 113240 213920 113268
rect 187108 113228 187114 113240
rect 213914 113228 213920 113240
rect 213972 113228 213978 113280
rect 245102 113228 245108 113280
rect 245160 113268 245166 113280
rect 265250 113268 265256 113280
rect 245160 113240 265256 113268
rect 245160 113228 245166 113240
rect 265250 113228 265256 113240
rect 265308 113228 265314 113280
rect 167822 113160 167828 113212
rect 167880 113200 167886 113212
rect 214006 113200 214012 113212
rect 167880 113172 214012 113200
rect 167880 113160 167886 113172
rect 214006 113160 214012 113172
rect 214064 113160 214070 113212
rect 235258 113160 235264 113212
rect 235316 113200 235322 113212
rect 265434 113200 265440 113212
rect 235316 113172 265440 113200
rect 235316 113160 235322 113172
rect 265434 113160 265440 113172
rect 265492 113160 265498 113212
rect 230934 113092 230940 113144
rect 230992 113132 230998 113144
rect 241146 113132 241152 113144
rect 230992 113104 241152 113132
rect 230992 113092 230998 113104
rect 241146 113092 241152 113104
rect 241204 113092 241210 113144
rect 282086 113092 282092 113144
rect 282144 113132 282150 113144
rect 294046 113132 294052 113144
rect 282144 113104 294052 113132
rect 282144 113092 282150 113104
rect 294046 113092 294052 113104
rect 294104 113092 294110 113144
rect 231670 112684 231676 112736
rect 231728 112724 231734 112736
rect 234154 112724 234160 112736
rect 231728 112696 234160 112724
rect 231728 112684 231734 112696
rect 234154 112684 234160 112696
rect 234212 112684 234218 112736
rect 231486 112412 231492 112464
rect 231544 112452 231550 112464
rect 258718 112452 258724 112464
rect 231544 112424 258724 112452
rect 231544 112412 231550 112424
rect 258718 112412 258724 112424
rect 258776 112412 258782 112464
rect 260282 111936 260288 111988
rect 260340 111976 260346 111988
rect 265710 111976 265716 111988
rect 260340 111948 265716 111976
rect 260340 111936 260346 111948
rect 265710 111936 265716 111948
rect 265768 111936 265774 111988
rect 211890 111868 211896 111920
rect 211948 111908 211954 111920
rect 214006 111908 214012 111920
rect 211948 111880 214012 111908
rect 211948 111868 211954 111880
rect 214006 111868 214012 111880
rect 214064 111868 214070 111920
rect 242158 111868 242164 111920
rect 242216 111908 242222 111920
rect 265526 111908 265532 111920
rect 242216 111880 265532 111908
rect 242216 111868 242222 111880
rect 265526 111868 265532 111880
rect 265584 111868 265590 111920
rect 166442 111800 166448 111852
rect 166500 111840 166506 111852
rect 213914 111840 213920 111852
rect 166500 111812 213920 111840
rect 166500 111800 166506 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 240962 111800 240968 111852
rect 241020 111840 241026 111852
rect 266078 111840 266084 111852
rect 241020 111812 266084 111840
rect 241020 111800 241026 111812
rect 266078 111800 266084 111812
rect 266136 111800 266142 111852
rect 231762 111732 231768 111784
rect 231820 111772 231826 111784
rect 261846 111772 261852 111784
rect 231820 111744 261852 111772
rect 231820 111732 231826 111744
rect 261846 111732 261852 111744
rect 261904 111732 261910 111784
rect 282822 111732 282828 111784
rect 282880 111772 282886 111784
rect 299566 111772 299572 111784
rect 282880 111744 299572 111772
rect 282880 111732 282886 111744
rect 299566 111732 299572 111744
rect 299624 111732 299630 111784
rect 231670 111664 231676 111716
rect 231728 111704 231734 111716
rect 241054 111704 241060 111716
rect 231728 111676 241060 111704
rect 231728 111664 231734 111676
rect 241054 111664 241060 111676
rect 241112 111664 241118 111716
rect 231670 111052 231676 111104
rect 231728 111092 231734 111104
rect 245010 111092 245016 111104
rect 231728 111064 245016 111092
rect 231728 111052 231734 111064
rect 245010 111052 245016 111064
rect 245068 111052 245074 111104
rect 3418 110848 3424 110900
rect 3476 110888 3482 110900
rect 7558 110888 7564 110900
rect 3476 110860 7564 110888
rect 3476 110848 3482 110860
rect 7558 110848 7564 110860
rect 7616 110848 7622 110900
rect 258902 110576 258908 110628
rect 258960 110616 258966 110628
rect 265526 110616 265532 110628
rect 258960 110588 265532 110616
rect 258960 110576 258966 110588
rect 265526 110576 265532 110588
rect 265584 110576 265590 110628
rect 196710 110508 196716 110560
rect 196768 110548 196774 110560
rect 213914 110548 213920 110560
rect 196768 110520 213920 110548
rect 196768 110508 196774 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 261570 110508 261576 110560
rect 261628 110548 261634 110560
rect 265158 110548 265164 110560
rect 261628 110520 265164 110548
rect 261628 110508 261634 110520
rect 265158 110508 265164 110520
rect 265216 110508 265222 110560
rect 173250 110440 173256 110492
rect 173308 110480 173314 110492
rect 214006 110480 214012 110492
rect 173308 110452 214012 110480
rect 173308 110440 173314 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 245194 110440 245200 110492
rect 245252 110480 245258 110492
rect 265710 110480 265716 110492
rect 245252 110452 265716 110480
rect 245252 110440 245258 110452
rect 265710 110440 265716 110452
rect 265768 110440 265774 110492
rect 167454 110372 167460 110424
rect 167512 110412 167518 110424
rect 170490 110412 170496 110424
rect 167512 110384 170496 110412
rect 167512 110372 167518 110384
rect 170490 110372 170496 110384
rect 170548 110372 170554 110424
rect 231762 110372 231768 110424
rect 231820 110412 231826 110424
rect 261754 110412 261760 110424
rect 231820 110384 261760 110412
rect 231820 110372 231826 110384
rect 261754 110372 261760 110384
rect 261812 110372 261818 110424
rect 231118 110304 231124 110356
rect 231176 110344 231182 110356
rect 254854 110344 254860 110356
rect 231176 110316 254860 110344
rect 231176 110304 231182 110316
rect 254854 110304 254860 110316
rect 254912 110304 254918 110356
rect 176102 109080 176108 109132
rect 176160 109120 176166 109132
rect 213914 109120 213920 109132
rect 176160 109092 213920 109120
rect 176160 109080 176166 109092
rect 213914 109080 213920 109092
rect 213972 109080 213978 109132
rect 231578 109080 231584 109132
rect 231636 109120 231642 109132
rect 235442 109120 235448 109132
rect 231636 109092 235448 109120
rect 231636 109080 231642 109092
rect 235442 109080 235448 109092
rect 235500 109080 235506 109132
rect 261846 109080 261852 109132
rect 261904 109120 261910 109132
rect 265526 109120 265532 109132
rect 261904 109092 265532 109120
rect 261904 109080 261910 109092
rect 265526 109080 265532 109092
rect 265584 109080 265590 109132
rect 173158 109012 173164 109064
rect 173216 109052 173222 109064
rect 214006 109052 214012 109064
rect 173216 109024 214012 109052
rect 173216 109012 173222 109024
rect 214006 109012 214012 109024
rect 214064 109012 214070 109064
rect 250622 109012 250628 109064
rect 250680 109052 250686 109064
rect 265710 109052 265716 109064
rect 250680 109024 265716 109052
rect 250680 109012 250686 109024
rect 265710 109012 265716 109024
rect 265768 109012 265774 109064
rect 167914 108944 167920 108996
rect 167972 108984 167978 108996
rect 173342 108984 173348 108996
rect 167972 108956 173348 108984
rect 167972 108944 167978 108956
rect 173342 108944 173348 108956
rect 173400 108944 173406 108996
rect 231118 108944 231124 108996
rect 231176 108984 231182 108996
rect 263134 108984 263140 108996
rect 231176 108956 263140 108984
rect 231176 108944 231182 108956
rect 263134 108944 263140 108956
rect 263192 108944 263198 108996
rect 282822 108944 282828 108996
rect 282880 108984 282886 108996
rect 306374 108984 306380 108996
rect 282880 108956 306380 108984
rect 282880 108944 282886 108956
rect 306374 108944 306380 108956
rect 306432 108944 306438 108996
rect 231762 108876 231768 108928
rect 231820 108916 231826 108928
rect 246574 108916 246580 108928
rect 231820 108888 246580 108916
rect 231820 108876 231826 108888
rect 246574 108876 246580 108888
rect 246632 108876 246638 108928
rect 230842 108128 230848 108180
rect 230900 108168 230906 108180
rect 232682 108168 232688 108180
rect 230900 108140 232688 108168
rect 230900 108128 230906 108140
rect 232682 108128 232688 108140
rect 232740 108128 232746 108180
rect 281534 107992 281540 108044
rect 281592 108032 281598 108044
rect 284386 108032 284392 108044
rect 281592 108004 284392 108032
rect 281592 107992 281598 108004
rect 284386 107992 284392 108004
rect 284444 107992 284450 108044
rect 241054 107856 241060 107908
rect 241112 107896 241118 107908
rect 265342 107896 265348 107908
rect 241112 107868 265348 107896
rect 241112 107856 241118 107868
rect 265342 107856 265348 107868
rect 265400 107856 265406 107908
rect 209038 107720 209044 107772
rect 209096 107760 209102 107772
rect 214006 107760 214012 107772
rect 209096 107732 214012 107760
rect 209096 107720 209102 107732
rect 214006 107720 214012 107732
rect 214064 107720 214070 107772
rect 260190 107720 260196 107772
rect 260248 107760 260254 107772
rect 265434 107760 265440 107772
rect 260248 107732 265440 107760
rect 260248 107720 260254 107732
rect 265434 107720 265440 107732
rect 265492 107720 265498 107772
rect 202230 107652 202236 107704
rect 202288 107692 202294 107704
rect 213914 107692 213920 107704
rect 202288 107664 213920 107692
rect 202288 107652 202294 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 263042 107652 263048 107704
rect 263100 107692 263106 107704
rect 265710 107692 265716 107704
rect 263100 107664 265716 107692
rect 263100 107652 263106 107664
rect 265710 107652 265716 107664
rect 265768 107652 265774 107704
rect 231762 107584 231768 107636
rect 231820 107624 231826 107636
rect 249334 107624 249340 107636
rect 231820 107596 249340 107624
rect 231820 107584 231826 107596
rect 249334 107584 249340 107596
rect 249392 107584 249398 107636
rect 282454 107584 282460 107636
rect 282512 107624 282518 107636
rect 298278 107624 298284 107636
rect 282512 107596 298284 107624
rect 282512 107584 282518 107596
rect 298278 107584 298284 107596
rect 298336 107584 298342 107636
rect 230566 107516 230572 107568
rect 230624 107556 230630 107568
rect 232590 107556 232596 107568
rect 230624 107528 232596 107556
rect 230624 107516 230630 107528
rect 232590 107516 232596 107528
rect 232648 107516 232654 107568
rect 231394 106904 231400 106956
rect 231452 106944 231458 106956
rect 264606 106944 264612 106956
rect 231452 106916 264612 106944
rect 231452 106904 231458 106916
rect 264606 106904 264612 106916
rect 264664 106904 264670 106956
rect 265434 106768 265440 106820
rect 265492 106808 265498 106820
rect 265802 106808 265808 106820
rect 265492 106780 265808 106808
rect 265492 106768 265498 106780
rect 265802 106768 265808 106780
rect 265860 106768 265866 106820
rect 259086 106428 259092 106480
rect 259144 106468 259150 106480
rect 265802 106468 265808 106480
rect 259144 106440 265808 106468
rect 259144 106428 259150 106440
rect 265802 106428 265808 106440
rect 265860 106428 265866 106480
rect 210510 106360 210516 106412
rect 210568 106400 210574 106412
rect 214006 106400 214012 106412
rect 210568 106372 214012 106400
rect 210568 106360 210574 106372
rect 214006 106360 214012 106372
rect 214064 106360 214070 106412
rect 263134 106360 263140 106412
rect 263192 106400 263198 106412
rect 265526 106400 265532 106412
rect 263192 106372 265532 106400
rect 263192 106360 263198 106372
rect 265526 106360 265532 106372
rect 265584 106360 265590 106412
rect 170490 106292 170496 106344
rect 170548 106332 170554 106344
rect 213914 106332 213920 106344
rect 170548 106304 213920 106332
rect 170548 106292 170554 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 249058 106292 249064 106344
rect 249116 106332 249122 106344
rect 265710 106332 265716 106344
rect 249116 106304 265716 106332
rect 249116 106292 249122 106304
rect 265710 106292 265716 106304
rect 265768 106292 265774 106344
rect 231762 106224 231768 106276
rect 231820 106264 231826 106276
rect 258994 106264 259000 106276
rect 231820 106236 259000 106264
rect 231820 106224 231826 106236
rect 258994 106224 259000 106236
rect 259052 106224 259058 106276
rect 282822 106224 282828 106276
rect 282880 106264 282886 106276
rect 305086 106264 305092 106276
rect 282880 106236 305092 106264
rect 282880 106224 282886 106236
rect 305086 106224 305092 106236
rect 305144 106224 305150 106276
rect 231670 106156 231676 106208
rect 231728 106196 231734 106208
rect 238386 106196 238392 106208
rect 231728 106168 238392 106196
rect 231728 106156 231734 106168
rect 238386 106156 238392 106168
rect 238444 106156 238450 106208
rect 230474 105544 230480 105596
rect 230532 105584 230538 105596
rect 256326 105584 256332 105596
rect 230532 105556 256332 105584
rect 230532 105544 230538 105556
rect 256326 105544 256332 105556
rect 256384 105544 256390 105596
rect 169294 105000 169300 105052
rect 169352 105040 169358 105052
rect 214006 105040 214012 105052
rect 169352 105012 214012 105040
rect 169352 105000 169358 105012
rect 214006 105000 214012 105012
rect 214064 105000 214070 105052
rect 258718 105000 258724 105052
rect 258776 105040 258782 105052
rect 266078 105040 266084 105052
rect 258776 105012 266084 105040
rect 258776 105000 258782 105012
rect 266078 105000 266084 105012
rect 266136 105000 266142 105052
rect 204990 104932 204996 104984
rect 205048 104972 205054 104984
rect 213914 104972 213920 104984
rect 205048 104944 213920 104972
rect 205048 104932 205054 104944
rect 213914 104932 213920 104944
rect 213972 104932 213978 104984
rect 255958 104932 255964 104984
rect 256016 104972 256022 104984
rect 265710 104972 265716 104984
rect 256016 104944 265716 104972
rect 256016 104932 256022 104944
rect 265710 104932 265716 104944
rect 265768 104932 265774 104984
rect 246574 104864 246580 104916
rect 246632 104904 246638 104916
rect 265802 104904 265808 104916
rect 246632 104876 265808 104904
rect 246632 104864 246638 104876
rect 265802 104864 265808 104876
rect 265860 104864 265866 104916
rect 231762 104796 231768 104848
rect 231820 104836 231826 104848
rect 245286 104836 245292 104848
rect 231820 104808 245292 104836
rect 231820 104796 231826 104808
rect 245286 104796 245292 104808
rect 245344 104796 245350 104848
rect 231578 104660 231584 104712
rect 231636 104700 231642 104712
rect 234062 104700 234068 104712
rect 231636 104672 234068 104700
rect 231636 104660 231642 104672
rect 234062 104660 234068 104672
rect 234120 104660 234126 104712
rect 235902 104116 235908 104168
rect 235960 104156 235966 104168
rect 265434 104156 265440 104168
rect 235960 104128 265440 104156
rect 235960 104116 235966 104128
rect 265434 104116 265440 104128
rect 265492 104116 265498 104168
rect 230658 103776 230664 103828
rect 230716 103816 230722 103828
rect 235350 103816 235356 103828
rect 230716 103788 235356 103816
rect 230716 103776 230722 103788
rect 235350 103776 235356 103788
rect 235408 103776 235414 103828
rect 205082 103504 205088 103556
rect 205140 103544 205146 103556
rect 213914 103544 213920 103556
rect 205140 103516 213920 103544
rect 205140 103504 205146 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 245010 103504 245016 103556
rect 245068 103544 245074 103556
rect 265802 103544 265808 103556
rect 245068 103516 265808 103544
rect 245068 103504 245074 103516
rect 265802 103504 265808 103516
rect 265860 103504 265866 103556
rect 231762 103436 231768 103488
rect 231820 103476 231826 103488
rect 252094 103476 252100 103488
rect 231820 103448 252100 103476
rect 231820 103436 231826 103448
rect 252094 103436 252100 103448
rect 252152 103436 252158 103488
rect 282822 103436 282828 103488
rect 282880 103476 282886 103488
rect 299658 103476 299664 103488
rect 282880 103448 299664 103476
rect 282880 103436 282886 103448
rect 299658 103436 299664 103448
rect 299716 103436 299722 103488
rect 231578 103300 231584 103352
rect 231636 103340 231642 103352
rect 233970 103340 233976 103352
rect 231636 103312 233976 103340
rect 231636 103300 231642 103312
rect 233970 103300 233976 103312
rect 234028 103300 234034 103352
rect 249334 102212 249340 102264
rect 249392 102252 249398 102264
rect 265802 102252 265808 102264
rect 249392 102224 265808 102252
rect 249392 102212 249398 102224
rect 265802 102212 265808 102224
rect 265860 102212 265866 102264
rect 232498 102144 232504 102196
rect 232556 102184 232562 102196
rect 265710 102184 265716 102196
rect 232556 102156 265716 102184
rect 232556 102144 232562 102156
rect 265710 102144 265716 102156
rect 265768 102144 265774 102196
rect 230566 102076 230572 102128
rect 230624 102116 230630 102128
rect 242250 102116 242256 102128
rect 230624 102088 242256 102116
rect 230624 102076 230630 102088
rect 242250 102076 242256 102088
rect 242308 102076 242314 102128
rect 231118 102008 231124 102060
rect 231176 102048 231182 102060
rect 235902 102048 235908 102060
rect 231176 102020 235908 102048
rect 231176 102008 231182 102020
rect 235902 102008 235908 102020
rect 235960 102008 235966 102060
rect 167914 101396 167920 101448
rect 167972 101436 167978 101448
rect 214558 101436 214564 101448
rect 167972 101408 214564 101436
rect 167972 101396 167978 101408
rect 214558 101396 214564 101408
rect 214616 101396 214622 101448
rect 254854 100852 254860 100904
rect 254912 100892 254918 100904
rect 265526 100892 265532 100904
rect 254912 100864 265532 100892
rect 254912 100852 254918 100864
rect 265526 100852 265532 100864
rect 265584 100852 265590 100904
rect 207750 100784 207756 100836
rect 207808 100824 207814 100836
rect 214006 100824 214012 100836
rect 207808 100796 214012 100824
rect 207808 100784 207814 100796
rect 214006 100784 214012 100796
rect 214064 100784 214070 100836
rect 242434 100784 242440 100836
rect 242492 100824 242498 100836
rect 265710 100824 265716 100836
rect 242492 100796 265716 100824
rect 242492 100784 242498 100796
rect 265710 100784 265716 100796
rect 265768 100784 265774 100836
rect 184290 100716 184296 100768
rect 184348 100756 184354 100768
rect 213914 100756 213920 100768
rect 184348 100728 213920 100756
rect 184348 100716 184354 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 238202 100716 238208 100768
rect 238260 100756 238266 100768
rect 265802 100756 265808 100768
rect 238260 100728 265808 100756
rect 238260 100716 238266 100728
rect 265802 100716 265808 100728
rect 265860 100716 265866 100768
rect 231670 100648 231676 100700
rect 231728 100688 231734 100700
rect 260374 100688 260380 100700
rect 231728 100660 260380 100688
rect 231728 100648 231734 100660
rect 260374 100648 260380 100660
rect 260432 100648 260438 100700
rect 385678 100648 385684 100700
rect 385736 100688 385742 100700
rect 580166 100688 580172 100700
rect 385736 100660 580172 100688
rect 385736 100648 385742 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 231762 100580 231768 100632
rect 231820 100620 231826 100632
rect 243722 100620 243728 100632
rect 231820 100592 243728 100620
rect 231820 100580 231826 100592
rect 243722 100580 243728 100592
rect 243780 100580 243786 100632
rect 260466 99492 260472 99544
rect 260524 99532 260530 99544
rect 265802 99532 265808 99544
rect 260524 99504 265808 99532
rect 260524 99492 260530 99504
rect 265802 99492 265808 99504
rect 265860 99492 265866 99544
rect 252094 99424 252100 99476
rect 252152 99464 252158 99476
rect 265710 99464 265716 99476
rect 252152 99436 265716 99464
rect 252152 99424 252158 99436
rect 265710 99424 265716 99436
rect 265768 99424 265774 99476
rect 164878 99356 164884 99408
rect 164936 99396 164942 99408
rect 213914 99396 213920 99408
rect 164936 99368 213920 99396
rect 164936 99356 164942 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 243630 99356 243636 99408
rect 243688 99396 243694 99408
rect 265526 99396 265532 99408
rect 243688 99368 265532 99396
rect 243688 99356 243694 99368
rect 265526 99356 265532 99368
rect 265584 99356 265590 99408
rect 265802 99356 265808 99408
rect 265860 99396 265866 99408
rect 266078 99396 266084 99408
rect 265860 99368 266084 99396
rect 265860 99356 265866 99368
rect 266078 99356 266084 99368
rect 266136 99356 266142 99408
rect 231486 99288 231492 99340
rect 231544 99328 231550 99340
rect 242526 99328 242532 99340
rect 231544 99300 242532 99328
rect 231544 99288 231550 99300
rect 242526 99288 242532 99300
rect 242584 99288 242590 99340
rect 282822 99288 282828 99340
rect 282880 99328 282886 99340
rect 299474 99328 299480 99340
rect 282880 99300 299480 99328
rect 282880 99288 282886 99300
rect 299474 99288 299480 99300
rect 299532 99288 299538 99340
rect 209222 98064 209228 98116
rect 209280 98104 209286 98116
rect 213914 98104 213920 98116
rect 209280 98076 213920 98104
rect 209280 98064 209286 98076
rect 213914 98064 213920 98076
rect 213972 98064 213978 98116
rect 242342 98064 242348 98116
rect 242400 98104 242406 98116
rect 265802 98104 265808 98116
rect 242400 98076 265808 98104
rect 242400 98064 242406 98076
rect 265802 98064 265808 98076
rect 265860 98064 265866 98116
rect 166534 97996 166540 98048
rect 166592 98036 166598 98048
rect 214006 98036 214012 98048
rect 166592 98008 214012 98036
rect 166592 97996 166598 98008
rect 214006 97996 214012 98008
rect 214064 97996 214070 98048
rect 235350 97996 235356 98048
rect 235408 98036 235414 98048
rect 265434 98036 265440 98048
rect 235408 98008 265440 98036
rect 235408 97996 235414 98008
rect 265434 97996 265440 98008
rect 265492 97996 265498 98048
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 21358 97968 21364 97980
rect 3476 97940 21364 97968
rect 3476 97928 3482 97940
rect 21358 97928 21364 97940
rect 21416 97928 21422 97980
rect 242250 96704 242256 96756
rect 242308 96744 242314 96756
rect 265158 96744 265164 96756
rect 242308 96716 265164 96744
rect 242308 96704 242314 96716
rect 265158 96704 265164 96716
rect 265216 96704 265222 96756
rect 207658 96636 207664 96688
rect 207716 96676 207722 96688
rect 213914 96676 213920 96688
rect 207716 96648 213920 96676
rect 207716 96636 207722 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 234062 96636 234068 96688
rect 234120 96676 234126 96688
rect 265802 96676 265808 96688
rect 234120 96648 265808 96676
rect 234120 96636 234126 96648
rect 265802 96636 265808 96648
rect 265860 96636 265866 96688
rect 193122 96568 193128 96620
rect 193180 96608 193186 96620
rect 229002 96608 229008 96620
rect 193180 96580 229008 96608
rect 193180 96568 193186 96580
rect 229002 96568 229008 96580
rect 229060 96568 229066 96620
rect 266998 96364 267004 96416
rect 267056 96404 267062 96416
rect 281534 96404 281540 96416
rect 267056 96376 281540 96404
rect 267056 96364 267062 96376
rect 281534 96364 281540 96376
rect 281592 96364 281598 96416
rect 229002 95888 229008 95940
rect 229060 95928 229066 95940
rect 230474 95928 230480 95940
rect 229060 95900 230480 95928
rect 229060 95888 229066 95900
rect 230474 95888 230480 95900
rect 230532 95928 230538 95940
rect 268010 95928 268016 95940
rect 230532 95900 268016 95928
rect 230532 95888 230538 95900
rect 268010 95888 268016 95900
rect 268068 95888 268074 95940
rect 228358 95208 228364 95260
rect 228416 95248 228422 95260
rect 265802 95248 265808 95260
rect 228416 95220 265808 95248
rect 228416 95208 228422 95220
rect 265802 95208 265808 95220
rect 265860 95208 265866 95260
rect 187602 95140 187608 95192
rect 187660 95180 187666 95192
rect 280154 95180 280160 95192
rect 187660 95152 280160 95180
rect 187660 95140 187666 95152
rect 280154 95140 280160 95152
rect 280212 95140 280218 95192
rect 215938 95072 215944 95124
rect 215996 95112 216002 95124
rect 281626 95112 281632 95124
rect 215996 95084 281632 95112
rect 215996 95072 216002 95084
rect 281626 95072 281632 95084
rect 281684 95072 281690 95124
rect 63402 95004 63408 95056
rect 63460 95044 63466 95056
rect 205082 95044 205088 95056
rect 63460 95016 205088 95044
rect 63460 95004 63466 95016
rect 205082 95004 205088 95016
rect 205140 95004 205146 95056
rect 267274 95004 267280 95056
rect 267332 95044 267338 95056
rect 279510 95044 279516 95056
rect 267332 95016 279516 95044
rect 267332 95004 267338 95016
rect 279510 95004 279516 95016
rect 279568 95004 279574 95056
rect 267090 94936 267096 94988
rect 267148 94976 267154 94988
rect 280338 94976 280344 94988
rect 267148 94948 280344 94976
rect 267148 94936 267154 94948
rect 280338 94936 280344 94948
rect 280396 94936 280402 94988
rect 122834 94460 122840 94512
rect 122892 94500 122898 94512
rect 214650 94500 214656 94512
rect 122892 94472 214656 94500
rect 122892 94460 122898 94472
rect 214650 94460 214656 94472
rect 214708 94460 214714 94512
rect 128078 93984 128084 94036
rect 128136 94024 128142 94036
rect 171870 94024 171876 94036
rect 128136 93996 171876 94024
rect 128136 93984 128142 93996
rect 171870 93984 171876 93996
rect 171928 93984 171934 94036
rect 112346 93916 112352 93968
rect 112404 93956 112410 93968
rect 173434 93956 173440 93968
rect 112404 93928 173440 93956
rect 112404 93916 112410 93928
rect 173434 93916 173440 93928
rect 173492 93916 173498 93968
rect 105722 93848 105728 93900
rect 105780 93888 105786 93900
rect 186958 93888 186964 93900
rect 105780 93860 186964 93888
rect 105780 93848 105786 93860
rect 186958 93848 186964 93860
rect 187016 93848 187022 93900
rect 231118 93780 231124 93832
rect 231176 93820 231182 93832
rect 253842 93820 253848 93832
rect 231176 93792 253848 93820
rect 231176 93780 231182 93792
rect 253842 93780 253848 93792
rect 253900 93820 253906 93832
rect 253900 93792 258074 93820
rect 253900 93780 253906 93792
rect 258046 93752 258074 93792
rect 268010 93780 268016 93832
rect 268068 93820 268074 93832
rect 276934 93820 276940 93832
rect 268068 93792 276940 93820
rect 268068 93780 268074 93792
rect 276934 93780 276940 93792
rect 276992 93780 276998 93832
rect 270954 93752 270960 93764
rect 258046 93724 270960 93752
rect 270954 93712 270960 93724
rect 271012 93712 271018 93764
rect 151722 93440 151728 93492
rect 151780 93480 151786 93492
rect 169018 93480 169024 93492
rect 151780 93452 169024 93480
rect 151780 93440 151786 93452
rect 169018 93440 169024 93452
rect 169076 93440 169082 93492
rect 134426 93372 134432 93424
rect 134484 93412 134490 93424
rect 174538 93412 174544 93424
rect 134484 93384 174544 93412
rect 134484 93372 134490 93384
rect 174538 93372 174544 93384
rect 174596 93372 174602 93424
rect 121730 93304 121736 93356
rect 121788 93344 121794 93356
rect 166350 93344 166356 93356
rect 121788 93316 166356 93344
rect 121788 93304 121794 93316
rect 166350 93304 166356 93316
rect 166408 93304 166414 93356
rect 88978 93236 88984 93288
rect 89036 93276 89042 93288
rect 164878 93276 164884 93288
rect 89036 93248 164884 93276
rect 89036 93236 89042 93248
rect 164878 93236 164884 93248
rect 164936 93236 164942 93288
rect 111242 93168 111248 93220
rect 111300 93208 111306 93220
rect 191190 93208 191196 93220
rect 111300 93180 191196 93208
rect 111300 93168 111306 93180
rect 191190 93168 191196 93180
rect 191248 93168 191254 93220
rect 230474 93168 230480 93220
rect 230532 93208 230538 93220
rect 233970 93208 233976 93220
rect 230532 93180 233976 93208
rect 230532 93168 230538 93180
rect 233970 93168 233976 93180
rect 234028 93168 234034 93220
rect 106458 93100 106464 93152
rect 106516 93140 106522 93152
rect 209130 93140 209136 93152
rect 106516 93112 209136 93140
rect 106516 93100 106522 93112
rect 209130 93100 209136 93112
rect 209188 93100 209194 93152
rect 216306 92556 216312 92608
rect 216364 92596 216370 92608
rect 220078 92596 220084 92608
rect 216364 92568 220084 92596
rect 216364 92556 216370 92568
rect 220078 92556 220084 92568
rect 220136 92556 220142 92608
rect 180610 92420 180616 92472
rect 180668 92460 180674 92472
rect 281810 92460 281816 92472
rect 180668 92432 281816 92460
rect 180668 92420 180674 92432
rect 281810 92420 281816 92432
rect 281868 92420 281874 92472
rect 98546 92352 98552 92404
rect 98604 92392 98610 92404
rect 196710 92392 196716 92404
rect 98604 92364 196716 92392
rect 98604 92352 98610 92364
rect 196710 92352 196716 92364
rect 196768 92352 196774 92404
rect 118050 92284 118056 92336
rect 118108 92324 118114 92336
rect 202138 92324 202144 92336
rect 118108 92296 202144 92324
rect 118108 92284 118114 92296
rect 202138 92284 202144 92296
rect 202196 92284 202202 92336
rect 110690 92216 110696 92268
rect 110748 92256 110754 92268
rect 122834 92256 122840 92268
rect 110748 92228 122840 92256
rect 110748 92216 110754 92228
rect 122834 92216 122840 92228
rect 122892 92216 122898 92268
rect 126698 92216 126704 92268
rect 126756 92256 126762 92268
rect 188338 92256 188344 92268
rect 126756 92228 188344 92256
rect 126756 92216 126762 92228
rect 188338 92216 188344 92228
rect 188396 92216 188402 92268
rect 133138 92148 133144 92200
rect 133196 92188 133202 92200
rect 167914 92188 167920 92200
rect 133196 92160 167920 92188
rect 133196 92148 133202 92160
rect 167914 92148 167920 92160
rect 167972 92148 167978 92200
rect 151538 92080 151544 92132
rect 151596 92120 151602 92132
rect 180058 92120 180064 92132
rect 151596 92092 180064 92120
rect 151596 92080 151602 92092
rect 180058 92080 180064 92092
rect 180116 92080 180122 92132
rect 106642 92012 106648 92064
rect 106700 92052 106706 92064
rect 184198 92052 184204 92064
rect 106700 92024 184204 92052
rect 106700 92012 106706 92024
rect 184198 92012 184204 92024
rect 184256 92012 184262 92064
rect 104618 91128 104624 91180
rect 104676 91168 104682 91180
rect 117958 91168 117964 91180
rect 104676 91140 117964 91168
rect 104676 91128 104682 91140
rect 117958 91128 117964 91140
rect 118016 91128 118022 91180
rect 86586 91060 86592 91112
rect 86644 91100 86650 91112
rect 110414 91100 110420 91112
rect 86644 91072 110420 91100
rect 86644 91060 86650 91072
rect 110414 91060 110420 91072
rect 110472 91060 110478 91112
rect 104342 90992 104348 91044
rect 104400 91032 104406 91044
rect 167822 91032 167828 91044
rect 104400 91004 167828 91032
rect 104400 90992 104406 91004
rect 167822 90992 167828 91004
rect 167880 90992 167886 91044
rect 126514 90924 126520 90976
rect 126572 90964 126578 90976
rect 188430 90964 188436 90976
rect 126572 90936 188436 90964
rect 126572 90924 126578 90936
rect 188430 90924 188436 90936
rect 188488 90924 188494 90976
rect 110138 90856 110144 90908
rect 110196 90896 110202 90908
rect 169202 90896 169208 90908
rect 110196 90868 169208 90896
rect 110196 90856 110202 90868
rect 169202 90856 169208 90868
rect 169260 90856 169266 90908
rect 151354 90788 151360 90840
rect 151412 90828 151418 90840
rect 177390 90828 177396 90840
rect 151412 90800 177396 90828
rect 151412 90788 151418 90800
rect 177390 90788 177396 90800
rect 177448 90788 177454 90840
rect 188338 90312 188344 90364
rect 188396 90352 188402 90364
rect 265986 90352 265992 90364
rect 188396 90324 265992 90352
rect 188396 90312 188402 90324
rect 265986 90312 265992 90324
rect 266044 90312 266050 90364
rect 67450 89632 67456 89684
rect 67508 89672 67514 89684
rect 207750 89672 207756 89684
rect 67508 89644 207756 89672
rect 67508 89632 67514 89644
rect 207750 89632 207756 89644
rect 207808 89632 207814 89684
rect 90358 89564 90364 89616
rect 90416 89604 90422 89616
rect 169294 89604 169300 89616
rect 90416 89576 169300 89604
rect 90416 89564 90422 89576
rect 169294 89564 169300 89576
rect 169352 89564 169358 89616
rect 119890 89496 119896 89548
rect 119948 89536 119954 89548
rect 197998 89536 198004 89548
rect 119948 89508 198004 89536
rect 119948 89496 119954 89508
rect 197998 89496 198004 89508
rect 198056 89496 198062 89548
rect 105998 89428 106004 89480
rect 106056 89468 106062 89480
rect 172054 89468 172060 89480
rect 106056 89440 172060 89468
rect 106056 89428 106062 89440
rect 172054 89428 172060 89440
rect 172112 89428 172118 89480
rect 132402 89360 132408 89412
rect 132460 89400 132466 89412
rect 178678 89400 178684 89412
rect 132460 89372 178684 89400
rect 132460 89360 132466 89372
rect 178678 89360 178684 89372
rect 178736 89360 178742 89412
rect 215938 88952 215944 89004
rect 215996 88992 216002 89004
rect 265894 88992 265900 89004
rect 215996 88964 265900 88992
rect 215996 88952 216002 88964
rect 265894 88952 265900 88964
rect 265952 88952 265958 89004
rect 84654 88272 84660 88324
rect 84712 88312 84718 88324
rect 184290 88312 184296 88324
rect 84712 88284 184296 88312
rect 84712 88272 84718 88284
rect 184290 88272 184296 88284
rect 184348 88272 184354 88324
rect 100570 88204 100576 88256
rect 100628 88244 100634 88256
rect 166442 88244 166448 88256
rect 100628 88216 166448 88244
rect 100628 88204 100634 88216
rect 166442 88204 166448 88216
rect 166500 88204 166506 88256
rect 117130 88136 117136 88188
rect 117188 88176 117194 88188
rect 170674 88176 170680 88188
rect 117188 88148 170680 88176
rect 117188 88136 117194 88148
rect 170674 88136 170680 88148
rect 170732 88136 170738 88188
rect 115566 88068 115572 88120
rect 115624 88108 115630 88120
rect 169110 88108 169116 88120
rect 115624 88080 169116 88108
rect 115624 88068 115630 88080
rect 169110 88068 169116 88080
rect 169168 88068 169174 88120
rect 123754 88000 123760 88052
rect 123812 88040 123818 88052
rect 175918 88040 175924 88052
rect 123812 88012 175924 88040
rect 123812 88000 123818 88012
rect 175918 88000 175924 88012
rect 175976 88000 175982 88052
rect 124030 87932 124036 87984
rect 124088 87972 124094 87984
rect 167730 87972 167736 87984
rect 124088 87944 167736 87972
rect 124088 87932 124094 87944
rect 167730 87932 167736 87944
rect 167788 87932 167794 87984
rect 101858 86912 101864 86964
rect 101916 86952 101922 86964
rect 211890 86952 211896 86964
rect 101916 86924 211896 86952
rect 101916 86912 101922 86924
rect 211890 86912 211896 86924
rect 211948 86912 211954 86964
rect 110414 86844 110420 86896
rect 110472 86884 110478 86896
rect 209222 86884 209228 86896
rect 110472 86856 209228 86884
rect 110472 86844 110478 86856
rect 209222 86844 209228 86856
rect 209280 86844 209286 86896
rect 97074 86776 97080 86828
rect 97132 86816 97138 86828
rect 174722 86816 174728 86828
rect 97132 86788 174728 86816
rect 97132 86776 97138 86788
rect 174722 86776 174728 86788
rect 174780 86776 174786 86828
rect 109494 86708 109500 86760
rect 109552 86748 109558 86760
rect 180150 86748 180156 86760
rect 109552 86720 180156 86748
rect 109552 86708 109558 86720
rect 180150 86708 180156 86720
rect 180208 86708 180214 86760
rect 120810 86640 120816 86692
rect 120868 86680 120874 86692
rect 170582 86680 170588 86692
rect 120868 86652 170588 86680
rect 120868 86640 120874 86652
rect 170582 86640 170588 86652
rect 170640 86640 170646 86692
rect 3418 85484 3424 85536
rect 3476 85524 3482 85536
rect 25498 85524 25504 85536
rect 3476 85496 25504 85524
rect 3476 85484 3482 85496
rect 25498 85484 25504 85496
rect 25556 85484 25562 85536
rect 64782 85484 64788 85536
rect 64840 85524 64846 85536
rect 207658 85524 207664 85536
rect 64840 85496 207664 85524
rect 64840 85484 64846 85496
rect 207658 85484 207664 85496
rect 207716 85484 207722 85536
rect 114370 85416 114376 85468
rect 114428 85456 114434 85468
rect 213178 85456 213184 85468
rect 114428 85428 213184 85456
rect 114428 85416 114434 85428
rect 213178 85416 213184 85428
rect 213236 85416 213242 85468
rect 103054 85348 103060 85400
rect 103112 85388 103118 85400
rect 187050 85388 187056 85400
rect 103112 85360 187056 85388
rect 103112 85348 103118 85360
rect 187050 85348 187056 85360
rect 187108 85348 187114 85400
rect 92290 85280 92296 85332
rect 92348 85320 92354 85332
rect 170490 85320 170496 85332
rect 92348 85292 170496 85320
rect 92348 85280 92354 85292
rect 170490 85280 170496 85292
rect 170548 85280 170554 85332
rect 152642 85212 152648 85264
rect 152700 85252 152706 85264
rect 196618 85252 196624 85264
rect 152700 85224 196624 85252
rect 152700 85212 152706 85224
rect 196618 85212 196624 85224
rect 196676 85212 196682 85264
rect 125410 85144 125416 85196
rect 125468 85184 125474 85196
rect 167638 85184 167644 85196
rect 125468 85156 167644 85184
rect 125468 85144 125474 85156
rect 167638 85144 167644 85156
rect 167696 85144 167702 85196
rect 108850 84124 108856 84176
rect 108908 84164 108914 84176
rect 213362 84164 213368 84176
rect 108908 84136 213368 84164
rect 108908 84124 108914 84136
rect 213362 84124 213368 84136
rect 213420 84124 213426 84176
rect 121362 84056 121368 84108
rect 121420 84096 121426 84108
rect 210418 84096 210424 84108
rect 121420 84068 210424 84096
rect 121420 84056 121426 84068
rect 210418 84056 210424 84068
rect 210476 84056 210482 84108
rect 86862 83988 86868 84040
rect 86920 84028 86926 84040
rect 166534 84028 166540 84040
rect 86920 84000 166540 84028
rect 86920 83988 86926 84000
rect 166534 83988 166540 84000
rect 166592 83988 166598 84040
rect 96522 83920 96528 83972
rect 96580 83960 96586 83972
rect 176102 83960 176108 83972
rect 96580 83932 176108 83960
rect 96580 83920 96586 83932
rect 176102 83920 176108 83932
rect 176160 83920 176166 83972
rect 115842 83852 115848 83904
rect 115900 83892 115906 83904
rect 178770 83892 178776 83904
rect 115900 83864 178776 83892
rect 115900 83852 115906 83864
rect 178770 83852 178776 83864
rect 178828 83852 178834 83904
rect 136542 83784 136548 83836
rect 136600 83824 136606 83836
rect 166258 83824 166264 83836
rect 136600 83796 166264 83824
rect 136600 83784 136606 83796
rect 166258 83784 166264 83796
rect 166316 83784 166322 83836
rect 75822 82764 75828 82816
rect 75880 82804 75886 82816
rect 214558 82804 214564 82816
rect 75880 82776 214564 82804
rect 75880 82764 75886 82776
rect 214558 82764 214564 82776
rect 214616 82764 214622 82816
rect 114462 82696 114468 82748
rect 114520 82736 114526 82748
rect 213270 82736 213276 82748
rect 114520 82708 213276 82736
rect 114520 82696 114526 82708
rect 213270 82696 213276 82708
rect 213328 82696 213334 82748
rect 103422 82628 103428 82680
rect 103480 82668 103486 82680
rect 176010 82668 176016 82680
rect 103480 82640 176016 82668
rect 103480 82628 103486 82640
rect 176010 82628 176016 82640
rect 176068 82628 176074 82680
rect 125502 82560 125508 82612
rect 125560 82600 125566 82612
rect 170398 82600 170404 82612
rect 125560 82572 170404 82600
rect 125560 82560 125566 82572
rect 170398 82560 170404 82572
rect 170456 82560 170462 82612
rect 95050 81336 95056 81388
rect 95108 81376 95114 81388
rect 202230 81376 202236 81388
rect 95108 81348 202236 81376
rect 95108 81336 95114 81348
rect 202230 81336 202236 81348
rect 202288 81336 202294 81388
rect 118602 81268 118608 81320
rect 118660 81308 118666 81320
rect 211798 81308 211804 81320
rect 118660 81280 211804 81308
rect 118660 81268 118666 81280
rect 211798 81268 211804 81280
rect 211856 81268 211862 81320
rect 129642 81200 129648 81252
rect 129700 81240 129706 81252
rect 177298 81240 177304 81252
rect 129700 81212 177304 81240
rect 129700 81200 129706 81212
rect 177298 81200 177304 81212
rect 177356 81200 177362 81252
rect 93762 79976 93768 80028
rect 93820 80016 93826 80028
rect 210510 80016 210516 80028
rect 93820 79988 210516 80016
rect 93820 79976 93826 79988
rect 210510 79976 210516 79988
rect 210568 79976 210574 80028
rect 117222 79908 117228 79960
rect 117280 79948 117286 79960
rect 206370 79948 206376 79960
rect 117280 79920 206376 79948
rect 117280 79908 117286 79920
rect 206370 79908 206376 79920
rect 206428 79908 206434 79960
rect 124122 79840 124128 79892
rect 124180 79880 124186 79892
rect 199378 79880 199384 79892
rect 124180 79852 199384 79880
rect 124180 79840 124186 79852
rect 199378 79840 199384 79852
rect 199436 79840 199442 79892
rect 100662 79772 100668 79824
rect 100720 79812 100726 79824
rect 173250 79812 173256 79824
rect 100720 79784 173256 79812
rect 100720 79772 100726 79784
rect 173250 79772 173256 79784
rect 173308 79772 173314 79824
rect 108942 79704 108948 79756
rect 109000 79744 109006 79756
rect 171778 79744 171784 79756
rect 109000 79716 171784 79744
rect 109000 79704 109006 79716
rect 171778 79704 171784 79716
rect 171836 79704 171842 79756
rect 95142 78616 95148 78668
rect 95200 78656 95206 78668
rect 209038 78656 209044 78668
rect 95200 78628 209044 78656
rect 95200 78616 95206 78628
rect 209038 78616 209044 78628
rect 209096 78616 209102 78668
rect 110322 78548 110328 78600
rect 110380 78588 110386 78600
rect 204898 78588 204904 78600
rect 110380 78560 204904 78588
rect 110380 78548 110386 78560
rect 204898 78548 204904 78560
rect 204956 78548 204962 78600
rect 99282 78480 99288 78532
rect 99340 78520 99346 78532
rect 177482 78520 177488 78532
rect 99340 78492 177488 78520
rect 99340 78480 99346 78492
rect 177482 78480 177488 78492
rect 177540 78480 177546 78532
rect 102042 78412 102048 78464
rect 102100 78452 102106 78464
rect 174630 78452 174636 78464
rect 102100 78424 174636 78452
rect 102100 78412 102106 78424
rect 174630 78412 174636 78424
rect 174688 78412 174694 78464
rect 67542 77188 67548 77240
rect 67600 77228 67606 77240
rect 214742 77228 214748 77240
rect 67600 77200 214748 77228
rect 67600 77188 67606 77200
rect 214742 77188 214748 77200
rect 214800 77188 214806 77240
rect 97902 77120 97908 77172
rect 97960 77160 97966 77172
rect 173158 77160 173164 77172
rect 97960 77132 173164 77160
rect 97960 77120 97966 77132
rect 173158 77120 173164 77132
rect 173216 77120 173222 77172
rect 13814 76508 13820 76560
rect 13872 76548 13878 76560
rect 252002 76548 252008 76560
rect 13872 76520 252008 76548
rect 13872 76508 13878 76520
rect 252002 76508 252008 76520
rect 252060 76508 252066 76560
rect 125594 75284 125600 75336
rect 125652 75324 125658 75336
rect 191098 75324 191104 75336
rect 125652 75296 191104 75324
rect 125652 75284 125658 75296
rect 191098 75284 191104 75296
rect 191156 75284 191162 75336
rect 95234 75216 95240 75268
rect 95292 75256 95298 75268
rect 253382 75256 253388 75268
rect 95292 75228 253388 75256
rect 95292 75216 95298 75228
rect 253382 75216 253388 75228
rect 253440 75216 253446 75268
rect 75914 75148 75920 75200
rect 75972 75188 75978 75200
rect 259086 75188 259092 75200
rect 75972 75160 259092 75188
rect 75972 75148 75978 75160
rect 259086 75148 259092 75160
rect 259144 75148 259150 75200
rect 117958 74468 117964 74520
rect 118016 74508 118022 74520
rect 206278 74508 206284 74520
rect 118016 74480 206284 74508
rect 118016 74468 118022 74480
rect 206278 74468 206284 74480
rect 206336 74468 206342 74520
rect 99374 73856 99380 73908
rect 99432 73896 99438 73908
rect 249242 73896 249248 73908
rect 99432 73868 249248 73896
rect 99432 73856 99438 73868
rect 249242 73856 249248 73868
rect 249300 73856 249306 73908
rect 78674 73788 78680 73840
rect 78732 73828 78738 73840
rect 263134 73828 263140 73840
rect 78732 73800 263140 73828
rect 78732 73788 78738 73800
rect 263134 73788 263140 73800
rect 263192 73788 263198 73840
rect 96614 72428 96620 72480
rect 96672 72468 96678 72480
rect 250622 72468 250628 72480
rect 96672 72440 250628 72468
rect 96672 72428 96678 72440
rect 250622 72428 250628 72440
rect 250680 72428 250686 72480
rect 74534 69708 74540 69760
rect 74592 69748 74598 69760
rect 229830 69748 229836 69760
rect 74592 69720 229836 69748
rect 74592 69708 74598 69720
rect 229830 69708 229836 69720
rect 229888 69708 229894 69760
rect 100754 69640 100760 69692
rect 100812 69680 100818 69692
rect 261846 69680 261852 69692
rect 100812 69652 261852 69680
rect 100812 69640 100818 69652
rect 261846 69640 261852 69652
rect 261904 69640 261910 69692
rect 107654 68348 107660 68400
rect 107712 68388 107718 68400
rect 245194 68388 245200 68400
rect 107712 68360 245200 68388
rect 107712 68348 107718 68360
rect 245194 68348 245200 68360
rect 245252 68348 245258 68400
rect 52454 68280 52460 68332
rect 52512 68320 52518 68332
rect 247862 68320 247868 68332
rect 52512 68292 247868 68320
rect 52512 68280 52518 68292
rect 247862 68280 247868 68292
rect 247920 68280 247926 68332
rect 103514 66920 103520 66972
rect 103572 66960 103578 66972
rect 264514 66960 264520 66972
rect 103572 66932 264520 66960
rect 103572 66920 103578 66932
rect 264514 66920 264520 66932
rect 264572 66920 264578 66972
rect 41414 66852 41420 66904
rect 41472 66892 41478 66904
rect 256234 66892 256240 66904
rect 41472 66864 256240 66892
rect 41472 66852 41478 66864
rect 256234 66852 256240 66864
rect 256292 66852 256298 66904
rect 110414 65560 110420 65612
rect 110472 65600 110478 65612
rect 247770 65600 247776 65612
rect 110472 65572 247776 65600
rect 110472 65560 110478 65572
rect 247770 65560 247776 65572
rect 247828 65560 247834 65612
rect 16574 65492 16580 65544
rect 16632 65532 16638 65544
rect 260466 65532 260472 65544
rect 16632 65504 260472 65532
rect 16632 65492 16638 65504
rect 260466 65492 260472 65504
rect 260524 65492 260530 65544
rect 121454 64200 121460 64252
rect 121512 64240 121518 64252
rect 260282 64240 260288 64252
rect 121512 64212 260288 64240
rect 121512 64200 121518 64212
rect 260282 64200 260288 64212
rect 260340 64200 260346 64252
rect 30374 64132 30380 64184
rect 30432 64172 30438 64184
rect 246482 64172 246488 64184
rect 30432 64144 246488 64172
rect 30432 64132 30438 64144
rect 246482 64132 246488 64144
rect 246540 64132 246546 64184
rect 20714 62772 20720 62824
rect 20772 62812 20778 62824
rect 252094 62812 252100 62824
rect 20772 62784 252100 62812
rect 20772 62772 20778 62784
rect 252094 62772 252100 62784
rect 252152 62772 252158 62824
rect 64874 61412 64880 61464
rect 64932 61452 64938 61464
rect 246574 61452 246580 61464
rect 64932 61424 246580 61452
rect 64932 61412 64938 61424
rect 246574 61412 246580 61424
rect 246632 61412 246638 61464
rect 28994 61344 29000 61396
rect 29052 61384 29058 61396
rect 242434 61384 242440 61396
rect 29052 61356 242440 61384
rect 29052 61344 29058 61356
rect 242434 61344 242440 61356
rect 242492 61344 242498 61396
rect 82814 60052 82820 60104
rect 82872 60092 82878 60104
rect 241054 60092 241060 60104
rect 82872 60064 241060 60092
rect 82872 60052 82878 60064
rect 241054 60052 241060 60064
rect 241112 60052 241118 60104
rect 33134 59984 33140 60036
rect 33192 60024 33198 60036
rect 254854 60024 254860 60036
rect 33192 59996 254860 60024
rect 33192 59984 33198 59996
rect 254854 59984 254860 59996
rect 254912 59984 254918 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 43438 59344 43444 59356
rect 3108 59316 43444 59344
rect 3108 59304 3114 59316
rect 43438 59304 43444 59316
rect 43496 59304 43502 59356
rect 122834 58692 122840 58744
rect 122892 58732 122898 58744
rect 257614 58732 257620 58744
rect 122892 58704 257620 58732
rect 122892 58692 122898 58704
rect 257614 58692 257620 58704
rect 257672 58692 257678 58744
rect 43530 58624 43536 58676
rect 43588 58664 43594 58676
rect 231118 58664 231124 58676
rect 43588 58636 231124 58664
rect 43588 58624 43594 58636
rect 231118 58624 231124 58636
rect 231176 58624 231182 58676
rect 93854 57196 93860 57248
rect 93912 57236 93918 57248
rect 263042 57236 263048 57248
rect 93912 57208 263048 57236
rect 93912 57196 93918 57208
rect 263042 57196 263048 57208
rect 263100 57196 263106 57248
rect 118694 55836 118700 55888
rect 118752 55876 118758 55888
rect 240962 55876 240968 55888
rect 118752 55848 240968 55876
rect 118752 55836 118758 55848
rect 240962 55836 240968 55848
rect 241020 55836 241026 55888
rect 97994 54544 98000 54596
rect 98052 54584 98058 54596
rect 250530 54584 250536 54596
rect 98052 54556 250536 54584
rect 98052 54544 98058 54556
rect 250530 54544 250536 54556
rect 250588 54544 250594 54596
rect 55214 54476 55220 54528
rect 55272 54516 55278 54528
rect 262950 54516 262956 54528
rect 55272 54488 262956 54516
rect 55272 54476 55278 54488
rect 262950 54476 262956 54488
rect 263008 54476 263014 54528
rect 109034 53116 109040 53168
rect 109092 53156 109098 53168
rect 251910 53156 251916 53168
rect 109092 53128 251916 53156
rect 109092 53116 109098 53128
rect 251910 53116 251916 53128
rect 251968 53116 251974 53168
rect 24854 53048 24860 53100
rect 24912 53088 24918 53100
rect 242342 53088 242348 53100
rect 24912 53060 242348 53088
rect 24912 53048 24918 53060
rect 242342 53048 242348 53060
rect 242400 53048 242406 53100
rect 35894 51688 35900 51740
rect 35952 51728 35958 51740
rect 249334 51728 249340 51740
rect 35952 51700 249340 51728
rect 35952 51688 35958 51700
rect 249334 51688 249340 51700
rect 249392 51688 249398 51740
rect 66254 50396 66260 50448
rect 66312 50436 66318 50448
rect 256142 50436 256148 50448
rect 66312 50408 256148 50436
rect 66312 50396 66318 50408
rect 256142 50396 256148 50408
rect 256200 50396 256206 50448
rect 19334 50328 19340 50380
rect 19392 50368 19398 50380
rect 235350 50368 235356 50380
rect 19392 50340 235356 50368
rect 19392 50328 19398 50340
rect 235350 50328 235356 50340
rect 235408 50328 235414 50380
rect 69014 49036 69020 49088
rect 69072 49076 69078 49088
rect 254762 49076 254768 49088
rect 69072 49048 254768 49076
rect 69072 49036 69078 49048
rect 254762 49036 254768 49048
rect 254820 49036 254826 49088
rect 15194 48968 15200 49020
rect 15252 49008 15258 49020
rect 234062 49008 234068 49020
rect 15252 48980 234068 49008
rect 15252 48968 15258 48980
rect 234062 48968 234068 48980
rect 234120 48968 234126 49020
rect 11054 47540 11060 47592
rect 11112 47580 11118 47592
rect 242250 47580 242256 47592
rect 11112 47552 242256 47580
rect 11112 47540 11118 47552
rect 242250 47540 242256 47552
rect 242308 47540 242314 47592
rect 322198 46860 322204 46912
rect 322256 46900 322262 46912
rect 580166 46900 580172 46912
rect 322256 46872 580172 46900
rect 322256 46860 322262 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 115934 46180 115940 46232
rect 115992 46220 115998 46232
rect 240870 46220 240876 46232
rect 115992 46192 240876 46220
rect 115992 46180 115998 46192
rect 240870 46180 240876 46192
rect 240928 46180 240934 46232
rect 2866 45500 2872 45552
rect 2924 45540 2930 45552
rect 4798 45540 4804 45552
rect 2924 45512 4804 45540
rect 2924 45500 2930 45512
rect 4798 45500 4804 45512
rect 4856 45500 4862 45552
rect 111794 44820 111800 44872
rect 111852 44860 111858 44872
rect 249150 44860 249156 44872
rect 111852 44832 249156 44860
rect 111852 44820 111858 44832
rect 249150 44820 249156 44832
rect 249208 44820 249214 44872
rect 56594 43392 56600 43444
rect 56652 43432 56658 43444
rect 250438 43432 250444 43444
rect 56652 43404 250444 43432
rect 56652 43392 56658 43404
rect 250438 43392 250444 43404
rect 250496 43392 250502 43444
rect 104894 42100 104900 42152
rect 104952 42140 104958 42152
rect 264330 42140 264336 42152
rect 104952 42112 264336 42140
rect 104952 42100 104958 42112
rect 264330 42100 264336 42112
rect 264388 42100 264394 42152
rect 35986 42032 35992 42084
rect 36044 42072 36050 42084
rect 257522 42072 257528 42084
rect 36044 42044 257528 42072
rect 36044 42032 36050 42044
rect 257522 42032 257528 42044
rect 257580 42032 257586 42084
rect 63494 40672 63500 40724
rect 63552 40712 63558 40724
rect 236638 40712 236644 40724
rect 63552 40684 236644 40712
rect 63552 40672 63558 40684
rect 236638 40672 236644 40684
rect 236696 40672 236702 40724
rect 67634 39380 67640 39432
rect 67692 39420 67698 39432
rect 262858 39420 262864 39432
rect 67692 39392 262864 39420
rect 67692 39380 67698 39392
rect 262858 39380 262864 39392
rect 262916 39380 262922 39432
rect 17954 39312 17960 39364
rect 18012 39352 18018 39364
rect 245102 39352 245108 39364
rect 18012 39324 245108 39352
rect 18012 39312 18018 39324
rect 245102 39312 245108 39324
rect 245160 39312 245166 39364
rect 102134 37952 102140 38004
rect 102192 37992 102198 38004
rect 254670 37992 254676 38004
rect 102192 37964 254676 37992
rect 102192 37952 102198 37964
rect 254670 37952 254676 37964
rect 254728 37952 254734 38004
rect 60734 37884 60740 37936
rect 60792 37924 60798 37936
rect 246298 37924 246304 37936
rect 60792 37896 246304 37924
rect 60792 37884 60798 37896
rect 246298 37884 246304 37896
rect 246356 37884 246362 37936
rect 81434 36524 81440 36576
rect 81492 36564 81498 36576
rect 253290 36564 253296 36576
rect 81492 36536 253296 36564
rect 81492 36524 81498 36536
rect 253290 36524 253296 36536
rect 253348 36524 253354 36576
rect 86954 35232 86960 35284
rect 87012 35272 87018 35284
rect 261662 35272 261668 35284
rect 87012 35244 261668 35272
rect 87012 35232 87018 35244
rect 261662 35232 261668 35244
rect 261720 35232 261726 35284
rect 12434 35164 12440 35216
rect 12492 35204 12498 35216
rect 235258 35204 235264 35216
rect 12492 35176 235264 35204
rect 12492 35164 12498 35176
rect 235258 35164 235264 35176
rect 235316 35164 235322 35216
rect 106918 33736 106924 33788
rect 106976 33776 106982 33788
rect 265618 33776 265624 33788
rect 106976 33748 265624 33776
rect 106976 33736 106982 33748
rect 265618 33736 265624 33748
rect 265676 33736 265682 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 18598 33096 18604 33108
rect 3568 33068 18604 33096
rect 3568 33056 3574 33068
rect 18598 33056 18604 33068
rect 18656 33056 18662 33108
rect 302878 33056 302884 33108
rect 302936 33096 302942 33108
rect 580166 33096 580172 33108
rect 302936 33068 580172 33096
rect 302936 33056 302942 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 85574 32444 85580 32496
rect 85632 32484 85638 32496
rect 238110 32484 238116 32496
rect 85632 32456 238116 32484
rect 85632 32444 85638 32456
rect 238110 32444 238116 32456
rect 238168 32444 238174 32496
rect 53834 32376 53840 32428
rect 53892 32416 53898 32428
rect 265710 32416 265716 32428
rect 53892 32388 265716 32416
rect 53892 32376 53898 32388
rect 265710 32376 265716 32388
rect 265768 32376 265774 32428
rect 52546 31084 52552 31136
rect 52604 31124 52610 31136
rect 239490 31124 239496 31136
rect 52604 31096 239496 31124
rect 52604 31084 52610 31096
rect 239490 31084 239496 31096
rect 239548 31084 239554 31136
rect 59354 31016 59360 31068
rect 59412 31056 59418 31068
rect 257430 31056 257436 31068
rect 59412 31028 257436 31056
rect 59412 31016 59418 31028
rect 257430 31016 257436 31028
rect 257488 31016 257494 31068
rect 80054 29656 80060 29708
rect 80112 29696 80118 29708
rect 258810 29696 258816 29708
rect 80112 29668 258816 29696
rect 80112 29656 80118 29668
rect 258810 29656 258816 29668
rect 258868 29656 258874 29708
rect 48314 29588 48320 29640
rect 48372 29628 48378 29640
rect 246390 29628 246396 29640
rect 48372 29600 246396 29628
rect 48372 29588 48378 29600
rect 246390 29588 246396 29600
rect 246448 29588 246454 29640
rect 88334 28296 88340 28348
rect 88392 28336 88398 28348
rect 261478 28336 261484 28348
rect 88392 28308 261484 28336
rect 88392 28296 88398 28308
rect 261478 28296 261484 28308
rect 261536 28296 261542 28348
rect 8294 28228 8300 28280
rect 8352 28268 8358 28280
rect 242158 28268 242164 28280
rect 8352 28240 242164 28268
rect 8352 28228 8358 28240
rect 242158 28228 242164 28240
rect 242216 28228 242222 28280
rect 57974 26936 57980 26988
rect 58032 26976 58038 26988
rect 264422 26976 264428 26988
rect 58032 26948 264428 26976
rect 58032 26936 58038 26948
rect 264422 26936 264428 26948
rect 264480 26936 264486 26988
rect 22094 26868 22100 26920
rect 22152 26908 22158 26920
rect 256050 26908 256056 26920
rect 22152 26880 256056 26908
rect 22152 26868 22158 26880
rect 256050 26868 256056 26880
rect 256108 26868 256114 26920
rect 114554 25576 114560 25628
rect 114612 25616 114618 25628
rect 258902 25616 258908 25628
rect 114612 25588 258908 25616
rect 114612 25576 114618 25588
rect 258902 25576 258908 25588
rect 258960 25576 258966 25628
rect 26234 25508 26240 25560
rect 26292 25548 26298 25560
rect 238202 25548 238208 25560
rect 26292 25520 238208 25548
rect 26292 25508 26298 25520
rect 238202 25508 238208 25520
rect 238260 25508 238266 25560
rect 110506 24148 110512 24200
rect 110564 24188 110570 24200
rect 261570 24188 261576 24200
rect 110564 24160 261576 24188
rect 110564 24148 110570 24160
rect 261570 24148 261576 24160
rect 261628 24148 261634 24200
rect 9674 24080 9680 24132
rect 9732 24120 9738 24132
rect 247678 24120 247684 24132
rect 9732 24092 247684 24120
rect 9732 24080 9738 24092
rect 247678 24080 247684 24092
rect 247736 24080 247742 24132
rect 92474 22720 92480 22772
rect 92532 22760 92538 22772
rect 260098 22760 260104 22772
rect 92532 22732 260104 22760
rect 92532 22720 92538 22732
rect 260098 22720 260104 22732
rect 260156 22720 260162 22772
rect 91094 21428 91100 21480
rect 91152 21468 91158 21480
rect 253198 21468 253204 21480
rect 91152 21440 253204 21468
rect 91152 21428 91158 21440
rect 253198 21428 253204 21440
rect 253256 21428 253262 21480
rect 23474 21360 23480 21412
rect 23532 21400 23538 21412
rect 240778 21400 240784 21412
rect 23532 21372 240784 21400
rect 23532 21360 23538 21372
rect 240778 21360 240784 21372
rect 240836 21360 240842 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 39298 20652 39304 20664
rect 3476 20624 39304 20652
rect 3476 20612 3482 20624
rect 39298 20612 39304 20624
rect 39356 20612 39362 20664
rect 44266 20000 44272 20052
rect 44324 20040 44330 20052
rect 251818 20040 251824 20052
rect 44324 20012 251824 20040
rect 44324 20000 44330 20012
rect 251818 20000 251824 20012
rect 251876 20000 251882 20052
rect 4154 19932 4160 19984
rect 4212 19972 4218 19984
rect 228358 19972 228364 19984
rect 4212 19944 228364 19972
rect 4212 19932 4218 19944
rect 228358 19932 228364 19944
rect 228416 19932 228422 19984
rect 85666 18640 85672 18692
rect 85724 18680 85730 18692
rect 264238 18680 264244 18692
rect 85724 18652 264244 18680
rect 85724 18640 85730 18652
rect 264238 18640 264244 18652
rect 264296 18640 264302 18692
rect 38654 18572 38660 18624
rect 38712 18612 38718 18624
rect 244918 18612 244924 18624
rect 38712 18584 244924 18612
rect 38712 18572 38718 18584
rect 244918 18572 244924 18584
rect 244976 18572 244982 18624
rect 84194 17212 84200 17264
rect 84252 17252 84258 17264
rect 233878 17252 233884 17264
rect 84252 17224 233884 17252
rect 84252 17212 84258 17224
rect 233878 17212 233884 17224
rect 233936 17212 233942 17264
rect 120626 15920 120632 15972
rect 120684 15960 120690 15972
rect 257338 15960 257344 15972
rect 120684 15932 257344 15960
rect 120684 15920 120690 15932
rect 257338 15920 257344 15932
rect 257396 15920 257402 15972
rect 11882 15852 11888 15904
rect 11940 15892 11946 15904
rect 243630 15892 243636 15904
rect 11940 15864 243636 15892
rect 11940 15852 11946 15864
rect 243630 15852 243636 15864
rect 243688 15852 243694 15904
rect 117314 14492 117320 14544
rect 117372 14532 117378 14544
rect 229738 14532 229744 14544
rect 117372 14504 229744 14532
rect 117372 14492 117378 14504
rect 229738 14492 229744 14504
rect 229796 14492 229802 14544
rect 69106 14424 69112 14476
rect 69164 14464 69170 14476
rect 255958 14464 255964 14476
rect 69164 14436 255964 14464
rect 69164 14424 69170 14436
rect 255958 14424 255964 14436
rect 256016 14424 256022 14476
rect 114002 13132 114008 13184
rect 114060 13172 114066 13184
rect 243538 13172 243544 13184
rect 114060 13144 243544 13172
rect 114060 13132 114066 13144
rect 243538 13132 243544 13144
rect 243596 13132 243602 13184
rect 61562 13064 61568 13116
rect 61620 13104 61626 13116
rect 258718 13104 258724 13116
rect 61620 13076 258724 13104
rect 61620 13064 61626 13076
rect 258718 13064 258724 13076
rect 258776 13064 258782 13116
rect 106458 11704 106464 11756
rect 106516 11744 106522 11756
rect 239398 11744 239404 11756
rect 106516 11716 239404 11744
rect 106516 11704 106522 11716
rect 239398 11704 239404 11716
rect 239456 11704 239462 11756
rect 78582 8984 78588 9036
rect 78640 9024 78646 9036
rect 254578 9024 254584 9036
rect 78640 8996 254584 9024
rect 78640 8984 78646 8996
rect 254578 8984 254584 8996
rect 254636 8984 254642 9036
rect 51350 8916 51356 8968
rect 51408 8956 51414 8968
rect 245010 8956 245016 8968
rect 51408 8928 245016 8956
rect 51408 8916 51414 8928
rect 245010 8916 245016 8928
rect 245068 8916 245074 8968
rect 90358 7556 90364 7608
rect 90416 7596 90422 7608
rect 260190 7596 260196 7608
rect 90416 7568 260196 7596
rect 90416 7556 90422 7568
rect 260190 7556 260196 7568
rect 260248 7556 260254 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 35158 6848 35164 6860
rect 3476 6820 35164 6848
rect 3476 6808 3482 6820
rect 35158 6808 35164 6820
rect 35216 6808 35222 6860
rect 220078 6808 220084 6860
rect 220136 6848 220142 6860
rect 580166 6848 580172 6860
rect 220136 6820 580172 6848
rect 220136 6808 220142 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 72602 6196 72608 6248
rect 72660 6236 72666 6248
rect 249058 6236 249064 6248
rect 72660 6208 249064 6236
rect 72660 6196 72666 6208
rect 249058 6196 249064 6208
rect 249116 6196 249122 6248
rect 47854 6128 47860 6180
rect 47912 6168 47918 6180
rect 232498 6168 232504 6180
rect 47912 6140 232504 6168
rect 47912 6128 47918 6140
rect 232498 6128 232504 6140
rect 232556 6128 232562 6180
rect 73798 4768 73804 4820
rect 73856 4808 73862 4820
rect 238018 4808 238024 4820
rect 73856 4780 238024 4808
rect 73856 4768 73862 4780
rect 238018 4768 238024 4780
rect 238076 4768 238082 4820
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3694 3516 3700 3528
rect 2832 3488 3700 3516
rect 2832 3476 2838 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 20254 3516 20260 3528
rect 19392 3488 20260 3516
rect 19392 3476 19398 3488
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 36814 3516 36820 3528
rect 35952 3488 36820 3516
rect 35952 3476 35958 3488
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 52454 3476 52460 3528
rect 52512 3516 52518 3528
rect 53374 3516 53380 3528
rect 52512 3488 53380 3516
rect 52512 3476 52518 3488
rect 53374 3476 53380 3488
rect 53432 3476 53438 3528
rect 69014 3476 69020 3528
rect 69072 3516 69078 3528
rect 69934 3516 69940 3528
rect 69072 3488 69940 3516
rect 69072 3476 69078 3488
rect 69934 3476 69940 3488
rect 69992 3476 69998 3528
rect 95142 3476 95148 3528
rect 95200 3516 95206 3528
rect 188338 3516 188344 3528
rect 95200 3488 188344 3516
rect 95200 3476 95206 3488
rect 188338 3476 188344 3488
rect 188396 3476 188402 3528
rect 233970 3476 233976 3528
rect 234028 3516 234034 3528
rect 235810 3516 235816 3528
rect 234028 3488 235816 3516
rect 234028 3476 234034 3488
rect 235810 3476 235816 3488
rect 235868 3476 235874 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 43530 3448 43536 3460
rect 624 3420 43536 3448
rect 624 3408 630 3420
rect 43530 3408 43536 3420
rect 43588 3408 43594 3460
rect 50154 3408 50160 3460
rect 50212 3448 50218 3460
rect 106918 3448 106924 3460
rect 50212 3420 106924 3448
rect 50212 3408 50218 3420
rect 106918 3408 106924 3420
rect 106976 3408 106982 3460
rect 119890 3408 119896 3460
rect 119948 3448 119954 3460
rect 215938 3448 215944 3460
rect 119948 3420 215944 3448
rect 119948 3408 119954 3420
rect 215938 3408 215944 3420
rect 215996 3408 216002 3460
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 177948 700340 178000 700392
rect 218980 700340 219032 700392
rect 268384 700340 268436 700392
rect 494796 700340 494848 700392
rect 24308 700272 24360 700324
rect 54484 700272 54536 700324
rect 137836 700272 137888 700324
rect 178684 700272 178736 700324
rect 184848 700272 184900 700324
rect 429844 700272 429896 700324
rect 504364 700272 504416 700324
rect 527180 700272 527232 700324
rect 547144 700272 547196 700324
rect 559656 700272 559708 700324
rect 235172 699660 235224 699712
rect 240784 699660 240836 699712
rect 258724 699660 258776 699712
rect 267648 699660 267700 699712
rect 359464 699660 359516 699712
rect 364984 699660 365036 699712
rect 154120 698912 154172 698964
rect 195244 698912 195296 698964
rect 260104 698912 260156 698964
rect 283840 698912 283892 698964
rect 180708 697552 180760 697604
rect 397460 697552 397512 697604
rect 367744 696940 367796 696992
rect 580172 696940 580224 696992
rect 264244 696192 264296 696244
rect 462320 696192 462372 696244
rect 237564 694764 237616 694816
rect 477500 694764 477552 694816
rect 215668 693404 215720 693456
rect 347780 693404 347832 693456
rect 411904 683136 411956 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 71044 670692 71096 670744
rect 222844 670692 222896 670744
rect 580172 670692 580224 670744
rect 3516 656888 3568 656940
rect 249064 656888 249116 656940
rect 262864 643084 262916 643136
rect 580172 643084 580224 643136
rect 6920 632680 6972 632732
rect 188344 632680 188396 632732
rect 3516 632068 3568 632120
rect 7564 632068 7616 632120
rect 269764 630640 269816 630692
rect 580172 630640 580224 630692
rect 3516 618264 3568 618316
rect 116584 618264 116636 618316
rect 3516 605820 3568 605872
rect 97264 605820 97316 605872
rect 3332 579640 3384 579692
rect 253204 579640 253256 579692
rect 3240 565836 3292 565888
rect 108304 565836 108356 565888
rect 232504 563048 232556 563100
rect 579804 563048 579856 563100
rect 3332 553392 3384 553444
rect 14464 553392 14516 553444
rect 2964 527144 3016 527196
rect 94504 527144 94556 527196
rect 267004 524424 267056 524476
rect 580172 524424 580224 524476
rect 3516 514768 3568 514820
rect 270500 514768 270552 514820
rect 200028 510620 200080 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 251824 500964 251876 501016
rect 428464 484372 428516 484424
rect 580172 484372 580224 484424
rect 3056 474716 3108 474768
rect 251916 474716 251968 474768
rect 410524 470568 410576 470620
rect 579988 470568 580040 470620
rect 3516 462340 3568 462392
rect 166264 462340 166316 462392
rect 3148 448536 3200 448588
rect 11704 448536 11756 448588
rect 425704 430584 425756 430636
rect 580172 430584 580224 430636
rect 2780 423512 2832 423564
rect 4804 423512 4856 423564
rect 226984 418140 227036 418192
rect 580172 418140 580224 418192
rect 2872 409844 2924 409896
rect 15844 409844 15896 409896
rect 206284 404336 206336 404388
rect 580172 404336 580224 404388
rect 407764 378156 407816 378208
rect 580172 378156 580224 378208
rect 3516 371220 3568 371272
rect 173164 371220 173216 371272
rect 3148 357416 3200 357468
rect 213184 357416 213236 357468
rect 204904 351908 204956 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 224224 345040 224276 345092
rect 257436 324300 257488 324352
rect 580172 324300 580224 324352
rect 54484 320832 54536 320884
rect 215024 320832 215076 320884
rect 3332 318792 3384 318844
rect 162124 318792 162176 318844
rect 88340 318044 88392 318096
rect 234988 318044 235040 318096
rect 71780 316684 71832 316736
rect 245292 316684 245344 316736
rect 198648 315256 198700 315308
rect 331220 315256 331272 315308
rect 201500 312536 201552 312588
rect 249984 312536 250036 312588
rect 254584 311856 254636 311908
rect 580172 311856 580224 311908
rect 225328 309748 225380 309800
rect 232504 309748 232556 309800
rect 238852 309748 238904 309800
rect 412640 309748 412692 309800
rect 208584 307028 208636 307080
rect 226984 307028 227036 307080
rect 3240 304988 3292 305040
rect 251272 304988 251324 305040
rect 97264 304308 97316 304360
rect 224684 304308 224736 304360
rect 224224 304240 224276 304292
rect 249892 304240 249944 304292
rect 206008 303628 206060 303680
rect 299480 303628 299532 303680
rect 162124 302880 162176 302932
rect 246580 302880 246632 302932
rect 249064 302608 249116 302660
rect 252560 302608 252612 302660
rect 236920 302268 236972 302320
rect 276664 302268 276716 302320
rect 218888 302200 218940 302252
rect 316040 302200 316092 302252
rect 198556 301452 198608 301504
rect 206284 301452 206336 301504
rect 207940 301452 207992 301504
rect 367744 301452 367796 301504
rect 233700 300976 233752 301028
rect 273904 300976 273956 301028
rect 203432 300908 203484 300960
rect 280804 300908 280856 300960
rect 204996 300840 205048 300892
rect 582840 300840 582892 300892
rect 3424 300092 3476 300144
rect 251180 300092 251232 300144
rect 253296 300092 253348 300144
rect 504364 300092 504416 300144
rect 239496 299616 239548 299668
rect 298100 299616 298152 299668
rect 202144 299548 202196 299600
rect 268476 299548 268528 299600
rect 219532 299480 219584 299532
rect 302240 299480 302292 299532
rect 221464 299412 221516 299464
rect 222844 299412 222896 299464
rect 4804 298732 4856 298784
rect 202788 298732 202840 298784
rect 231124 298460 231176 298512
rect 259552 298460 259604 298512
rect 223396 298392 223448 298444
rect 260840 298392 260892 298444
rect 216312 298324 216364 298376
rect 263692 298324 263744 298376
rect 227904 298256 227956 298308
rect 278044 298256 278096 298308
rect 206652 298188 206704 298240
rect 299572 298188 299624 298240
rect 197268 298120 197320 298172
rect 303620 298120 303672 298172
rect 247868 296964 247920 297016
rect 267096 296964 267148 297016
rect 240140 296896 240192 296948
rect 269856 296896 269908 296948
rect 232412 296828 232464 296880
rect 265072 296828 265124 296880
rect 213736 296760 213788 296812
rect 262312 296760 262364 296812
rect 210516 296692 210568 296744
rect 583024 296692 583076 296744
rect 11704 295944 11756 295996
rect 201500 295944 201552 295996
rect 213184 295944 213236 295996
rect 228548 295944 228600 295996
rect 233056 295672 233108 295724
rect 258172 295672 258224 295724
rect 224040 295604 224092 295656
rect 264980 295604 265032 295656
rect 213092 295536 213144 295588
rect 260932 295536 260984 295588
rect 204076 295468 204128 295520
rect 204904 295468 204956 295520
rect 247224 295468 247276 295520
rect 296720 295468 296772 295520
rect 193128 295400 193180 295452
rect 226616 295400 226668 295452
rect 241428 295400 241480 295452
rect 291200 295400 291252 295452
rect 180524 295332 180576 295384
rect 214380 295332 214432 295384
rect 229192 295332 229244 295384
rect 309140 295332 309192 295384
rect 240784 294652 240836 294704
rect 255504 294652 255556 294704
rect 211804 294584 211856 294636
rect 240140 294584 240192 294636
rect 43444 294312 43496 294364
rect 227260 294312 227312 294364
rect 234344 294312 234396 294364
rect 273996 294312 274048 294364
rect 196624 294244 196676 294296
rect 222752 294244 222804 294296
rect 225972 294244 226024 294296
rect 267188 294244 267240 294296
rect 218244 294176 218296 294228
rect 244280 294176 244332 294228
rect 222108 294108 222160 294160
rect 254032 294108 254084 294160
rect 193864 294040 193916 294092
rect 231768 294040 231820 294092
rect 240140 294040 240192 294092
rect 250536 294040 250588 294092
rect 197084 293972 197136 294024
rect 204720 293972 204772 294024
rect 245936 293972 245988 294024
rect 250444 293972 250496 294024
rect 244280 293224 244332 293276
rect 258080 293224 258132 293276
rect 242716 292816 242768 292868
rect 262220 292816 262272 292868
rect 220820 292748 220872 292800
rect 250168 292748 250220 292800
rect 217600 292680 217652 292732
rect 253388 292680 253440 292732
rect 212448 292612 212500 292664
rect 253940 292612 253992 292664
rect 3424 292544 3476 292596
rect 21364 292544 21416 292596
rect 195796 292544 195848 292596
rect 205364 292544 205416 292596
rect 207296 292544 207348 292596
rect 271236 292544 271288 292596
rect 201408 292476 201460 292528
rect 204996 292476 205048 292528
rect 210240 292068 210292 292120
rect 11704 291184 11756 291236
rect 197360 291184 197412 291236
rect 241152 292068 241204 292120
rect 253756 291320 253808 291372
rect 259460 291320 259512 291372
rect 255412 291252 255464 291304
rect 256700 291184 256752 291236
rect 253756 291116 253808 291168
rect 407764 291116 407816 291168
rect 188988 289824 189040 289876
rect 197360 289824 197412 289876
rect 195244 289756 195296 289808
rect 197728 289756 197780 289808
rect 253756 288464 253808 288516
rect 272524 288464 272576 288516
rect 186228 288396 186280 288448
rect 197360 288396 197412 288448
rect 252928 288396 252980 288448
rect 296812 288396 296864 288448
rect 190368 287104 190420 287156
rect 197360 287104 197412 287156
rect 182088 287036 182140 287088
rect 197452 287036 197504 287088
rect 253756 287036 253808 287088
rect 305644 287036 305696 287088
rect 71044 286968 71096 287020
rect 197360 286968 197412 287020
rect 253756 285676 253808 285728
rect 381544 285676 381596 285728
rect 253848 285608 253900 285660
rect 410524 285608 410576 285660
rect 3516 284928 3568 284980
rect 196624 284928 196676 284980
rect 188896 284316 188948 284368
rect 197360 284316 197412 284368
rect 253756 282888 253808 282940
rect 278136 282888 278188 282940
rect 250444 282140 250496 282192
rect 580264 282140 580316 282192
rect 252560 280304 252612 280356
rect 255596 280304 255648 280356
rect 183468 280168 183520 280220
rect 197360 280168 197412 280220
rect 253756 280168 253808 280220
rect 295340 280168 295392 280220
rect 35164 278740 35216 278792
rect 197360 278740 197412 278792
rect 253388 277992 253440 278044
rect 263600 277992 263652 278044
rect 190092 277448 190144 277500
rect 197452 277448 197504 277500
rect 187424 277380 187476 277432
rect 197360 277380 197412 277432
rect 253848 277380 253900 277432
rect 283104 277380 283156 277432
rect 251916 276972 251968 277024
rect 252560 276972 252612 277024
rect 195888 276088 195940 276140
rect 197728 276088 197780 276140
rect 190276 276020 190328 276072
rect 197360 276020 197412 276072
rect 253296 276020 253348 276072
rect 566464 276020 566516 276072
rect 187516 274728 187568 274780
rect 197360 274728 197412 274780
rect 184756 274660 184808 274712
rect 197452 274660 197504 274712
rect 253296 274660 253348 274712
rect 385684 274660 385736 274712
rect 116584 274592 116636 274644
rect 197360 274592 197412 274644
rect 252652 274252 252704 274304
rect 254584 274252 254636 274304
rect 253756 273912 253808 273964
rect 283012 273912 283064 273964
rect 253480 272484 253532 272536
rect 287060 272484 287112 272536
rect 252652 272144 252704 272196
rect 254216 272144 254268 272196
rect 251824 271872 251876 271924
rect 252652 271872 252704 271924
rect 574744 271872 574796 271924
rect 580172 271872 580224 271924
rect 169760 271804 169812 271856
rect 197360 271804 197412 271856
rect 250536 271124 250588 271176
rect 580356 271124 580408 271176
rect 192852 270512 192904 270564
rect 197452 270512 197504 270564
rect 192944 269152 192996 269204
rect 197452 269152 197504 269204
rect 186136 269084 186188 269136
rect 197360 269084 197412 269136
rect 18604 267724 18656 267776
rect 197360 267724 197412 267776
rect 253204 267724 253256 267776
rect 271144 267724 271196 267776
rect 108304 267656 108356 267708
rect 197452 267656 197504 267708
rect 188344 267588 188396 267640
rect 197360 267588 197412 267640
rect 253756 266432 253808 266484
rect 276756 266432 276808 266484
rect 253296 266364 253348 266416
rect 290096 266364 290148 266416
rect 7564 266296 7616 266348
rect 197360 266296 197412 266348
rect 253756 265004 253808 265056
rect 267280 265004 267332 265056
rect 187608 264936 187660 264988
rect 197452 264936 197504 264988
rect 253848 264936 253900 264988
rect 303712 264936 303764 264988
rect 253756 264868 253808 264920
rect 428464 264868 428516 264920
rect 188712 263644 188764 263696
rect 197360 263644 197412 263696
rect 17224 263576 17276 263628
rect 197452 263576 197504 263628
rect 14464 263508 14516 263560
rect 197360 263508 197412 263560
rect 191656 262216 191708 262268
rect 197360 262216 197412 262268
rect 253756 262216 253808 262268
rect 300860 262216 300912 262268
rect 195704 260924 195756 260976
rect 197544 260924 197596 260976
rect 172428 260856 172480 260908
rect 197452 260856 197504 260908
rect 253388 260856 253440 260908
rect 293960 260856 294012 260908
rect 94504 260788 94556 260840
rect 197360 260788 197412 260840
rect 253204 259496 253256 259548
rect 256792 259496 256844 259548
rect 175188 259428 175240 259480
rect 197360 259428 197412 259480
rect 252836 259428 252888 259480
rect 382924 259428 382976 259480
rect 271236 259360 271288 259412
rect 579620 259360 579672 259412
rect 252560 259020 252612 259072
rect 255504 259020 255556 259072
rect 191748 258272 191800 258324
rect 197452 258272 197504 258324
rect 188804 258068 188856 258120
rect 197360 258068 197412 258120
rect 253848 258068 253900 258120
rect 276848 258068 276900 258120
rect 250352 258000 250404 258052
rect 253756 258000 253808 258052
rect 253020 257524 253072 257576
rect 257436 257524 257488 257576
rect 184664 256776 184716 256828
rect 197360 256776 197412 256828
rect 14464 256708 14516 256760
rect 197452 256708 197504 256760
rect 253112 256640 253164 256692
rect 582380 256640 582432 256692
rect 253756 256572 253808 256624
rect 425704 256572 425756 256624
rect 177856 255280 177908 255332
rect 197452 255280 197504 255332
rect 184848 255212 184900 255264
rect 197360 255212 197412 255264
rect 253020 253988 253072 254040
rect 256884 253988 256936 254040
rect 3148 253920 3200 253972
rect 169024 253920 169076 253972
rect 193036 253920 193088 253972
rect 197360 253920 197412 253972
rect 253756 253920 253808 253972
rect 271236 253920 271288 253972
rect 25504 252560 25556 252612
rect 197360 252560 197412 252612
rect 253848 252560 253900 252612
rect 305000 252560 305052 252612
rect 253756 252492 253808 252544
rect 411904 252492 411956 252544
rect 181996 251268 182048 251320
rect 197452 251268 197504 251320
rect 180616 251200 180668 251252
rect 197360 251200 197412 251252
rect 187332 250452 187384 250504
rect 198096 250452 198148 250504
rect 253480 250452 253532 250504
rect 284300 250452 284352 250504
rect 253388 249976 253440 250028
rect 259644 249976 259696 250028
rect 191564 249772 191616 249824
rect 197452 249772 197504 249824
rect 178684 249704 178736 249756
rect 197360 249704 197412 249756
rect 253756 249704 253808 249756
rect 267004 249704 267056 249756
rect 194508 248684 194560 248736
rect 197360 248684 197412 248736
rect 253756 248412 253808 248464
rect 306380 248412 306432 248464
rect 180708 248344 180760 248396
rect 197452 248344 197504 248396
rect 253848 248344 253900 248396
rect 270500 248344 270552 248396
rect 194416 247052 194468 247104
rect 197544 247052 197596 247104
rect 253756 247052 253808 247104
rect 263784 247052 263836 247104
rect 15844 246984 15896 247036
rect 197360 246984 197412 247036
rect 253756 245624 253808 245676
rect 298192 245624 298244 245676
rect 253848 245556 253900 245608
rect 264244 245556 264296 245608
rect 3608 244876 3660 244928
rect 191104 244876 191156 244928
rect 195612 244264 195664 244316
rect 197452 244264 197504 244316
rect 253756 244264 253808 244316
rect 292856 244264 292908 244316
rect 21364 244196 21416 244248
rect 197360 244196 197412 244248
rect 253388 244196 253440 244248
rect 579896 244264 579948 244316
rect 253756 242972 253808 243024
rect 260104 242972 260156 243024
rect 192852 242836 192904 242888
rect 198740 242836 198792 242888
rect 253756 242836 253808 242888
rect 547144 242836 547196 242888
rect 252560 241544 252612 241596
rect 255504 241544 255556 241596
rect 190184 241476 190236 241528
rect 197360 241476 197412 241528
rect 3056 240116 3108 240168
rect 191840 240116 191892 240168
rect 249064 240116 249116 240168
rect 250260 240116 250312 240168
rect 253756 240116 253808 240168
rect 311900 240116 311952 240168
rect 206016 240048 206068 240100
rect 582472 240048 582524 240100
rect 169024 239980 169076 240032
rect 242716 239980 242768 240032
rect 244012 239980 244064 240032
rect 268384 239980 268436 240032
rect 200764 239912 200816 239964
rect 206376 239912 206428 239964
rect 236920 239912 236972 239964
rect 258724 239912 258776 239964
rect 190552 239844 190604 239896
rect 212448 239844 212500 239896
rect 195796 239776 195848 239828
rect 238760 239776 238812 239828
rect 249248 239776 249300 239828
rect 254124 239776 254176 239828
rect 198740 239368 198792 239420
rect 215944 239368 215996 239420
rect 245016 239368 245068 239420
rect 252744 239368 252796 239420
rect 246304 238756 246356 238808
rect 250168 238756 250220 238808
rect 177948 238688 178000 238740
rect 211804 238688 211856 238740
rect 222108 238688 222160 238740
rect 583116 238688 583168 238740
rect 191104 238620 191156 238672
rect 216956 238620 217008 238672
rect 221464 238620 221516 238672
rect 574744 238620 574796 238672
rect 228548 238552 228600 238604
rect 359464 238552 359516 238604
rect 191840 238484 191892 238536
rect 233700 238484 233752 238536
rect 247224 238484 247276 238536
rect 269764 238484 269816 238536
rect 173164 238416 173216 238468
rect 229192 238416 229244 238468
rect 235632 238076 235684 238128
rect 267004 238076 267056 238128
rect 218888 238008 218940 238060
rect 300952 238008 301004 238060
rect 202788 237804 202840 237856
rect 205548 237804 205600 237856
rect 200212 237396 200264 237448
rect 206284 237396 206336 237448
rect 233056 237396 233108 237448
rect 237380 237396 237432 237448
rect 245292 237328 245344 237380
rect 582564 237328 582616 237380
rect 244924 236716 244976 236768
rect 251088 236716 251140 236768
rect 199844 236648 199896 236700
rect 281632 236648 281684 236700
rect 205548 235900 205600 235952
rect 582932 235900 582984 235952
rect 166264 235832 166316 235884
rect 244648 235832 244700 235884
rect 242164 235356 242216 235408
rect 252836 235356 252888 235408
rect 243544 235288 243596 235340
rect 265072 235288 265124 235340
rect 247868 235220 247920 235272
rect 322204 235220 322256 235272
rect 237564 234540 237616 234592
rect 542360 234540 542412 234592
rect 253848 233928 253900 233980
rect 255504 233928 255556 233980
rect 188712 233860 188764 233912
rect 306472 233860 306524 233912
rect 231124 233180 231176 233232
rect 233240 233180 233292 233232
rect 566464 233180 566516 233232
rect 580172 233180 580224 233232
rect 249800 232636 249852 232688
rect 287152 232636 287204 232688
rect 191104 232568 191156 232620
rect 254216 232568 254268 232620
rect 206652 232500 206704 232552
rect 302884 232500 302936 232552
rect 200856 231072 200908 231124
rect 284484 231072 284536 231124
rect 190092 228420 190144 228472
rect 269764 228420 269816 228472
rect 21364 228352 21416 228404
rect 213736 228352 213788 228404
rect 230480 225700 230532 225752
rect 231860 225700 231912 225752
rect 196992 225564 197044 225616
rect 230480 225564 230532 225616
rect 235264 225564 235316 225616
rect 252652 225564 252704 225616
rect 200028 224204 200080 224256
rect 230572 224204 230624 224256
rect 231768 223524 231820 223576
rect 233332 223524 233384 223576
rect 199936 222844 199988 222896
rect 230664 222844 230716 222896
rect 7564 220056 7616 220108
rect 240784 220056 240836 220108
rect 4804 218696 4856 218748
rect 240140 218696 240192 218748
rect 3332 215228 3384 215280
rect 17224 215228 17276 215280
rect 211160 211760 211212 211812
rect 287244 211760 287296 211812
rect 257344 206932 257396 206984
rect 579896 206932 579948 206984
rect 198556 206252 198608 206304
rect 285772 206252 285824 206304
rect 195704 204892 195756 204944
rect 281724 204892 281776 204944
rect 3056 202784 3108 202836
rect 259644 202784 259696 202836
rect 229836 202104 229888 202156
rect 284576 202104 284628 202156
rect 215024 200744 215076 200796
rect 287336 200744 287388 200796
rect 202144 196596 202196 196648
rect 280160 196596 280212 196648
rect 181996 195236 182048 195288
rect 292764 195236 292816 195288
rect 234344 193808 234396 193860
rect 305092 193808 305144 193860
rect 188896 193128 188948 193180
rect 580172 193128 580224 193180
rect 224040 191156 224092 191208
rect 233424 191156 233476 191208
rect 217600 191088 217652 191140
rect 299664 191088 299716 191140
rect 172428 189864 172480 189916
rect 288624 189864 288676 189916
rect 175188 189796 175240 189848
rect 295524 189796 295576 189848
rect 177856 189728 177908 189780
rect 299756 189728 299808 189780
rect 245936 188436 245988 188488
rect 284392 188436 284444 188488
rect 210516 188368 210568 188420
rect 276940 188368 276992 188420
rect 184664 188300 184716 188352
rect 296904 188300 296956 188352
rect 236276 187008 236328 187060
rect 292672 187008 292724 187060
rect 238852 186940 238904 186992
rect 303804 186940 303856 186992
rect 190276 185852 190328 185904
rect 236000 185852 236052 185904
rect 186228 185784 186280 185836
rect 240232 185784 240284 185836
rect 201500 185716 201552 185768
rect 231952 185716 232004 185768
rect 232412 185716 232464 185768
rect 294144 185716 294196 185768
rect 184756 185648 184808 185700
rect 291384 185648 291436 185700
rect 3516 185580 3568 185632
rect 193864 185580 193916 185632
rect 223396 185580 223448 185632
rect 285864 185580 285916 185632
rect 197268 184288 197320 184340
rect 230756 184288 230808 184340
rect 278136 184288 278188 184340
rect 307760 184288 307812 184340
rect 227904 184220 227956 184272
rect 288440 184220 288492 184272
rect 225328 184152 225380 184204
rect 289912 184152 289964 184204
rect 100668 183540 100720 183592
rect 209044 183540 209096 183592
rect 220176 183132 220228 183184
rect 232136 183132 232188 183184
rect 191656 183064 191708 183116
rect 234620 183064 234672 183116
rect 188988 182996 189040 183048
rect 244372 182996 244424 183048
rect 187332 182928 187384 182980
rect 247040 182928 247092 182980
rect 214380 182860 214432 182912
rect 298284 182860 298336 182912
rect 203432 182792 203484 182844
rect 296996 182792 297048 182844
rect 127072 182384 127124 182436
rect 170588 182384 170640 182436
rect 108120 182316 108172 182368
rect 169024 182316 169076 182368
rect 105912 182248 105964 182300
rect 167644 182248 167696 182300
rect 130752 182180 130804 182232
rect 204904 182180 204956 182232
rect 215668 181432 215720 181484
rect 232044 181432 232096 181484
rect 243360 181432 243412 181484
rect 295432 181432 295484 181484
rect 132408 181092 132460 181144
rect 166540 181092 166592 181144
rect 124956 181024 125008 181076
rect 167828 181024 167880 181076
rect 103336 180956 103388 181008
rect 166264 180956 166316 181008
rect 114468 180888 114520 180940
rect 178684 180888 178736 180940
rect 119528 180820 119580 180872
rect 213276 180820 213328 180872
rect 180524 180412 180576 180464
rect 227628 180412 227680 180464
rect 190184 180344 190236 180396
rect 237472 180344 237524 180396
rect 187424 180276 187476 180328
rect 234712 180276 234764 180328
rect 276756 180276 276808 180328
rect 288716 180276 288768 180328
rect 226616 180208 226668 180260
rect 280344 180208 280396 180260
rect 188804 180140 188856 180192
rect 242992 180140 243044 180192
rect 272524 180140 272576 180192
rect 301044 180140 301096 180192
rect 224684 180072 224736 180124
rect 291292 180072 291344 180124
rect 123760 179596 123812 179648
rect 169208 179596 169260 179648
rect 97540 179528 97592 179580
rect 173164 179528 173216 179580
rect 129464 179460 129516 179512
rect 214196 179460 214248 179512
rect 114376 179392 114428 179444
rect 211804 179392 211856 179444
rect 218244 178916 218296 178968
rect 229100 178916 229152 178968
rect 208584 178848 208636 178900
rect 238852 178848 238904 178900
rect 273904 178848 273956 178900
rect 295616 178848 295668 178900
rect 191564 178780 191616 178832
rect 244280 178780 244332 178832
rect 271144 178780 271196 178832
rect 294052 178780 294104 178832
rect 206284 178712 206336 178764
rect 291476 178712 291528 178764
rect 204076 178644 204128 178696
rect 301136 178644 301188 178696
rect 118424 178304 118476 178356
rect 166356 178304 166408 178356
rect 110696 178236 110748 178288
rect 169116 178236 169168 178288
rect 112260 178168 112312 178220
rect 177304 178168 177356 178220
rect 133144 178100 133196 178152
rect 214012 178100 214064 178152
rect 109592 178032 109644 178084
rect 213184 178032 213236 178084
rect 227260 177964 227312 178016
rect 229192 177964 229244 178016
rect 268476 177964 268528 178016
rect 296628 177964 296680 178016
rect 222752 177488 222804 177540
rect 236092 177488 236144 177540
rect 220820 177420 220872 177472
rect 238760 177420 238812 177472
rect 271236 177420 271288 177472
rect 288532 177420 288584 177472
rect 194416 177352 194468 177404
rect 236276 177352 236328 177404
rect 276848 177352 276900 177404
rect 302332 177352 302384 177404
rect 195612 177284 195664 177336
rect 292580 177284 292632 177336
rect 128176 177012 128228 177064
rect 214104 177012 214156 177064
rect 107016 176944 107068 176996
rect 165344 176944 165396 176996
rect 148232 176876 148284 176928
rect 214564 176876 214616 176928
rect 104624 176808 104676 176860
rect 170496 176808 170548 176860
rect 125876 176740 125928 176792
rect 198004 176740 198056 176792
rect 136088 176672 136140 176724
rect 158996 176672 159048 176724
rect 165436 176672 165488 176724
rect 213920 176604 213972 176656
rect 134432 176196 134484 176248
rect 165528 176196 165580 176248
rect 121920 176128 121972 176180
rect 166448 176128 166500 176180
rect 194508 176128 194560 176180
rect 242900 176128 242952 176180
rect 276664 176128 276716 176180
rect 279332 176128 279384 176180
rect 116952 176060 117004 176112
rect 169300 176060 169352 176112
rect 187516 176060 187568 176112
rect 236184 176060 236236 176112
rect 278044 176060 278096 176112
rect 290004 176060 290056 176112
rect 120816 175992 120868 176044
rect 180064 175992 180116 176044
rect 183468 175992 183520 176044
rect 237564 175992 237616 176044
rect 276940 175992 276992 176044
rect 289820 175992 289872 176044
rect 115756 175924 115808 175976
rect 211896 175924 211948 175976
rect 238208 175924 238260 175976
rect 280252 175924 280304 175976
rect 235356 175244 235408 175296
rect 265808 175244 265860 175296
rect 165528 175176 165580 175228
rect 213920 175176 213972 175228
rect 231124 175176 231176 175228
rect 250444 175176 250496 175228
rect 231768 175108 231820 175160
rect 245016 175108 245068 175160
rect 165436 174496 165488 174548
rect 214656 174496 214708 174548
rect 256056 174020 256108 174072
rect 265348 174020 265400 174072
rect 247868 173952 247920 174004
rect 265808 173952 265860 174004
rect 238024 173884 238076 173936
rect 265624 173884 265676 173936
rect 166540 173816 166592 173868
rect 213920 173816 213972 173868
rect 231216 173816 231268 173868
rect 265256 173816 265308 173868
rect 204904 173748 204956 173800
rect 214012 173748 214064 173800
rect 231768 173748 231820 173800
rect 252008 173748 252060 173800
rect 231676 173680 231728 173732
rect 236000 173680 236052 173732
rect 254676 173136 254728 173188
rect 265900 173136 265952 173188
rect 243636 172592 243688 172644
rect 265900 172592 265952 172644
rect 236828 172524 236880 172576
rect 265808 172524 265860 172576
rect 231768 172456 231820 172508
rect 251272 172456 251324 172508
rect 231676 172388 231728 172440
rect 251364 172388 251416 172440
rect 231676 171708 231728 171760
rect 235264 171708 235316 171760
rect 258816 171504 258868 171556
rect 265348 171504 265400 171556
rect 251824 171164 251876 171216
rect 265900 171164 265952 171216
rect 247684 171096 247736 171148
rect 265808 171096 265860 171148
rect 170588 171028 170640 171080
rect 213920 171028 213972 171080
rect 231768 171028 231820 171080
rect 263692 171028 263744 171080
rect 282736 171028 282788 171080
rect 296996 171028 297048 171080
rect 198004 170960 198056 171012
rect 214012 170960 214064 171012
rect 282828 170960 282880 171012
rect 290004 170960 290056 171012
rect 231308 170552 231360 170604
rect 236184 170552 236236 170604
rect 231768 170484 231820 170536
rect 236276 170484 236328 170536
rect 236644 170348 236696 170400
rect 265716 170348 265768 170400
rect 168012 169736 168064 169788
rect 170404 169736 170456 169788
rect 246396 169736 246448 169788
rect 265348 169736 265400 169788
rect 167828 169668 167880 169720
rect 213920 169668 213972 169720
rect 231768 169668 231820 169720
rect 258080 169668 258132 169720
rect 282828 169668 282880 169720
rect 289820 169668 289872 169720
rect 169208 169600 169260 169652
rect 214012 169600 214064 169652
rect 231676 169532 231728 169584
rect 237380 169532 237432 169584
rect 240876 168512 240928 168564
rect 245016 168444 245068 168496
rect 246580 168444 246632 168496
rect 260288 168512 260340 168564
rect 265624 168512 265676 168564
rect 265808 168444 265860 168496
rect 235540 168376 235592 168428
rect 264428 168376 264480 168428
rect 166448 168308 166500 168360
rect 213920 168308 213972 168360
rect 231768 168308 231820 168360
rect 260932 168308 260984 168360
rect 282460 168308 282512 168360
rect 292580 168308 292632 168360
rect 180064 168240 180116 168292
rect 214012 168240 214064 168292
rect 231676 168240 231728 168292
rect 254032 168240 254084 168292
rect 231584 168172 231636 168224
rect 250076 168172 250128 168224
rect 246488 167628 246540 167680
rect 265440 167628 265492 167680
rect 262956 167084 263008 167136
rect 265164 167084 265216 167136
rect 239680 167016 239732 167068
rect 265808 167016 265860 167068
rect 231768 166948 231820 167000
rect 244924 166948 244976 167000
rect 282092 166948 282144 167000
rect 294236 166948 294288 167000
rect 382924 166948 382976 167000
rect 580172 166948 580224 167000
rect 169300 166880 169352 166932
rect 214012 166880 214064 166932
rect 231124 166880 231176 166932
rect 234620 166880 234672 166932
rect 166356 166812 166408 166864
rect 213920 166812 213972 166864
rect 240784 166268 240836 166320
rect 265348 166268 265400 166320
rect 231492 166064 231544 166116
rect 236092 166064 236144 166116
rect 261484 165656 261536 165708
rect 265808 165656 265860 165708
rect 245108 165588 245160 165640
rect 265716 165588 265768 165640
rect 178684 165520 178736 165572
rect 213920 165520 213972 165572
rect 231768 165520 231820 165572
rect 255412 165520 255464 165572
rect 282000 165520 282052 165572
rect 294144 165520 294196 165572
rect 211896 165452 211948 165504
rect 214656 165452 214708 165504
rect 231308 165452 231360 165504
rect 234712 165452 234764 165504
rect 282828 165452 282880 165504
rect 291476 165452 291528 165504
rect 236920 164840 236972 164892
rect 261392 164840 261444 164892
rect 230664 164568 230716 164620
rect 232136 164568 232188 164620
rect 257436 164296 257488 164348
rect 265808 164296 265860 164348
rect 242256 164228 242308 164280
rect 265440 164228 265492 164280
rect 177304 164160 177356 164212
rect 213920 164160 213972 164212
rect 231676 164160 231728 164212
rect 242164 164160 242216 164212
rect 282828 164160 282880 164212
rect 295524 164160 295576 164212
rect 211804 164092 211856 164144
rect 214472 164092 214524 164144
rect 282092 163208 282144 163260
rect 288624 163208 288676 163260
rect 250628 163004 250680 163056
rect 265532 163004 265584 163056
rect 242348 162936 242400 162988
rect 265348 162936 265400 162988
rect 235264 162868 235316 162920
rect 265900 162868 265952 162920
rect 169116 162800 169168 162852
rect 213920 162800 213972 162852
rect 231768 162800 231820 162852
rect 249984 162800 250036 162852
rect 282092 162800 282144 162852
rect 298100 162800 298152 162852
rect 231676 162732 231728 162784
rect 238852 162732 238904 162784
rect 282828 162732 282880 162784
rect 292856 162732 292908 162784
rect 260196 162120 260248 162172
rect 265808 162120 265860 162172
rect 231768 161984 231820 162036
rect 237564 161984 237616 162036
rect 249524 161508 249576 161560
rect 265348 161508 265400 161560
rect 238300 161440 238352 161492
rect 265808 161440 265860 161492
rect 169024 161372 169076 161424
rect 213920 161372 213972 161424
rect 231768 161372 231820 161424
rect 262312 161372 262364 161424
rect 282828 161372 282880 161424
rect 291200 161372 291252 161424
rect 231400 161304 231452 161356
rect 245016 161304 245068 161356
rect 167736 160692 167788 160744
rect 214104 160692 214156 160744
rect 281540 160624 281592 160676
rect 283196 160624 283248 160676
rect 255964 160216 256016 160268
rect 265624 160216 265676 160268
rect 244924 160148 244976 160200
rect 265348 160148 265400 160200
rect 239496 160080 239548 160132
rect 265808 160080 265860 160132
rect 167644 160012 167696 160064
rect 213920 160012 213972 160064
rect 231492 160012 231544 160064
rect 249248 160012 249300 160064
rect 281540 160012 281592 160064
rect 284484 160012 284536 160064
rect 170496 159944 170548 159996
rect 214012 159944 214064 159996
rect 231768 159944 231820 159996
rect 240232 159944 240284 159996
rect 263048 158856 263100 158908
rect 265624 158856 265676 158908
rect 249432 158788 249484 158840
rect 265348 158788 265400 158840
rect 242164 158720 242216 158772
rect 265808 158720 265860 158772
rect 166264 158652 166316 158704
rect 213920 158652 213972 158704
rect 231768 158652 231820 158704
rect 260840 158652 260892 158704
rect 282736 158652 282788 158704
rect 295616 158652 295668 158704
rect 282828 158584 282880 158636
rect 288716 158584 288768 158636
rect 254768 157972 254820 158024
rect 265992 157972 266044 158024
rect 236736 157428 236788 157480
rect 265624 157428 265676 157480
rect 232504 157360 232556 157412
rect 265532 157360 265584 157412
rect 209044 157292 209096 157344
rect 213920 157292 213972 157344
rect 231768 157292 231820 157344
rect 259552 157292 259604 157344
rect 231676 157224 231728 157276
rect 256792 157224 256844 157276
rect 281724 156544 281776 156596
rect 284576 156544 284628 156596
rect 253204 156068 253256 156120
rect 265900 156068 265952 156120
rect 246672 156000 246724 156052
rect 265532 156000 265584 156052
rect 238208 155932 238260 155984
rect 265808 155932 265860 155984
rect 173164 155864 173216 155916
rect 213920 155864 213972 155916
rect 231124 155796 231176 155848
rect 233240 155796 233292 155848
rect 231768 155728 231820 155780
rect 246304 155728 246356 155780
rect 258908 155524 258960 155576
rect 261668 155524 261720 155576
rect 230572 155388 230624 155440
rect 232044 155388 232096 155440
rect 250720 154640 250772 154692
rect 265808 154640 265860 154692
rect 239588 154572 239640 154624
rect 265716 154572 265768 154624
rect 281724 154504 281776 154556
rect 300952 154504 301004 154556
rect 252192 153824 252244 153876
rect 265256 153824 265308 153876
rect 282828 153416 282880 153468
rect 287244 153416 287296 153468
rect 180064 153280 180116 153332
rect 213920 153280 213972 153332
rect 241152 153280 241204 153332
rect 265900 153280 265952 153332
rect 169024 153212 169076 153264
rect 214012 153212 214064 153264
rect 234160 153212 234212 153264
rect 265808 153212 265860 153264
rect 231768 153144 231820 153196
rect 262220 153144 262272 153196
rect 282736 153144 282788 153196
rect 305000 153144 305052 153196
rect 381544 153144 381596 153196
rect 579804 153144 579856 153196
rect 231676 153076 231728 153128
rect 244372 153076 244424 153128
rect 234528 152464 234580 152516
rect 242072 152464 242124 152516
rect 245200 152464 245252 152516
rect 265992 152464 266044 152516
rect 241060 151920 241112 151972
rect 265716 151920 265768 151972
rect 196624 151852 196676 151904
rect 213920 151852 213972 151904
rect 177396 151784 177448 151836
rect 214012 151784 214064 151836
rect 261760 151784 261812 151836
rect 265808 151784 265860 151836
rect 282828 151716 282880 151768
rect 301136 151716 301188 151768
rect 231676 151648 231728 151700
rect 234528 151648 234580 151700
rect 231768 151580 231820 151632
rect 238760 151580 238812 151632
rect 258724 150560 258776 150612
rect 265900 150560 265952 150612
rect 198096 150492 198148 150544
rect 213920 150492 213972 150544
rect 254860 150492 254912 150544
rect 265992 150492 266044 150544
rect 170496 150424 170548 150476
rect 214012 150424 214064 150476
rect 246580 150424 246632 150476
rect 265808 150424 265860 150476
rect 3424 150356 3476 150408
rect 11704 150356 11756 150408
rect 170404 150356 170456 150408
rect 213920 150356 213972 150408
rect 282828 150356 282880 150408
rect 291384 150356 291436 150408
rect 231676 150288 231728 150340
rect 249064 150288 249116 150340
rect 231768 150220 231820 150272
rect 253940 150220 253992 150272
rect 230940 150016 230992 150068
rect 233424 150016 233476 150068
rect 231216 149676 231268 149728
rect 245108 149676 245160 149728
rect 281540 149608 281592 149660
rect 284300 149608 284352 149660
rect 263140 149200 263192 149252
rect 265348 149200 265400 149252
rect 249340 149132 249392 149184
rect 265808 149132 265860 149184
rect 245016 149064 245068 149116
rect 265900 149064 265952 149116
rect 231768 148996 231820 149048
rect 243544 148996 243596 149048
rect 282828 148996 282880 149048
rect 290096 148996 290148 149048
rect 282276 148588 282328 148640
rect 287336 148588 287388 148640
rect 232780 148316 232832 148368
rect 266084 148316 266136 148368
rect 259000 147704 259052 147756
rect 265808 147704 265860 147756
rect 166264 147636 166316 147688
rect 213920 147636 213972 147688
rect 235448 147636 235500 147688
rect 265440 147636 265492 147688
rect 231768 147568 231820 147620
rect 263600 147568 263652 147620
rect 281724 147568 281776 147620
rect 316040 147568 316092 147620
rect 230940 147024 230992 147076
rect 233332 147024 233384 147076
rect 232596 146888 232648 146940
rect 265164 146888 265216 146940
rect 234068 146344 234120 146396
rect 265808 146344 265860 146396
rect 174544 146276 174596 146328
rect 213920 146276 213972 146328
rect 232688 146276 232740 146328
rect 265532 146276 265584 146328
rect 231768 146208 231820 146260
rect 244280 146208 244332 146260
rect 282000 146208 282052 146260
rect 299756 146208 299808 146260
rect 231676 146140 231728 146192
rect 242992 146140 243044 146192
rect 282828 146140 282880 146192
rect 296720 146140 296772 146192
rect 231032 146072 231084 146124
rect 237472 146072 237524 146124
rect 238392 145528 238444 145580
rect 261576 145528 261628 145580
rect 233976 145052 234028 145104
rect 265808 145052 265860 145104
rect 252100 144984 252152 145036
rect 265532 144984 265584 145036
rect 178684 144916 178736 144968
rect 213920 144916 213972 144968
rect 231584 144848 231636 144900
rect 261852 144848 261904 144900
rect 265716 144848 265768 144900
rect 263784 144780 263836 144832
rect 282552 144780 282604 144832
rect 285772 144780 285824 144832
rect 282828 143692 282880 143744
rect 287060 143692 287112 143744
rect 177304 143624 177356 143676
rect 214012 143624 214064 143676
rect 250812 143624 250864 143676
rect 265440 143624 265492 143676
rect 171876 143556 171928 143608
rect 213920 143556 213972 143608
rect 229928 143556 229980 143608
rect 265808 143556 265860 143608
rect 231676 143488 231728 143540
rect 259460 143488 259512 143540
rect 281632 143488 281684 143540
rect 301044 143488 301096 143540
rect 231768 143420 231820 143472
rect 251180 143420 251232 143472
rect 231124 143352 231176 143404
rect 233792 143352 233844 143404
rect 233884 142808 233936 142860
rect 265624 142808 265676 142860
rect 260380 142332 260432 142384
rect 264336 142332 264388 142384
rect 243728 142264 243780 142316
rect 265348 142264 265400 142316
rect 188344 142128 188396 142180
rect 213920 142128 213972 142180
rect 231768 142060 231820 142112
rect 255596 142060 255648 142112
rect 282828 142060 282880 142112
rect 303712 142060 303764 142112
rect 231308 141448 231360 141500
rect 251824 141448 251876 141500
rect 245292 141380 245344 141432
rect 266084 141380 266136 141432
rect 175924 140836 175976 140888
rect 213920 140836 213972 140888
rect 170404 140768 170456 140820
rect 214012 140768 214064 140820
rect 256332 140768 256384 140820
rect 265808 140768 265860 140820
rect 231676 140700 231728 140752
rect 256700 140700 256752 140752
rect 281908 140700 281960 140752
rect 296812 140700 296864 140752
rect 231768 140632 231820 140684
rect 247040 140632 247092 140684
rect 210424 139408 210476 139460
rect 213920 139408 213972 139460
rect 257344 139408 257396 139460
rect 265440 139408 265492 139460
rect 282828 139340 282880 139392
rect 313280 139340 313332 139392
rect 282736 139272 282788 139324
rect 292764 139272 292816 139324
rect 231216 138660 231268 138712
rect 244924 138660 244976 138712
rect 247776 138116 247828 138168
rect 265624 138116 265676 138168
rect 202144 138048 202196 138100
rect 213920 138048 213972 138100
rect 243544 138048 243596 138100
rect 265164 138048 265216 138100
rect 171968 137980 172020 138032
rect 214012 137980 214064 138032
rect 229744 137980 229796 138032
rect 265440 137980 265492 138032
rect 3424 137912 3476 137964
rect 14464 137912 14516 137964
rect 231400 137912 231452 137964
rect 262404 137912 262456 137964
rect 282184 137912 282236 137964
rect 298376 137912 298428 137964
rect 231768 137844 231820 137896
rect 242900 137844 242952 137896
rect 282828 137844 282880 137896
rect 293960 137844 294012 137896
rect 231584 137232 231636 137284
rect 243636 137232 243688 137284
rect 249248 136688 249300 136740
rect 265532 136688 265584 136740
rect 206376 136620 206428 136672
rect 213920 136620 213972 136672
rect 239404 136620 239456 136672
rect 265624 136620 265676 136672
rect 231400 136552 231452 136604
rect 256056 136552 256108 136604
rect 231768 136484 231820 136536
rect 247868 136484 247920 136536
rect 260104 135464 260156 135516
rect 265348 135464 265400 135516
rect 261484 135396 261536 135448
rect 266084 135396 266136 135448
rect 253388 135328 253440 135380
rect 265624 135328 265676 135380
rect 238116 135260 238168 135312
rect 265900 135260 265952 135312
rect 231492 135192 231544 135244
rect 254676 135192 254728 135244
rect 231032 135056 231084 135108
rect 236644 135056 236696 135108
rect 173348 134512 173400 134564
rect 214840 134512 214892 134564
rect 254584 134036 254636 134088
rect 265900 134036 265952 134088
rect 253296 133968 253348 134020
rect 265532 133968 265584 134020
rect 204904 133900 204956 133952
rect 213920 133900 213972 133952
rect 229836 133900 229888 133952
rect 265900 133900 265952 133952
rect 231676 133832 231728 133884
rect 258816 133832 258868 133884
rect 282828 133832 282880 133884
rect 311900 133832 311952 133884
rect 230940 133764 230992 133816
rect 236828 133764 236880 133816
rect 262864 132608 262916 132660
rect 265624 132608 265676 132660
rect 184204 132540 184256 132592
rect 213920 132540 213972 132592
rect 171784 132472 171836 132524
rect 214012 132472 214064 132524
rect 236644 132472 236696 132524
rect 265900 132472 265952 132524
rect 231768 132404 231820 132456
rect 247684 132404 247736 132456
rect 282828 132404 282880 132456
rect 307760 132404 307812 132456
rect 231676 132336 231728 132388
rect 246396 132336 246448 132388
rect 250444 131248 250496 131300
rect 265164 131248 265216 131300
rect 206284 131180 206336 131232
rect 213920 131180 213972 131232
rect 247868 131180 247920 131232
rect 265624 131180 265676 131232
rect 186964 131112 187016 131164
rect 214012 131112 214064 131164
rect 231492 131112 231544 131164
rect 235540 131112 235592 131164
rect 246304 131112 246356 131164
rect 265900 131112 265952 131164
rect 231768 131044 231820 131096
rect 264244 131044 264296 131096
rect 282828 131044 282880 131096
rect 302332 131044 302384 131096
rect 231400 130976 231452 131028
rect 260288 130976 260340 131028
rect 231676 130908 231728 130960
rect 246488 130908 246540 130960
rect 282276 130568 282328 130620
rect 285864 130568 285916 130620
rect 176016 129820 176068 129872
rect 214012 129820 214064 129872
rect 174636 129752 174688 129804
rect 213920 129752 213972 129804
rect 231308 129684 231360 129736
rect 240784 129684 240836 129736
rect 231584 129004 231636 129056
rect 257436 129004 257488 129056
rect 282828 128460 282880 128512
rect 287152 128460 287204 128512
rect 257528 128392 257580 128444
rect 265624 128392 265676 128444
rect 177488 128324 177540 128376
rect 213920 128324 213972 128376
rect 244924 128324 244976 128376
rect 265900 128324 265952 128376
rect 231676 128256 231728 128308
rect 262956 128256 263008 128308
rect 281724 128256 281776 128308
rect 303804 128256 303856 128308
rect 231768 128188 231820 128240
rect 240876 128188 240928 128240
rect 231676 127780 231728 127832
rect 236920 127780 236972 127832
rect 252008 127032 252060 127084
rect 265900 127032 265952 127084
rect 174728 126964 174780 127016
rect 213920 126964 213972 127016
rect 240784 126964 240836 127016
rect 265348 126964 265400 127016
rect 231124 126896 231176 126948
rect 254768 126896 254820 126948
rect 305644 126896 305696 126948
rect 580172 126896 580224 126948
rect 231768 126828 231820 126880
rect 239680 126828 239732 126880
rect 231492 126216 231544 126268
rect 242348 126216 242400 126268
rect 242532 126216 242584 126268
rect 265992 126216 266044 126268
rect 188436 125672 188488 125724
rect 214012 125672 214064 125724
rect 257620 125672 257672 125724
rect 265256 125672 265308 125724
rect 63408 125604 63460 125656
rect 65156 125604 65208 125656
rect 167644 125604 167696 125656
rect 213920 125604 213972 125656
rect 247684 125604 247736 125656
rect 265900 125604 265952 125656
rect 231768 125536 231820 125588
rect 242256 125536 242308 125588
rect 282092 125536 282144 125588
rect 285680 125536 285732 125588
rect 231308 124924 231360 124976
rect 233884 124924 233936 124976
rect 230848 124856 230900 124908
rect 249524 124856 249576 124908
rect 282828 124652 282880 124704
rect 288532 124652 288584 124704
rect 251916 124312 251968 124364
rect 265992 124312 266044 124364
rect 199384 124244 199436 124296
rect 213920 124244 213972 124296
rect 249156 124244 249208 124296
rect 265532 124244 265584 124296
rect 167736 124176 167788 124228
rect 214012 124176 214064 124228
rect 240876 124176 240928 124228
rect 265900 124176 265952 124228
rect 231768 124108 231820 124160
rect 250628 124108 250680 124160
rect 282736 124108 282788 124160
rect 300860 124108 300912 124160
rect 282828 124040 282880 124092
rect 295340 124040 295392 124092
rect 231584 123564 231636 123616
rect 235264 123564 235316 123616
rect 230756 123496 230808 123548
rect 253204 123496 253256 123548
rect 242256 123428 242308 123480
rect 265716 123428 265768 123480
rect 250536 122952 250588 123004
rect 265072 122952 265124 123004
rect 170588 122884 170640 122936
rect 213920 122884 213972 122936
rect 254676 122884 254728 122936
rect 265532 122884 265584 122936
rect 166356 122816 166408 122868
rect 214012 122816 214064 122868
rect 231308 122748 231360 122800
rect 260196 122748 260248 122800
rect 282092 122748 282144 122800
rect 309140 122748 309192 122800
rect 167920 122068 167972 122120
rect 198096 122068 198148 122120
rect 231676 122068 231728 122120
rect 250720 122068 250772 122120
rect 211804 121524 211856 121576
rect 214472 121524 214524 121576
rect 253204 121524 253256 121576
rect 265992 121524 266044 121576
rect 198004 121456 198056 121508
rect 213920 121456 213972 121508
rect 233884 121456 233936 121508
rect 265900 121456 265952 121508
rect 231768 121388 231820 121440
rect 258908 121388 258960 121440
rect 282460 121388 282512 121440
rect 302240 121388 302292 121440
rect 230940 121320 230992 121372
rect 238300 121320 238352 121372
rect 281724 121320 281776 121372
rect 291292 121320 291344 121372
rect 231216 120708 231268 120760
rect 264520 120708 264572 120760
rect 178776 120164 178828 120216
rect 213920 120164 213972 120216
rect 258816 120164 258868 120216
rect 265992 120164 266044 120216
rect 170680 120096 170732 120148
rect 214012 120096 214064 120148
rect 238024 120096 238076 120148
rect 265900 120096 265952 120148
rect 230940 120028 230992 120080
rect 255964 120028 256016 120080
rect 282092 120028 282144 120080
rect 298192 120028 298244 120080
rect 231492 119960 231544 120012
rect 249432 119960 249484 120012
rect 231768 119892 231820 119944
rect 239496 119892 239548 119944
rect 169116 118804 169168 118856
rect 214012 118804 214064 118856
rect 173440 118736 173492 118788
rect 213920 118736 213972 118788
rect 256148 118736 256200 118788
rect 265256 118736 265308 118788
rect 254768 118668 254820 118720
rect 265716 118668 265768 118720
rect 230664 118600 230716 118652
rect 263048 118600 263100 118652
rect 282828 118600 282880 118652
rect 292672 118600 292724 118652
rect 231768 118532 231820 118584
rect 242164 118532 242216 118584
rect 282736 118532 282788 118584
rect 289912 118532 289964 118584
rect 230940 117512 230992 117564
rect 236736 117512 236788 117564
rect 262956 117444 263008 117496
rect 265164 117444 265216 117496
rect 191196 117376 191248 117428
rect 214012 117376 214064 117428
rect 257436 117376 257488 117428
rect 265532 117376 265584 117428
rect 169208 117308 169260 117360
rect 213920 117308 213972 117360
rect 239496 117308 239548 117360
rect 265716 117308 265768 117360
rect 230664 117240 230716 117292
rect 252192 117240 252244 117292
rect 282828 117240 282880 117292
rect 306472 117240 306524 117292
rect 282736 117172 282788 117224
rect 295432 117172 295484 117224
rect 231216 116560 231268 116612
rect 250812 116560 250864 116612
rect 230572 116492 230624 116544
rect 232504 116492 232556 116544
rect 256240 116084 256292 116136
rect 264520 116084 264572 116136
rect 251824 116016 251876 116068
rect 266084 116016 266136 116068
rect 180156 115948 180208 116000
rect 213920 115948 213972 116000
rect 246396 115948 246448 116000
rect 266176 115948 266228 116000
rect 231768 115880 231820 115932
rect 246672 115880 246724 115932
rect 281724 115880 281776 115932
rect 303620 115880 303672 115932
rect 282092 115812 282144 115864
rect 296904 115812 296956 115864
rect 231584 115200 231636 115252
rect 264428 115200 264480 115252
rect 231768 115132 231820 115184
rect 238208 115132 238260 115184
rect 209136 114588 209188 114640
rect 214012 114588 214064 114640
rect 172060 114520 172112 114572
rect 213920 114520 213972 114572
rect 246488 114520 246540 114572
rect 265256 114520 265308 114572
rect 230572 114452 230624 114504
rect 232780 114452 232832 114504
rect 230664 114384 230716 114436
rect 239588 114384 239640 114436
rect 231492 114316 231544 114368
rect 245200 114316 245252 114368
rect 282828 113908 282880 113960
rect 288440 113908 288492 113960
rect 256056 113296 256108 113348
rect 265716 113296 265768 113348
rect 187056 113228 187108 113280
rect 213920 113228 213972 113280
rect 245108 113228 245160 113280
rect 265256 113228 265308 113280
rect 167828 113160 167880 113212
rect 214012 113160 214064 113212
rect 235264 113160 235316 113212
rect 265440 113160 265492 113212
rect 230940 113092 230992 113144
rect 241152 113092 241204 113144
rect 282092 113092 282144 113144
rect 294052 113092 294104 113144
rect 231676 112684 231728 112736
rect 234160 112684 234212 112736
rect 231492 112412 231544 112464
rect 258724 112412 258776 112464
rect 260288 111936 260340 111988
rect 265716 111936 265768 111988
rect 211896 111868 211948 111920
rect 214012 111868 214064 111920
rect 242164 111868 242216 111920
rect 265532 111868 265584 111920
rect 166448 111800 166500 111852
rect 213920 111800 213972 111852
rect 240968 111800 241020 111852
rect 266084 111800 266136 111852
rect 231768 111732 231820 111784
rect 261852 111732 261904 111784
rect 282828 111732 282880 111784
rect 299572 111732 299624 111784
rect 231676 111664 231728 111716
rect 241060 111664 241112 111716
rect 231676 111052 231728 111104
rect 245016 111052 245068 111104
rect 3424 110848 3476 110900
rect 7564 110848 7616 110900
rect 258908 110576 258960 110628
rect 265532 110576 265584 110628
rect 196716 110508 196768 110560
rect 213920 110508 213972 110560
rect 261576 110508 261628 110560
rect 265164 110508 265216 110560
rect 173256 110440 173308 110492
rect 214012 110440 214064 110492
rect 245200 110440 245252 110492
rect 265716 110440 265768 110492
rect 167460 110372 167512 110424
rect 170496 110372 170548 110424
rect 231768 110372 231820 110424
rect 261760 110372 261812 110424
rect 231124 110304 231176 110356
rect 254860 110304 254912 110356
rect 176108 109080 176160 109132
rect 213920 109080 213972 109132
rect 231584 109080 231636 109132
rect 235448 109080 235500 109132
rect 261852 109080 261904 109132
rect 265532 109080 265584 109132
rect 173164 109012 173216 109064
rect 214012 109012 214064 109064
rect 250628 109012 250680 109064
rect 265716 109012 265768 109064
rect 167920 108944 167972 108996
rect 173348 108944 173400 108996
rect 231124 108944 231176 108996
rect 263140 108944 263192 108996
rect 282828 108944 282880 108996
rect 306380 108944 306432 108996
rect 231768 108876 231820 108928
rect 246580 108876 246632 108928
rect 230848 108128 230900 108180
rect 232688 108128 232740 108180
rect 281540 107992 281592 108044
rect 284392 107992 284444 108044
rect 241060 107856 241112 107908
rect 265348 107856 265400 107908
rect 209044 107720 209096 107772
rect 214012 107720 214064 107772
rect 260196 107720 260248 107772
rect 265440 107720 265492 107772
rect 202236 107652 202288 107704
rect 213920 107652 213972 107704
rect 263048 107652 263100 107704
rect 265716 107652 265768 107704
rect 231768 107584 231820 107636
rect 249340 107584 249392 107636
rect 282460 107584 282512 107636
rect 298284 107584 298336 107636
rect 230572 107516 230624 107568
rect 232596 107516 232648 107568
rect 231400 106904 231452 106956
rect 264612 106904 264664 106956
rect 265440 106768 265492 106820
rect 265808 106768 265860 106820
rect 259092 106428 259144 106480
rect 265808 106428 265860 106480
rect 210516 106360 210568 106412
rect 214012 106360 214064 106412
rect 263140 106360 263192 106412
rect 265532 106360 265584 106412
rect 170496 106292 170548 106344
rect 213920 106292 213972 106344
rect 249064 106292 249116 106344
rect 265716 106292 265768 106344
rect 231768 106224 231820 106276
rect 259000 106224 259052 106276
rect 282828 106224 282880 106276
rect 305092 106224 305144 106276
rect 231676 106156 231728 106208
rect 238392 106156 238444 106208
rect 230480 105544 230532 105596
rect 256332 105544 256384 105596
rect 169300 105000 169352 105052
rect 214012 105000 214064 105052
rect 258724 105000 258776 105052
rect 266084 105000 266136 105052
rect 204996 104932 205048 104984
rect 213920 104932 213972 104984
rect 255964 104932 256016 104984
rect 265716 104932 265768 104984
rect 246580 104864 246632 104916
rect 265808 104864 265860 104916
rect 231768 104796 231820 104848
rect 245292 104796 245344 104848
rect 231584 104660 231636 104712
rect 234068 104660 234120 104712
rect 235908 104116 235960 104168
rect 265440 104116 265492 104168
rect 230664 103776 230716 103828
rect 235356 103776 235408 103828
rect 205088 103504 205140 103556
rect 213920 103504 213972 103556
rect 245016 103504 245068 103556
rect 265808 103504 265860 103556
rect 231768 103436 231820 103488
rect 252100 103436 252152 103488
rect 282828 103436 282880 103488
rect 299664 103436 299716 103488
rect 231584 103300 231636 103352
rect 233976 103300 234028 103352
rect 249340 102212 249392 102264
rect 265808 102212 265860 102264
rect 232504 102144 232556 102196
rect 265716 102144 265768 102196
rect 230572 102076 230624 102128
rect 242256 102076 242308 102128
rect 231124 102008 231176 102060
rect 235908 102008 235960 102060
rect 167920 101396 167972 101448
rect 214564 101396 214616 101448
rect 254860 100852 254912 100904
rect 265532 100852 265584 100904
rect 207756 100784 207808 100836
rect 214012 100784 214064 100836
rect 242440 100784 242492 100836
rect 265716 100784 265768 100836
rect 184296 100716 184348 100768
rect 213920 100716 213972 100768
rect 238208 100716 238260 100768
rect 265808 100716 265860 100768
rect 231676 100648 231728 100700
rect 260380 100648 260432 100700
rect 385684 100648 385736 100700
rect 580172 100648 580224 100700
rect 231768 100580 231820 100632
rect 243728 100580 243780 100632
rect 260472 99492 260524 99544
rect 265808 99492 265860 99544
rect 252100 99424 252152 99476
rect 265716 99424 265768 99476
rect 164884 99356 164936 99408
rect 213920 99356 213972 99408
rect 243636 99356 243688 99408
rect 265532 99356 265584 99408
rect 265808 99356 265860 99408
rect 266084 99356 266136 99408
rect 231492 99288 231544 99340
rect 242532 99288 242584 99340
rect 282828 99288 282880 99340
rect 299480 99288 299532 99340
rect 209228 98064 209280 98116
rect 213920 98064 213972 98116
rect 242348 98064 242400 98116
rect 265808 98064 265860 98116
rect 166540 97996 166592 98048
rect 214012 97996 214064 98048
rect 235356 97996 235408 98048
rect 265440 97996 265492 98048
rect 3424 97928 3476 97980
rect 21364 97928 21416 97980
rect 242256 96704 242308 96756
rect 265164 96704 265216 96756
rect 207664 96636 207716 96688
rect 213920 96636 213972 96688
rect 234068 96636 234120 96688
rect 265808 96636 265860 96688
rect 193128 96568 193180 96620
rect 229008 96568 229060 96620
rect 267004 96364 267056 96416
rect 281540 96364 281592 96416
rect 229008 95888 229060 95940
rect 230480 95888 230532 95940
rect 268016 95888 268068 95940
rect 228364 95208 228416 95260
rect 265808 95208 265860 95260
rect 187608 95140 187660 95192
rect 280160 95140 280212 95192
rect 215944 95072 215996 95124
rect 281632 95072 281684 95124
rect 63408 95004 63460 95056
rect 205088 95004 205140 95056
rect 267280 95004 267332 95056
rect 279516 95004 279568 95056
rect 267096 94936 267148 94988
rect 280344 94936 280396 94988
rect 122840 94460 122892 94512
rect 214656 94460 214708 94512
rect 128084 93984 128136 94036
rect 171876 93984 171928 94036
rect 112352 93916 112404 93968
rect 173440 93916 173492 93968
rect 105728 93848 105780 93900
rect 186964 93848 187016 93900
rect 231124 93780 231176 93832
rect 253848 93780 253900 93832
rect 268016 93780 268068 93832
rect 276940 93780 276992 93832
rect 270960 93712 271012 93764
rect 151728 93440 151780 93492
rect 169024 93440 169076 93492
rect 134432 93372 134484 93424
rect 174544 93372 174596 93424
rect 121736 93304 121788 93356
rect 166356 93304 166408 93356
rect 88984 93236 89036 93288
rect 164884 93236 164936 93288
rect 111248 93168 111300 93220
rect 191196 93168 191248 93220
rect 230480 93168 230532 93220
rect 233976 93168 234028 93220
rect 106464 93100 106516 93152
rect 209136 93100 209188 93152
rect 216312 92556 216364 92608
rect 220084 92556 220136 92608
rect 180616 92420 180668 92472
rect 281816 92420 281868 92472
rect 98552 92352 98604 92404
rect 196716 92352 196768 92404
rect 118056 92284 118108 92336
rect 202144 92284 202196 92336
rect 110696 92216 110748 92268
rect 122840 92216 122892 92268
rect 126704 92216 126756 92268
rect 188344 92216 188396 92268
rect 133144 92148 133196 92200
rect 167920 92148 167972 92200
rect 151544 92080 151596 92132
rect 180064 92080 180116 92132
rect 106648 92012 106700 92064
rect 184204 92012 184256 92064
rect 104624 91128 104676 91180
rect 117964 91128 118016 91180
rect 86592 91060 86644 91112
rect 110420 91060 110472 91112
rect 104348 90992 104400 91044
rect 167828 90992 167880 91044
rect 126520 90924 126572 90976
rect 188436 90924 188488 90976
rect 110144 90856 110196 90908
rect 169208 90856 169260 90908
rect 151360 90788 151412 90840
rect 177396 90788 177448 90840
rect 188344 90312 188396 90364
rect 265992 90312 266044 90364
rect 67456 89632 67508 89684
rect 207756 89632 207808 89684
rect 90364 89564 90416 89616
rect 169300 89564 169352 89616
rect 119896 89496 119948 89548
rect 198004 89496 198056 89548
rect 106004 89428 106056 89480
rect 172060 89428 172112 89480
rect 132408 89360 132460 89412
rect 178684 89360 178736 89412
rect 215944 88952 215996 89004
rect 265900 88952 265952 89004
rect 84660 88272 84712 88324
rect 184296 88272 184348 88324
rect 100576 88204 100628 88256
rect 166448 88204 166500 88256
rect 117136 88136 117188 88188
rect 170680 88136 170732 88188
rect 115572 88068 115624 88120
rect 169116 88068 169168 88120
rect 123760 88000 123812 88052
rect 175924 88000 175976 88052
rect 124036 87932 124088 87984
rect 167736 87932 167788 87984
rect 101864 86912 101916 86964
rect 211896 86912 211948 86964
rect 110420 86844 110472 86896
rect 209228 86844 209280 86896
rect 97080 86776 97132 86828
rect 174728 86776 174780 86828
rect 109500 86708 109552 86760
rect 180156 86708 180208 86760
rect 120816 86640 120868 86692
rect 170588 86640 170640 86692
rect 3424 85484 3476 85536
rect 25504 85484 25556 85536
rect 64788 85484 64840 85536
rect 207664 85484 207716 85536
rect 114376 85416 114428 85468
rect 213184 85416 213236 85468
rect 103060 85348 103112 85400
rect 187056 85348 187108 85400
rect 92296 85280 92348 85332
rect 170496 85280 170548 85332
rect 152648 85212 152700 85264
rect 196624 85212 196676 85264
rect 125416 85144 125468 85196
rect 167644 85144 167696 85196
rect 108856 84124 108908 84176
rect 213368 84124 213420 84176
rect 121368 84056 121420 84108
rect 210424 84056 210476 84108
rect 86868 83988 86920 84040
rect 166540 83988 166592 84040
rect 96528 83920 96580 83972
rect 176108 83920 176160 83972
rect 115848 83852 115900 83904
rect 178776 83852 178828 83904
rect 136548 83784 136600 83836
rect 166264 83784 166316 83836
rect 75828 82764 75880 82816
rect 214564 82764 214616 82816
rect 114468 82696 114520 82748
rect 213276 82696 213328 82748
rect 103428 82628 103480 82680
rect 176016 82628 176068 82680
rect 125508 82560 125560 82612
rect 170404 82560 170456 82612
rect 95056 81336 95108 81388
rect 202236 81336 202288 81388
rect 118608 81268 118660 81320
rect 211804 81268 211856 81320
rect 129648 81200 129700 81252
rect 177304 81200 177356 81252
rect 93768 79976 93820 80028
rect 210516 79976 210568 80028
rect 117228 79908 117280 79960
rect 206376 79908 206428 79960
rect 124128 79840 124180 79892
rect 199384 79840 199436 79892
rect 100668 79772 100720 79824
rect 173256 79772 173308 79824
rect 108948 79704 109000 79756
rect 171784 79704 171836 79756
rect 95148 78616 95200 78668
rect 209044 78616 209096 78668
rect 110328 78548 110380 78600
rect 204904 78548 204956 78600
rect 99288 78480 99340 78532
rect 177488 78480 177540 78532
rect 102048 78412 102100 78464
rect 174636 78412 174688 78464
rect 67548 77188 67600 77240
rect 214748 77188 214800 77240
rect 97908 77120 97960 77172
rect 173164 77120 173216 77172
rect 13820 76508 13872 76560
rect 252008 76508 252060 76560
rect 125600 75284 125652 75336
rect 191104 75284 191156 75336
rect 95240 75216 95292 75268
rect 253388 75216 253440 75268
rect 75920 75148 75972 75200
rect 259092 75148 259144 75200
rect 117964 74468 118016 74520
rect 206284 74468 206336 74520
rect 99380 73856 99432 73908
rect 249248 73856 249300 73908
rect 78680 73788 78732 73840
rect 263140 73788 263192 73840
rect 96620 72428 96672 72480
rect 250628 72428 250680 72480
rect 74540 69708 74592 69760
rect 229836 69708 229888 69760
rect 100760 69640 100812 69692
rect 261852 69640 261904 69692
rect 107660 68348 107712 68400
rect 245200 68348 245252 68400
rect 52460 68280 52512 68332
rect 247868 68280 247920 68332
rect 103520 66920 103572 66972
rect 264520 66920 264572 66972
rect 41420 66852 41472 66904
rect 256240 66852 256292 66904
rect 110420 65560 110472 65612
rect 247776 65560 247828 65612
rect 16580 65492 16632 65544
rect 260472 65492 260524 65544
rect 121460 64200 121512 64252
rect 260288 64200 260340 64252
rect 30380 64132 30432 64184
rect 246488 64132 246540 64184
rect 20720 62772 20772 62824
rect 252100 62772 252152 62824
rect 64880 61412 64932 61464
rect 246580 61412 246632 61464
rect 29000 61344 29052 61396
rect 242440 61344 242492 61396
rect 82820 60052 82872 60104
rect 241060 60052 241112 60104
rect 33140 59984 33192 60036
rect 254860 59984 254912 60036
rect 3056 59304 3108 59356
rect 43444 59304 43496 59356
rect 122840 58692 122892 58744
rect 257620 58692 257672 58744
rect 43536 58624 43588 58676
rect 231124 58624 231176 58676
rect 93860 57196 93912 57248
rect 263048 57196 263100 57248
rect 118700 55836 118752 55888
rect 240968 55836 241020 55888
rect 98000 54544 98052 54596
rect 250536 54544 250588 54596
rect 55220 54476 55272 54528
rect 262956 54476 263008 54528
rect 109040 53116 109092 53168
rect 251916 53116 251968 53168
rect 24860 53048 24912 53100
rect 242348 53048 242400 53100
rect 35900 51688 35952 51740
rect 249340 51688 249392 51740
rect 66260 50396 66312 50448
rect 256148 50396 256200 50448
rect 19340 50328 19392 50380
rect 235356 50328 235408 50380
rect 69020 49036 69072 49088
rect 254768 49036 254820 49088
rect 15200 48968 15252 49020
rect 234068 48968 234120 49020
rect 11060 47540 11112 47592
rect 242256 47540 242308 47592
rect 322204 46860 322256 46912
rect 580172 46860 580224 46912
rect 115940 46180 115992 46232
rect 240876 46180 240928 46232
rect 2872 45500 2924 45552
rect 4804 45500 4856 45552
rect 111800 44820 111852 44872
rect 249156 44820 249208 44872
rect 56600 43392 56652 43444
rect 250444 43392 250496 43444
rect 104900 42100 104952 42152
rect 264336 42100 264388 42152
rect 35992 42032 36044 42084
rect 257528 42032 257580 42084
rect 63500 40672 63552 40724
rect 236644 40672 236696 40724
rect 67640 39380 67692 39432
rect 262864 39380 262916 39432
rect 17960 39312 18012 39364
rect 245108 39312 245160 39364
rect 102140 37952 102192 38004
rect 254676 37952 254728 38004
rect 60740 37884 60792 37936
rect 246304 37884 246356 37936
rect 81440 36524 81492 36576
rect 253296 36524 253348 36576
rect 86960 35232 87012 35284
rect 261668 35232 261720 35284
rect 12440 35164 12492 35216
rect 235264 35164 235316 35216
rect 106924 33736 106976 33788
rect 265624 33736 265676 33788
rect 3516 33056 3568 33108
rect 18604 33056 18656 33108
rect 302884 33056 302936 33108
rect 580172 33056 580224 33108
rect 85580 32444 85632 32496
rect 238116 32444 238168 32496
rect 53840 32376 53892 32428
rect 265716 32376 265768 32428
rect 52552 31084 52604 31136
rect 239496 31084 239548 31136
rect 59360 31016 59412 31068
rect 257436 31016 257488 31068
rect 80060 29656 80112 29708
rect 258816 29656 258868 29708
rect 48320 29588 48372 29640
rect 246396 29588 246448 29640
rect 88340 28296 88392 28348
rect 261484 28296 261536 28348
rect 8300 28228 8352 28280
rect 242164 28228 242216 28280
rect 57980 26936 58032 26988
rect 264428 26936 264480 26988
rect 22100 26868 22152 26920
rect 256056 26868 256108 26920
rect 114560 25576 114612 25628
rect 258908 25576 258960 25628
rect 26240 25508 26292 25560
rect 238208 25508 238260 25560
rect 110512 24148 110564 24200
rect 261576 24148 261628 24200
rect 9680 24080 9732 24132
rect 247684 24080 247736 24132
rect 92480 22720 92532 22772
rect 260104 22720 260156 22772
rect 91100 21428 91152 21480
rect 253204 21428 253256 21480
rect 23480 21360 23532 21412
rect 240784 21360 240836 21412
rect 3424 20612 3476 20664
rect 39304 20612 39356 20664
rect 44272 20000 44324 20052
rect 251824 20000 251876 20052
rect 4160 19932 4212 19984
rect 228364 19932 228416 19984
rect 85672 18640 85724 18692
rect 264244 18640 264296 18692
rect 38660 18572 38712 18624
rect 244924 18572 244976 18624
rect 84200 17212 84252 17264
rect 233884 17212 233936 17264
rect 120632 15920 120684 15972
rect 257344 15920 257396 15972
rect 11888 15852 11940 15904
rect 243636 15852 243688 15904
rect 117320 14492 117372 14544
rect 229744 14492 229796 14544
rect 69112 14424 69164 14476
rect 255964 14424 256016 14476
rect 114008 13132 114060 13184
rect 243544 13132 243596 13184
rect 61568 13064 61620 13116
rect 258724 13064 258776 13116
rect 106464 11704 106516 11756
rect 239404 11704 239456 11756
rect 78588 8984 78640 9036
rect 254584 8984 254636 9036
rect 51356 8916 51408 8968
rect 245016 8916 245068 8968
rect 90364 7556 90416 7608
rect 260196 7556 260248 7608
rect 3424 6808 3476 6860
rect 35164 6808 35216 6860
rect 220084 6808 220136 6860
rect 580172 6808 580224 6860
rect 72608 6196 72660 6248
rect 249064 6196 249116 6248
rect 47860 6128 47912 6180
rect 232504 6128 232556 6180
rect 73804 4768 73856 4820
rect 238024 4768 238076 4820
rect 2780 3476 2832 3528
rect 3700 3476 3752 3528
rect 19340 3476 19392 3528
rect 20260 3476 20312 3528
rect 35900 3476 35952 3528
rect 36820 3476 36872 3528
rect 52460 3476 52512 3528
rect 53380 3476 53432 3528
rect 69020 3476 69072 3528
rect 69940 3476 69992 3528
rect 95148 3476 95200 3528
rect 188344 3476 188396 3528
rect 233976 3476 234028 3528
rect 235816 3476 235868 3528
rect 572 3408 624 3460
rect 43536 3408 43588 3460
rect 50160 3408 50212 3460
rect 106924 3408 106976 3460
rect 119896 3408 119948 3460
rect 215944 3408 215996 3460
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2778 423600 2834 423609
rect 2778 423535 2780 423544
rect 2832 423535 2834 423544
rect 2780 423506 2832 423512
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3436 300150 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 6932 632738 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700330 24348 703520
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 6920 632732 6972 632738
rect 6920 632674 6972 632680
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 7564 632120 7616 632126
rect 3568 632088 3570 632097
rect 7564 632062 7616 632068
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 4804 423564 4856 423570
rect 4804 423506 4856 423512
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3528 371278 3556 371311
rect 3516 371272 3568 371278
rect 3516 371214 3568 371220
rect 3424 300144 3476 300150
rect 3424 300086 3476 300092
rect 4816 298790 4844 423506
rect 4804 298784 4856 298790
rect 4804 298726 4856 298732
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3422 290864 3478 290873
rect 3422 290799 3478 290808
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3160 253978 3188 254079
rect 3148 253972 3200 253978
rect 3148 253914 3200 253920
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240174 3096 241023
rect 3056 240168 3108 240174
rect 3056 240110 3108 240116
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3436 162897 3464 290799
rect 3516 284980 3568 284986
rect 3516 284922 3568 284928
rect 3528 188873 3556 284922
rect 3606 267200 3662 267209
rect 3606 267135 3662 267144
rect 3620 244934 3648 267135
rect 7576 266354 7604 632062
rect 14464 553444 14516 553450
rect 14464 553386 14516 553392
rect 11704 448588 11756 448594
rect 11704 448530 11756 448536
rect 11716 296002 11744 448530
rect 11704 295996 11756 296002
rect 11704 295938 11756 295944
rect 11704 291236 11756 291242
rect 11704 291178 11756 291184
rect 7564 266348 7616 266354
rect 7564 266290 7616 266296
rect 3608 244928 3660 244934
rect 3608 244870 3660 244876
rect 7564 220108 7616 220114
rect 7564 220050 7616 220056
rect 4804 218748 4856 218754
rect 4804 218690 4856 218696
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 3516 185632 3568 185638
rect 3516 185574 3568 185580
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3424 137964 3476 137970
rect 3424 137906 3476 137912
rect 3436 136785 3464 137906
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3424 110900 3476 110906
rect 3424 110842 3476 110848
rect 3436 110673 3464 110842
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3424 85536 3476 85542
rect 3424 85478 3476 85484
rect 3436 84697 3464 85478
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3528 71641 3556 185574
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 2778 55856 2834 55865
rect 2778 55791 2834 55800
rect 1398 44840 1454 44849
rect 1398 44775 1454 44784
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 542 -960 654 480
rect 1412 354 1440 44775
rect 2792 3534 2820 55791
rect 4816 45558 4844 218690
rect 7576 110906 7604 220050
rect 11716 150414 11744 291178
rect 14476 263566 14504 553386
rect 15844 409896 15896 409902
rect 15844 409838 15896 409844
rect 14464 263560 14516 263566
rect 14464 263502 14516 263508
rect 14464 256760 14516 256766
rect 14464 256702 14516 256708
rect 11704 150408 11756 150414
rect 11704 150350 11756 150356
rect 14476 137970 14504 256702
rect 15856 247042 15884 409838
rect 39302 292904 39358 292913
rect 39302 292839 39358 292848
rect 21364 292596 21416 292602
rect 21364 292538 21416 292544
rect 18604 267776 18656 267782
rect 18604 267718 18656 267724
rect 17224 263628 17276 263634
rect 17224 263570 17276 263576
rect 15844 247036 15896 247042
rect 15844 246978 15896 246984
rect 17236 215286 17264 263570
rect 17224 215280 17276 215286
rect 17224 215222 17276 215228
rect 14464 137964 14516 137970
rect 14464 137906 14516 137912
rect 7564 110900 7616 110906
rect 7564 110842 7616 110848
rect 13820 76560 13872 76566
rect 13820 76502 13872 76508
rect 11060 47592 11112 47598
rect 11060 47534 11112 47540
rect 2872 45552 2924 45558
rect 2870 45520 2872 45529
rect 4804 45552 4856 45558
rect 2924 45520 2926 45529
rect 4804 45494 4856 45500
rect 2870 45455 2926 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 8300 28280 8352 28286
rect 8300 28222 8352 28228
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 19926
rect 8312 16574 8340 28222
rect 9680 24132 9732 24138
rect 9680 24074 9732 24080
rect 4172 16546 5304 16574
rect 8312 16546 8800 16574
rect 2870 10296 2926 10305
rect 2870 10231 2926 10240
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 480 2912 10231
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 3712 354 3740 3470
rect 5276 480 5304 16546
rect 7654 11656 7710 11665
rect 7654 11591 7710 11600
rect 6458 4856 6514 4865
rect 6458 4791 6514 4800
rect 6472 480 6500 4791
rect 7668 480 7696 11591
rect 8772 480 8800 16546
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 24074
rect 11072 16574 11100 47534
rect 12440 35216 12492 35222
rect 12440 35158 12492 35164
rect 12452 16574 12480 35158
rect 13832 16574 13860 76502
rect 16580 65544 16632 65550
rect 16580 65486 16632 65492
rect 15200 49020 15252 49026
rect 15200 48962 15252 48968
rect 15212 16574 15240 48962
rect 16592 16574 16620 65486
rect 17960 39364 18012 39370
rect 17960 39306 18012 39312
rect 11072 16546 11192 16574
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 11164 480 11192 16546
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 15846
rect 13556 480 13584 16546
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 39306
rect 18616 33114 18644 267718
rect 21376 244254 21404 292538
rect 35164 278792 35216 278798
rect 35164 278734 35216 278740
rect 25504 252612 25556 252618
rect 25504 252554 25556 252560
rect 21364 244248 21416 244254
rect 21364 244190 21416 244196
rect 21364 228404 21416 228410
rect 21364 228346 21416 228352
rect 21376 97986 21404 228346
rect 21364 97980 21416 97986
rect 21364 97922 21416 97928
rect 25516 85542 25544 252554
rect 25504 85536 25556 85542
rect 25504 85478 25556 85484
rect 27618 71088 27674 71097
rect 27618 71023 27674 71032
rect 20720 62824 20772 62830
rect 20720 62766 20772 62772
rect 19340 50380 19392 50386
rect 19340 50322 19392 50328
rect 18604 33108 18656 33114
rect 18604 33050 18656 33056
rect 19352 3534 19380 50322
rect 19430 36544 19486 36553
rect 19430 36479 19486 36488
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19444 480 19472 36479
rect 20732 16574 20760 62766
rect 24860 53100 24912 53106
rect 24860 53042 24912 53048
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22112 16574 22140 26862
rect 23480 21412 23532 21418
rect 23480 21354 23532 21360
rect 23492 16574 23520 21354
rect 24872 16574 24900 53042
rect 26240 25560 26292 25566
rect 26240 25502 26292 25508
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20272 354 20300 3470
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20272 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 25502
rect 27632 6914 27660 71023
rect 30380 64184 30432 64190
rect 30380 64126 30432 64132
rect 29000 61396 29052 61402
rect 29000 61338 29052 61344
rect 27710 40624 27766 40633
rect 27710 40559 27766 40568
rect 27724 16574 27752 40559
rect 29012 16574 29040 61338
rect 30392 16574 30420 64126
rect 33140 60036 33192 60042
rect 33140 59978 33192 59984
rect 31758 43480 31814 43489
rect 31758 43415 31814 43424
rect 31772 16574 31800 43415
rect 33152 16574 33180 59978
rect 27724 16546 28488 16574
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 27632 6886 27752 6914
rect 27724 480 27752 6886
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 34794 7576 34850 7585
rect 34794 7511 34850 7520
rect 34808 480 34836 7511
rect 35176 6866 35204 278734
rect 35900 51740 35952 51746
rect 35900 51682 35952 51688
rect 35164 6860 35216 6866
rect 35164 6802 35216 6808
rect 35912 3534 35940 51682
rect 35992 42084 36044 42090
rect 35992 42026 36044 42032
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36004 480 36032 42026
rect 37278 33824 37334 33833
rect 37278 33759 37334 33768
rect 37292 16574 37320 33759
rect 39316 20670 39344 292839
rect 40052 238649 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 54484 700324 54536 700330
rect 54484 700266 54536 700272
rect 54496 320890 54524 700266
rect 71044 670744 71096 670750
rect 71044 670686 71096 670692
rect 54484 320884 54536 320890
rect 54484 320826 54536 320832
rect 43444 294364 43496 294370
rect 43444 294306 43496 294312
rect 40038 238640 40094 238649
rect 40038 238575 40094 238584
rect 41420 66904 41472 66910
rect 41420 66846 41472 66852
rect 40038 57216 40094 57225
rect 40038 57151 40094 57160
rect 39304 20664 39356 20670
rect 39304 20606 39356 20612
rect 38660 18624 38712 18630
rect 38660 18566 38712 18572
rect 38672 16574 38700 18566
rect 40052 16574 40080 57151
rect 41432 16574 41460 66846
rect 43456 59362 43484 294306
rect 71056 287026 71084 670686
rect 71792 316742 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 318102 88380 702406
rect 97264 605872 97316 605878
rect 97264 605814 97316 605820
rect 94504 527196 94556 527202
rect 94504 527138 94556 527144
rect 88340 318096 88392 318102
rect 88340 318038 88392 318044
rect 71780 316736 71832 316742
rect 71780 316678 71832 316684
rect 71044 287020 71096 287026
rect 71044 286962 71096 286968
rect 94516 260846 94544 527138
rect 97276 304366 97304 605814
rect 97264 304360 97316 304366
rect 97264 304302 97316 304308
rect 94504 260840 94556 260846
rect 94504 260782 94556 260788
rect 104912 242185 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 137848 700330 137876 703520
rect 137836 700324 137888 700330
rect 137836 700266 137888 700272
rect 154132 698970 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 698964 154172 698970
rect 154120 698906 154172 698912
rect 116584 618316 116636 618322
rect 116584 618258 116636 618264
rect 108304 565888 108356 565894
rect 108304 565830 108356 565836
rect 108316 267714 108344 565830
rect 116596 274650 116624 618258
rect 166264 462392 166316 462398
rect 166264 462334 166316 462340
rect 162124 318844 162176 318850
rect 162124 318786 162176 318792
rect 162136 302938 162164 318786
rect 162124 302932 162176 302938
rect 162124 302874 162176 302880
rect 116584 274644 116636 274650
rect 116584 274586 116636 274592
rect 108304 267708 108356 267714
rect 108304 267650 108356 267656
rect 104898 242176 104954 242185
rect 104898 242111 104954 242120
rect 166276 235890 166304 462334
rect 169772 271862 169800 702406
rect 177948 700392 178000 700398
rect 177948 700334 178000 700340
rect 173164 371272 173216 371278
rect 173164 371214 173216 371220
rect 169760 271856 169812 271862
rect 169760 271798 169812 271804
rect 172428 260908 172480 260914
rect 172428 260850 172480 260856
rect 169024 253972 169076 253978
rect 169024 253914 169076 253920
rect 169036 240038 169064 253914
rect 169024 240032 169076 240038
rect 169024 239974 169076 239980
rect 166264 235884 166316 235890
rect 166264 235826 166316 235832
rect 172440 189922 172468 260850
rect 173176 238474 173204 371214
rect 175188 259480 175240 259486
rect 175188 259422 175240 259428
rect 173164 238468 173216 238474
rect 173164 238410 173216 238416
rect 172428 189916 172480 189922
rect 172428 189858 172480 189864
rect 175200 189854 175228 259422
rect 177856 255332 177908 255338
rect 177856 255274 177908 255280
rect 175188 189848 175240 189854
rect 175188 189790 175240 189796
rect 177868 189786 177896 255274
rect 177960 238746 177988 700334
rect 178684 700324 178736 700330
rect 178684 700266 178736 700272
rect 184848 700324 184900 700330
rect 184848 700266 184900 700272
rect 178696 249762 178724 700266
rect 180708 697604 180760 697610
rect 180708 697546 180760 697552
rect 180524 295384 180576 295390
rect 180524 295326 180576 295332
rect 179326 273864 179382 273873
rect 179326 273799 179382 273808
rect 178684 249756 178736 249762
rect 178684 249698 178736 249704
rect 177948 238740 178000 238746
rect 177948 238682 178000 238688
rect 177856 189780 177908 189786
rect 177856 189722 177908 189728
rect 100668 183592 100720 183598
rect 100668 183534 100720 183540
rect 97540 179580 97592 179586
rect 97540 179522 97592 179528
rect 97552 177041 97580 179522
rect 99102 179480 99158 179489
rect 99102 179415 99158 179424
rect 99116 177041 99144 179415
rect 97538 177032 97594 177041
rect 97538 176967 97594 176976
rect 99102 177032 99158 177041
rect 99102 176967 99158 176976
rect 100680 176769 100708 183534
rect 127072 182436 127124 182442
rect 127072 182378 127124 182384
rect 170588 182436 170640 182442
rect 170588 182378 170640 182384
rect 108120 182368 108172 182374
rect 108120 182310 108172 182316
rect 105912 182300 105964 182306
rect 105912 182242 105964 182248
rect 103336 181008 103388 181014
rect 103336 180950 103388 180956
rect 103348 176769 103376 180950
rect 105924 177721 105952 182242
rect 108132 177721 108160 182310
rect 124956 181076 125008 181082
rect 124956 181018 125008 181024
rect 114468 180940 114520 180946
rect 114468 180882 114520 180888
rect 114376 179444 114428 179450
rect 114376 179386 114428 179392
rect 110696 178288 110748 178294
rect 110696 178230 110748 178236
rect 109592 178084 109644 178090
rect 109592 178026 109644 178032
rect 105910 177712 105966 177721
rect 105910 177647 105966 177656
rect 108118 177712 108174 177721
rect 108118 177647 108174 177656
rect 107016 176996 107068 177002
rect 107016 176938 107068 176944
rect 104624 176860 104676 176866
rect 104624 176802 104676 176808
rect 104636 176769 104664 176802
rect 107028 176769 107056 176938
rect 109604 176769 109632 178026
rect 110708 176769 110736 178230
rect 112260 178220 112312 178226
rect 112260 178162 112312 178168
rect 112272 176769 112300 178162
rect 114388 177177 114416 179386
rect 114480 177721 114508 180882
rect 119528 180872 119580 180878
rect 119528 180814 119580 180820
rect 118424 178356 118476 178362
rect 118424 178298 118476 178304
rect 114466 177712 114522 177721
rect 114466 177647 114522 177656
rect 114374 177168 114430 177177
rect 114374 177103 114430 177112
rect 118436 176769 118464 178298
rect 119540 177721 119568 180814
rect 123760 179648 123812 179654
rect 123760 179590 123812 179596
rect 119526 177712 119582 177721
rect 119526 177647 119582 177656
rect 123772 177177 123800 179590
rect 124968 177721 124996 181018
rect 127084 177721 127112 182378
rect 169024 182368 169076 182374
rect 169024 182310 169076 182316
rect 167644 182300 167696 182306
rect 167644 182242 167696 182248
rect 130752 182232 130804 182238
rect 130752 182174 130804 182180
rect 129464 179512 129516 179518
rect 129464 179454 129516 179460
rect 124954 177712 125010 177721
rect 124954 177647 125010 177656
rect 127070 177712 127126 177721
rect 127070 177647 127126 177656
rect 129476 177177 129504 179454
rect 130764 177721 130792 182174
rect 132408 181144 132460 181150
rect 132408 181086 132460 181092
rect 166540 181144 166592 181150
rect 166540 181086 166592 181092
rect 132420 177721 132448 181086
rect 166264 181008 166316 181014
rect 166264 180950 166316 180956
rect 133144 178152 133196 178158
rect 133144 178094 133196 178100
rect 130750 177712 130806 177721
rect 130750 177647 130806 177656
rect 132406 177712 132462 177721
rect 132406 177647 132462 177656
rect 123758 177168 123814 177177
rect 123758 177103 123814 177112
rect 129462 177168 129518 177177
rect 129462 177103 129518 177112
rect 128176 177064 128228 177070
rect 128176 177006 128228 177012
rect 125876 176792 125928 176798
rect 100666 176760 100722 176769
rect 100666 176695 100722 176704
rect 103334 176760 103390 176769
rect 103334 176695 103390 176704
rect 104622 176760 104678 176769
rect 104622 176695 104678 176704
rect 107014 176760 107070 176769
rect 107014 176695 107070 176704
rect 109590 176760 109646 176769
rect 109590 176695 109646 176704
rect 110694 176760 110750 176769
rect 110694 176695 110750 176704
rect 112258 176760 112314 176769
rect 112258 176695 112314 176704
rect 118422 176760 118478 176769
rect 118422 176695 118478 176704
rect 125874 176760 125876 176769
rect 128188 176769 128216 177006
rect 133156 176769 133184 178094
rect 165344 176996 165396 177002
rect 165344 176938 165396 176944
rect 148232 176928 148284 176934
rect 148232 176870 148284 176876
rect 148244 176769 148272 176870
rect 125928 176760 125930 176769
rect 125874 176695 125930 176704
rect 128174 176760 128230 176769
rect 128174 176695 128230 176704
rect 133142 176760 133198 176769
rect 133142 176695 133198 176704
rect 136086 176760 136142 176769
rect 136086 176695 136088 176704
rect 136140 176695 136142 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 158994 176760 159050 176769
rect 158994 176695 158996 176704
rect 136088 176666 136140 176672
rect 159048 176695 159050 176704
rect 158996 176666 159048 176672
rect 134432 176248 134484 176254
rect 134432 176190 134484 176196
rect 121920 176180 121972 176186
rect 121920 176122 121972 176128
rect 116952 176112 117004 176118
rect 116952 176054 117004 176060
rect 115756 175976 115808 175982
rect 115756 175918 115808 175924
rect 115768 175001 115796 175918
rect 116964 175409 116992 176054
rect 120816 176044 120868 176050
rect 120816 175986 120868 175992
rect 120828 175409 120856 175986
rect 121932 175409 121960 176122
rect 134444 175409 134472 176190
rect 116950 175400 117006 175409
rect 116950 175335 117006 175344
rect 120814 175400 120870 175409
rect 120814 175335 120870 175344
rect 121918 175400 121974 175409
rect 121918 175335 121974 175344
rect 134430 175400 134486 175409
rect 134430 175335 134486 175344
rect 115754 174992 115810 175001
rect 115754 174927 115810 174936
rect 165356 173233 165384 176938
rect 165436 176724 165488 176730
rect 165436 176666 165488 176672
rect 165448 174554 165476 176666
rect 165528 176248 165580 176254
rect 165528 176190 165580 176196
rect 165540 175234 165568 176190
rect 165528 175228 165580 175234
rect 165528 175170 165580 175176
rect 165436 174548 165488 174554
rect 165436 174490 165488 174496
rect 165342 173224 165398 173233
rect 165342 173159 165398 173168
rect 166276 158710 166304 180950
rect 166356 178356 166408 178362
rect 166356 178298 166408 178304
rect 166368 166870 166396 178298
rect 166448 176180 166500 176186
rect 166448 176122 166500 176128
rect 166460 168366 166488 176122
rect 166552 173874 166580 181086
rect 166540 173868 166592 173874
rect 166540 173810 166592 173816
rect 166448 168360 166500 168366
rect 166448 168302 166500 168308
rect 166356 166864 166408 166870
rect 166356 166806 166408 166812
rect 167656 160070 167684 182242
rect 167828 181076 167880 181082
rect 167828 181018 167880 181024
rect 167734 177032 167790 177041
rect 167734 176967 167790 176976
rect 167748 160750 167776 176967
rect 167840 169726 167868 181018
rect 168010 171592 168066 171601
rect 168010 171527 168066 171536
rect 168024 169794 168052 171527
rect 168012 169788 168064 169794
rect 168012 169730 168064 169736
rect 167828 169720 167880 169726
rect 167828 169662 167880 169668
rect 169036 161430 169064 182310
rect 169208 179648 169260 179654
rect 169208 179590 169260 179596
rect 169116 178288 169168 178294
rect 169116 178230 169168 178236
rect 169128 162858 169156 178230
rect 169220 169658 169248 179590
rect 170496 176860 170548 176866
rect 170496 176802 170548 176808
rect 169300 176112 169352 176118
rect 169300 176054 169352 176060
rect 169208 169652 169260 169658
rect 169208 169594 169260 169600
rect 169312 166938 169340 176054
rect 170404 169788 170456 169794
rect 170404 169730 170456 169736
rect 169300 166932 169352 166938
rect 169300 166874 169352 166880
rect 169116 162852 169168 162858
rect 169116 162794 169168 162800
rect 169024 161424 169076 161430
rect 169024 161366 169076 161372
rect 167736 160744 167788 160750
rect 167736 160686 167788 160692
rect 167644 160064 167696 160070
rect 167644 160006 167696 160012
rect 166264 158704 166316 158710
rect 166264 158646 166316 158652
rect 169024 153264 169076 153270
rect 169024 153206 169076 153212
rect 166264 147688 166316 147694
rect 166264 147630 166316 147636
rect 66074 129296 66130 129305
rect 66074 129231 66130 129240
rect 65154 126304 65210 126313
rect 65154 126239 65210 126248
rect 65168 125662 65196 126239
rect 63408 125656 63460 125662
rect 63408 125598 63460 125604
rect 65156 125656 65208 125662
rect 65156 125598 65208 125604
rect 63420 95062 63448 125598
rect 65982 123584 66038 123593
rect 65982 123519 66038 123528
rect 64786 102232 64842 102241
rect 64786 102167 64842 102176
rect 63408 95056 63460 95062
rect 63408 94998 63460 95004
rect 64800 85542 64828 102167
rect 65996 90953 66024 123519
rect 66088 94897 66116 129231
rect 66166 128072 66222 128081
rect 66166 128007 66222 128016
rect 66074 94888 66130 94897
rect 66074 94823 66130 94832
rect 66180 93809 66208 128007
rect 67638 125216 67694 125225
rect 67638 125151 67694 125160
rect 67546 122632 67602 122641
rect 67546 122567 67602 122576
rect 67454 120864 67510 120873
rect 67454 120799 67510 120808
rect 66166 93800 66222 93809
rect 66166 93735 66222 93744
rect 65982 90944 66038 90953
rect 65982 90879 66038 90888
rect 67468 89690 67496 120799
rect 67456 89684 67508 89690
rect 67456 89626 67508 89632
rect 64788 85536 64840 85542
rect 64788 85478 64840 85484
rect 67560 77246 67588 122567
rect 67652 91089 67680 125151
rect 67730 100736 67786 100745
rect 67730 100671 67786 100680
rect 67638 91080 67694 91089
rect 67638 91015 67694 91024
rect 67744 88233 67772 100671
rect 164884 99408 164936 99414
rect 164884 99350 164936 99356
rect 105726 94752 105782 94761
rect 105726 94687 105782 94696
rect 112350 94752 112406 94761
rect 112350 94687 112406 94696
rect 128082 94752 128138 94761
rect 128082 94687 128138 94696
rect 151726 94752 151782 94761
rect 151726 94687 151782 94696
rect 105740 93906 105768 94687
rect 106462 94072 106518 94081
rect 106462 94007 106518 94016
rect 105728 93900 105780 93906
rect 105728 93842 105780 93848
rect 88982 93528 89038 93537
rect 88982 93463 89038 93472
rect 88996 93294 89024 93463
rect 88984 93288 89036 93294
rect 88984 93230 89036 93236
rect 103426 93256 103482 93265
rect 103426 93191 103482 93200
rect 86590 92440 86646 92449
rect 86590 92375 86646 92384
rect 98550 92440 98606 92449
rect 98550 92375 98552 92384
rect 75826 91216 75882 91225
rect 75826 91151 75882 91160
rect 84658 91216 84714 91225
rect 84658 91151 84714 91160
rect 67730 88224 67786 88233
rect 67730 88159 67786 88168
rect 75840 82822 75868 91151
rect 84672 88330 84700 91151
rect 86604 91118 86632 92375
rect 98604 92375 98606 92384
rect 98552 92346 98604 92352
rect 90362 91760 90418 91769
rect 90362 91695 90418 91704
rect 86866 91216 86922 91225
rect 86866 91151 86922 91160
rect 86592 91112 86644 91118
rect 86592 91054 86644 91060
rect 84660 88324 84712 88330
rect 84660 88266 84712 88272
rect 86880 84046 86908 91151
rect 90376 89622 90404 91695
rect 101862 91488 101918 91497
rect 101862 91423 101918 91432
rect 95054 91352 95110 91361
rect 95054 91287 95110 91296
rect 99194 91352 99250 91361
rect 99194 91287 99250 91296
rect 100574 91352 100630 91361
rect 100574 91287 100630 91296
rect 92294 91216 92350 91225
rect 92294 91151 92350 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 90364 89616 90416 89622
rect 90364 89558 90416 89564
rect 92308 85338 92336 91151
rect 92296 85332 92348 85338
rect 92296 85274 92348 85280
rect 86868 84040 86920 84046
rect 86868 83982 86920 83988
rect 75828 82816 75880 82822
rect 75828 82758 75880 82764
rect 93780 80034 93808 91151
rect 95068 81394 95096 91287
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 97078 91216 97134 91225
rect 97078 91151 97134 91160
rect 97906 91216 97962 91225
rect 97906 91151 97962 91160
rect 95056 81388 95108 81394
rect 95056 81330 95108 81336
rect 93768 80028 93820 80034
rect 93768 79970 93820 79976
rect 95160 78674 95188 91151
rect 96540 83978 96568 91151
rect 97092 86834 97120 91151
rect 97080 86828 97132 86834
rect 97080 86770 97132 86776
rect 96528 83972 96580 83978
rect 96528 83914 96580 83920
rect 95148 78668 95200 78674
rect 95148 78610 95200 78616
rect 67548 77240 67600 77246
rect 67548 77182 67600 77188
rect 97920 77178 97948 91151
rect 99208 82793 99236 91287
rect 99286 91216 99342 91225
rect 99286 91151 99342 91160
rect 99194 82784 99250 82793
rect 99194 82719 99250 82728
rect 99300 78538 99328 91151
rect 100588 88262 100616 91287
rect 100666 91216 100722 91225
rect 100666 91151 100722 91160
rect 100576 88256 100628 88262
rect 100576 88198 100628 88204
rect 100680 79830 100708 91151
rect 101876 86970 101904 91423
rect 101954 91352 102010 91361
rect 101954 91287 102010 91296
rect 101864 86964 101916 86970
rect 101864 86906 101916 86912
rect 101968 81433 101996 91287
rect 102046 91216 102102 91225
rect 102046 91151 102102 91160
rect 103058 91216 103114 91225
rect 103058 91151 103114 91160
rect 101954 81424 102010 81433
rect 101954 81359 102010 81368
rect 100668 79824 100720 79830
rect 100668 79766 100720 79772
rect 99288 78532 99340 78538
rect 99288 78474 99340 78480
rect 102060 78470 102088 91151
rect 103072 85406 103100 91151
rect 103060 85400 103112 85406
rect 103060 85342 103112 85348
rect 103440 82686 103468 93191
rect 106476 93158 106504 94007
rect 112364 93974 112392 94687
rect 122840 94512 122892 94518
rect 122840 94454 122892 94460
rect 112352 93968 112404 93974
rect 112352 93910 112404 93916
rect 121734 93664 121790 93673
rect 121734 93599 121790 93608
rect 111246 93528 111302 93537
rect 111246 93463 111302 93472
rect 110142 93256 110198 93265
rect 111260 93226 111288 93463
rect 121748 93362 121776 93599
rect 121736 93356 121788 93362
rect 121736 93298 121788 93304
rect 110142 93191 110198 93200
rect 111248 93220 111300 93226
rect 106464 93152 106516 93158
rect 106464 93094 106516 93100
rect 104346 92440 104402 92449
rect 104346 92375 104402 92384
rect 104622 92440 104678 92449
rect 104622 92375 104678 92384
rect 106646 92440 106702 92449
rect 106646 92375 106702 92384
rect 104360 91050 104388 92375
rect 104636 91186 104664 92375
rect 106660 92070 106688 92375
rect 106648 92064 106700 92070
rect 106648 92006 106700 92012
rect 106002 91624 106058 91633
rect 106002 91559 106058 91568
rect 104624 91180 104676 91186
rect 104624 91122 104676 91128
rect 104348 91044 104400 91050
rect 104348 90986 104400 90992
rect 106016 89486 106044 91559
rect 109498 91488 109554 91497
rect 109498 91423 109554 91432
rect 108854 91352 108910 91361
rect 108854 91287 108910 91296
rect 106004 89480 106056 89486
rect 106004 89422 106056 89428
rect 108868 84182 108896 91287
rect 108946 91216 109002 91225
rect 108946 91151 109002 91160
rect 108856 84176 108908 84182
rect 108856 84118 108908 84124
rect 103428 82680 103480 82686
rect 103428 82622 103480 82628
rect 108960 79762 108988 91151
rect 109512 86766 109540 91423
rect 110156 90914 110184 93191
rect 111248 93162 111300 93168
rect 110694 92440 110750 92449
rect 110694 92375 110750 92384
rect 118054 92440 118110 92449
rect 118054 92375 118110 92384
rect 110708 92274 110736 92375
rect 118068 92342 118096 92375
rect 118056 92336 118108 92342
rect 118056 92278 118108 92284
rect 122852 92274 122880 94454
rect 128096 94042 128124 94687
rect 128084 94036 128136 94042
rect 128084 93978 128136 93984
rect 134430 93528 134486 93537
rect 151740 93498 151768 94687
rect 134430 93463 134486 93472
rect 151728 93492 151780 93498
rect 134444 93430 134472 93463
rect 151728 93434 151780 93440
rect 134432 93424 134484 93430
rect 134432 93366 134484 93372
rect 164896 93294 164924 99350
rect 164884 93288 164936 93294
rect 164884 93230 164936 93236
rect 126702 92440 126758 92449
rect 126702 92375 126758 92384
rect 133142 92440 133198 92449
rect 133142 92375 133198 92384
rect 151542 92440 151598 92449
rect 151542 92375 151598 92384
rect 126716 92274 126744 92375
rect 110696 92268 110748 92274
rect 110696 92210 110748 92216
rect 122840 92268 122892 92274
rect 122840 92210 122892 92216
rect 126704 92268 126756 92274
rect 126704 92210 126756 92216
rect 133156 92206 133184 92375
rect 133144 92200 133196 92206
rect 133144 92142 133196 92148
rect 151556 92138 151584 92375
rect 151544 92132 151596 92138
rect 151544 92074 151596 92080
rect 115478 92032 115534 92041
rect 115478 91967 115534 91976
rect 126518 92032 126574 92041
rect 126518 91967 126574 91976
rect 151358 92032 151414 92041
rect 151358 91967 151414 91976
rect 114374 91352 114430 91361
rect 114374 91287 114430 91296
rect 110326 91216 110382 91225
rect 110326 91151 110382 91160
rect 113086 91216 113142 91225
rect 113086 91151 113142 91160
rect 110144 90908 110196 90914
rect 110144 90850 110196 90856
rect 109500 86760 109552 86766
rect 109500 86702 109552 86708
rect 108948 79756 109000 79762
rect 108948 79698 109000 79704
rect 110340 78606 110368 91151
rect 110420 91112 110472 91118
rect 110420 91054 110472 91060
rect 110432 86902 110460 91054
rect 110420 86896 110472 86902
rect 110420 86838 110472 86844
rect 113100 81297 113128 91151
rect 114388 85474 114416 91287
rect 114466 91216 114522 91225
rect 114466 91151 114522 91160
rect 114376 85468 114428 85474
rect 114376 85410 114428 85416
rect 114480 82754 114508 91151
rect 115492 89729 115520 91967
rect 119894 91760 119950 91769
rect 119894 91695 119950 91704
rect 117134 91352 117190 91361
rect 117134 91287 117190 91296
rect 115570 91216 115626 91225
rect 115570 91151 115626 91160
rect 115846 91216 115902 91225
rect 115846 91151 115902 91160
rect 115478 89720 115534 89729
rect 115478 89655 115534 89664
rect 115584 88126 115612 91151
rect 115572 88120 115624 88126
rect 115572 88062 115624 88068
rect 115860 83910 115888 91151
rect 117148 88194 117176 91287
rect 117226 91216 117282 91225
rect 118606 91216 118662 91225
rect 117226 91151 117282 91160
rect 117964 91180 118016 91186
rect 117136 88188 117188 88194
rect 117136 88130 117188 88136
rect 115848 83904 115900 83910
rect 115848 83846 115900 83852
rect 114468 82748 114520 82754
rect 114468 82690 114520 82696
rect 113086 81288 113142 81297
rect 113086 81223 113142 81232
rect 117240 79966 117268 91151
rect 118606 91151 118662 91160
rect 117964 91122 118016 91128
rect 117228 79960 117280 79966
rect 117228 79902 117280 79908
rect 110328 78600 110380 78606
rect 110328 78542 110380 78548
rect 102048 78464 102100 78470
rect 102048 78406 102100 78412
rect 97908 77172 97960 77178
rect 97908 77114 97960 77120
rect 95240 75268 95292 75274
rect 95240 75210 95292 75216
rect 75920 75200 75972 75206
rect 75920 75142 75972 75148
rect 70398 72448 70454 72457
rect 70398 72383 70454 72392
rect 52460 68332 52512 68338
rect 52460 68274 52512 68280
rect 43444 59356 43496 59362
rect 43444 59298 43496 59304
rect 43536 58676 43588 58682
rect 43536 58618 43588 58624
rect 42798 46200 42854 46209
rect 42798 46135 42854 46144
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 36832 354 36860 3470
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 46135
rect 43548 3466 43576 58618
rect 48320 29640 48372 29646
rect 48320 29582 48372 29588
rect 44178 22672 44234 22681
rect 44178 22607 44234 22616
rect 44192 6914 44220 22607
rect 44272 20052 44324 20058
rect 44272 19994 44324 20000
rect 44284 16574 44312 19994
rect 45558 17232 45614 17241
rect 45558 17167 45614 17176
rect 45572 16574 45600 17167
rect 48332 16574 48360 29582
rect 44284 16546 45048 16574
rect 45572 16546 46704 16574
rect 48332 16546 48544 16574
rect 44192 6886 44312 6914
rect 43536 3460 43588 3466
rect 43536 3402 43588 3408
rect 44284 480 44312 6886
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 47860 6180 47912 6186
rect 47860 6122 47912 6128
rect 47872 480 47900 6122
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48516 354 48544 16546
rect 51356 8968 51408 8974
rect 51356 8910 51408 8916
rect 50160 3460 50212 3466
rect 50160 3402 50212 3408
rect 50172 480 50200 3402
rect 51368 480 51396 8910
rect 52472 3534 52500 68274
rect 64880 61464 64932 61470
rect 64880 61406 64932 61412
rect 55220 54528 55272 54534
rect 55220 54470 55272 54476
rect 53840 32428 53892 32434
rect 53840 32370 53892 32376
rect 52552 31136 52604 31142
rect 52552 31078 52604 31084
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 52564 480 52592 31078
rect 53852 16574 53880 32370
rect 55232 16574 55260 54470
rect 62118 51776 62174 51785
rect 62118 51711 62174 51720
rect 56600 43444 56652 43450
rect 56600 43386 56652 43392
rect 56612 16574 56640 43386
rect 60740 37936 60792 37942
rect 60740 37878 60792 37884
rect 59360 31068 59412 31074
rect 59360 31010 59412 31016
rect 57980 26988 58032 26994
rect 57980 26930 58032 26936
rect 57992 16574 58020 26930
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 53380 3528 53432 3534
rect 53380 3470 53432 3476
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3470
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 31010
rect 60752 16574 60780 37878
rect 62132 16574 62160 51711
rect 63500 40724 63552 40730
rect 63500 40666 63552 40672
rect 63512 16574 63540 40666
rect 64892 16574 64920 61406
rect 66260 50448 66312 50454
rect 66260 50390 66312 50396
rect 66272 16574 66300 50390
rect 69020 49088 69072 49094
rect 69020 49030 69072 49036
rect 67640 39432 67692 39438
rect 67640 39374 67692 39380
rect 60752 16546 60872 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 60844 480 60872 16546
rect 61568 13116 61620 13122
rect 61568 13058 61620 13064
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 13058
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 39374
rect 69032 3534 69060 49030
rect 70412 16574 70440 72383
rect 74540 69760 74592 69766
rect 74540 69702 74592 69708
rect 74552 16574 74580 69702
rect 70412 16546 71544 16574
rect 74552 16546 75040 16574
rect 69112 14476 69164 14482
rect 69112 14418 69164 14424
rect 69020 3528 69072 3534
rect 69020 3470 69072 3476
rect 69124 480 69152 14418
rect 69940 3528 69992 3534
rect 69940 3470 69992 3476
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3470
rect 71516 480 71544 16546
rect 72608 6248 72660 6254
rect 72608 6190 72660 6196
rect 72620 480 72648 6190
rect 73804 4820 73856 4826
rect 73804 4762 73856 4768
rect 73816 480 73844 4762
rect 75012 480 75040 16546
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 75142
rect 78680 73840 78732 73846
rect 78680 73782 78732 73788
rect 77298 47560 77354 47569
rect 77298 47495 77354 47504
rect 77312 16574 77340 47495
rect 78692 16574 78720 73782
rect 82820 60104 82872 60110
rect 82820 60046 82872 60052
rect 81440 36576 81492 36582
rect 81440 36518 81492 36524
rect 80060 29708 80112 29714
rect 80060 29650 80112 29656
rect 80072 16574 80100 29650
rect 81452 16574 81480 36518
rect 82832 16574 82860 60046
rect 93860 57248 93912 57254
rect 93860 57190 93912 57196
rect 86960 35284 87012 35290
rect 86960 35226 87012 35232
rect 85580 32496 85632 32502
rect 85580 32438 85632 32444
rect 84200 17264 84252 17270
rect 84200 17206 84252 17212
rect 77312 16546 77432 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77404 480 77432 16546
rect 78588 9036 78640 9042
rect 78588 8978 78640 8984
rect 78600 480 78628 8978
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 17206
rect 85592 6914 85620 32438
rect 85672 18692 85724 18698
rect 85672 18634 85724 18640
rect 85684 16574 85712 18634
rect 86972 16574 87000 35226
rect 88340 28348 88392 28354
rect 88340 28290 88392 28296
rect 88352 16574 88380 28290
rect 92480 22772 92532 22778
rect 92480 22714 92532 22720
rect 91100 21480 91152 21486
rect 91100 21422 91152 21428
rect 91112 16574 91140 21422
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 91112 16546 91600 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 90364 7608 90416 7614
rect 90364 7550 90416 7556
rect 90376 480 90404 7550
rect 91572 480 91600 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 22714
rect 93872 16574 93900 57190
rect 95252 16574 95280 75210
rect 117976 74526 118004 91122
rect 118620 81326 118648 91151
rect 119908 89554 119936 91695
rect 124126 91488 124182 91497
rect 124126 91423 124182 91432
rect 120814 91352 120870 91361
rect 120814 91287 120870 91296
rect 119896 89548 119948 89554
rect 119896 89490 119948 89496
rect 120828 86698 120856 91287
rect 121366 91216 121422 91225
rect 121366 91151 121422 91160
rect 123758 91216 123814 91225
rect 123758 91151 123814 91160
rect 124034 91216 124090 91225
rect 124034 91151 124090 91160
rect 120816 86692 120868 86698
rect 120816 86634 120868 86640
rect 121380 84114 121408 91151
rect 123772 88058 123800 91151
rect 123760 88052 123812 88058
rect 123760 87994 123812 88000
rect 124048 87990 124076 91151
rect 124036 87984 124088 87990
rect 124036 87926 124088 87932
rect 121368 84108 121420 84114
rect 121368 84050 121420 84056
rect 118608 81320 118660 81326
rect 118608 81262 118660 81268
rect 124140 79898 124168 91423
rect 125414 91352 125470 91361
rect 125414 91287 125470 91296
rect 125428 85202 125456 91287
rect 125506 91216 125562 91225
rect 125506 91151 125562 91160
rect 125416 85196 125468 85202
rect 125416 85138 125468 85144
rect 125520 82618 125548 91151
rect 126532 90982 126560 91967
rect 132406 91624 132462 91633
rect 132406 91559 132462 91568
rect 126702 91216 126758 91225
rect 126702 91151 126758 91160
rect 129646 91216 129702 91225
rect 129646 91151 129702 91160
rect 130750 91216 130806 91225
rect 130750 91151 130806 91160
rect 126520 90976 126572 90982
rect 126520 90918 126572 90924
rect 126716 86873 126744 91151
rect 126702 86864 126758 86873
rect 126702 86799 126758 86808
rect 125508 82612 125560 82618
rect 125508 82554 125560 82560
rect 129660 81258 129688 91151
rect 130764 85513 130792 91151
rect 132420 89418 132448 91559
rect 136546 91216 136602 91225
rect 136546 91151 136602 91160
rect 132408 89412 132460 89418
rect 132408 89354 132460 89360
rect 130750 85504 130806 85513
rect 130750 85439 130806 85448
rect 136560 83842 136588 91151
rect 151372 90846 151400 91967
rect 152646 91216 152702 91225
rect 152646 91151 152702 91160
rect 151360 90840 151412 90846
rect 151360 90782 151412 90788
rect 152660 85270 152688 91151
rect 152648 85264 152700 85270
rect 152648 85206 152700 85212
rect 166276 83842 166304 147630
rect 167644 125656 167696 125662
rect 167644 125598 167696 125604
rect 166356 122868 166408 122874
rect 166356 122810 166408 122816
rect 166368 93362 166396 122810
rect 166448 111852 166500 111858
rect 166448 111794 166500 111800
rect 166356 93356 166408 93362
rect 166356 93298 166408 93304
rect 166460 88262 166488 111794
rect 167460 110424 167512 110430
rect 167460 110366 167512 110372
rect 167472 110129 167500 110366
rect 167458 110120 167514 110129
rect 167458 110055 167514 110064
rect 166540 98048 166592 98054
rect 166540 97990 166592 97996
rect 166448 88256 166500 88262
rect 166448 88198 166500 88204
rect 166552 84046 166580 97990
rect 167656 85202 167684 125598
rect 167736 124228 167788 124234
rect 167736 124170 167788 124176
rect 167748 87990 167776 124170
rect 167920 122120 167972 122126
rect 167920 122062 167972 122068
rect 167828 113212 167880 113218
rect 167828 113154 167880 113160
rect 167840 91050 167868 113154
rect 167932 111761 167960 122062
rect 167918 111752 167974 111761
rect 167918 111687 167974 111696
rect 167920 108996 167972 109002
rect 167920 108938 167972 108944
rect 167932 108769 167960 108938
rect 167918 108760 167974 108769
rect 167918 108695 167974 108704
rect 167920 101448 167972 101454
rect 167920 101390 167972 101396
rect 167932 92206 167960 101390
rect 169036 93498 169064 153206
rect 170416 150414 170444 169730
rect 170508 160002 170536 176802
rect 170600 171086 170628 182378
rect 179340 181529 179368 273799
rect 179326 181520 179382 181529
rect 179326 181455 179382 181464
rect 178684 180940 178736 180946
rect 178684 180882 178736 180888
rect 173164 179580 173216 179586
rect 173164 179522 173216 179528
rect 170588 171080 170640 171086
rect 170588 171022 170640 171028
rect 170496 159996 170548 160002
rect 170496 159938 170548 159944
rect 173176 155922 173204 179522
rect 177304 178220 177356 178226
rect 177304 178162 177356 178168
rect 177316 164218 177344 178162
rect 178696 165578 178724 180882
rect 180536 180470 180564 295326
rect 180616 251252 180668 251258
rect 180616 251194 180668 251200
rect 180524 180464 180576 180470
rect 180524 180406 180576 180412
rect 180064 176044 180116 176050
rect 180064 175986 180116 175992
rect 180076 168298 180104 175986
rect 180064 168292 180116 168298
rect 180064 168234 180116 168240
rect 178684 165572 178736 165578
rect 178684 165514 178736 165520
rect 177304 164212 177356 164218
rect 177304 164154 177356 164160
rect 173164 155916 173216 155922
rect 173164 155858 173216 155864
rect 180064 153332 180116 153338
rect 180064 153274 180116 153280
rect 177396 151836 177448 151842
rect 177396 151778 177448 151784
rect 170496 150476 170548 150482
rect 170496 150418 170548 150424
rect 170404 150408 170456 150414
rect 170404 150350 170456 150356
rect 170404 140820 170456 140826
rect 170404 140762 170456 140768
rect 169116 118856 169168 118862
rect 169116 118798 169168 118804
rect 169024 93492 169076 93498
rect 169024 93434 169076 93440
rect 167920 92200 167972 92206
rect 167920 92142 167972 92148
rect 167828 91044 167880 91050
rect 167828 90986 167880 90992
rect 169128 88126 169156 118798
rect 169208 117360 169260 117366
rect 169208 117302 169260 117308
rect 169220 90914 169248 117302
rect 169300 105052 169352 105058
rect 169300 104994 169352 105000
rect 169208 90908 169260 90914
rect 169208 90850 169260 90856
rect 169312 89622 169340 104994
rect 169300 89616 169352 89622
rect 169300 89558 169352 89564
rect 169116 88120 169168 88126
rect 169116 88062 169168 88068
rect 167736 87984 167788 87990
rect 167736 87926 167788 87932
rect 167644 85196 167696 85202
rect 167644 85138 167696 85144
rect 166540 84040 166592 84046
rect 166540 83982 166592 83988
rect 136548 83836 136600 83842
rect 136548 83778 136600 83784
rect 166264 83836 166316 83842
rect 166264 83778 166316 83784
rect 170416 82618 170444 140762
rect 170508 110430 170536 150418
rect 174544 146328 174596 146334
rect 174544 146270 174596 146276
rect 171876 143608 171928 143614
rect 171876 143550 171928 143556
rect 171784 132524 171836 132530
rect 171784 132466 171836 132472
rect 170588 122936 170640 122942
rect 170588 122878 170640 122884
rect 170496 110424 170548 110430
rect 170496 110366 170548 110372
rect 170496 106344 170548 106350
rect 170496 106286 170548 106292
rect 170508 85338 170536 106286
rect 170600 86698 170628 122878
rect 170680 120148 170732 120154
rect 170680 120090 170732 120096
rect 170692 88194 170720 120090
rect 170680 88188 170732 88194
rect 170680 88130 170732 88136
rect 170588 86692 170640 86698
rect 170588 86634 170640 86640
rect 170496 85332 170548 85338
rect 170496 85274 170548 85280
rect 170404 82612 170456 82618
rect 170404 82554 170456 82560
rect 129648 81252 129700 81258
rect 129648 81194 129700 81200
rect 124128 79892 124180 79898
rect 124128 79834 124180 79840
rect 171796 79762 171824 132466
rect 171888 94042 171916 143550
rect 171968 138032 172020 138038
rect 171968 137974 172020 137980
rect 171876 94036 171928 94042
rect 171876 93978 171928 93984
rect 171980 93673 172008 137974
rect 173348 134564 173400 134570
rect 173348 134506 173400 134512
rect 172060 114572 172112 114578
rect 172060 114514 172112 114520
rect 171966 93664 172022 93673
rect 171966 93599 172022 93608
rect 172072 89486 172100 114514
rect 173256 110492 173308 110498
rect 173256 110434 173308 110440
rect 173164 109064 173216 109070
rect 173164 109006 173216 109012
rect 172060 89480 172112 89486
rect 172060 89422 172112 89428
rect 171784 79756 171836 79762
rect 171784 79698 171836 79704
rect 173176 77178 173204 109006
rect 173268 79830 173296 110434
rect 173360 109002 173388 134506
rect 173440 118788 173492 118794
rect 173440 118730 173492 118736
rect 173348 108996 173400 109002
rect 173348 108938 173400 108944
rect 173452 93974 173480 118730
rect 173440 93968 173492 93974
rect 173440 93910 173492 93916
rect 174556 93430 174584 146270
rect 177304 143676 177356 143682
rect 177304 143618 177356 143624
rect 175924 140888 175976 140894
rect 175924 140830 175976 140836
rect 174636 129804 174688 129810
rect 174636 129746 174688 129752
rect 174544 93424 174596 93430
rect 174544 93366 174596 93372
rect 173256 79824 173308 79830
rect 173256 79766 173308 79772
rect 174648 78470 174676 129746
rect 174728 127016 174780 127022
rect 174728 126958 174780 126964
rect 174740 86834 174768 126958
rect 175936 88058 175964 140830
rect 176016 129872 176068 129878
rect 176016 129814 176068 129820
rect 175924 88052 175976 88058
rect 175924 87994 175976 88000
rect 174728 86828 174780 86834
rect 174728 86770 174780 86776
rect 176028 82686 176056 129814
rect 176108 109132 176160 109138
rect 176108 109074 176160 109080
rect 176120 83978 176148 109074
rect 176108 83972 176160 83978
rect 176108 83914 176160 83920
rect 176016 82680 176068 82686
rect 176016 82622 176068 82628
rect 177316 81258 177344 143618
rect 177408 90846 177436 151778
rect 178684 144968 178736 144974
rect 178684 144910 178736 144916
rect 177488 128376 177540 128382
rect 177488 128318 177540 128324
rect 177396 90840 177448 90846
rect 177396 90782 177448 90788
rect 177304 81252 177356 81258
rect 177304 81194 177356 81200
rect 177500 78538 177528 128318
rect 178696 89418 178724 144910
rect 178776 120216 178828 120222
rect 178776 120158 178828 120164
rect 178684 89412 178736 89418
rect 178684 89354 178736 89360
rect 178788 83910 178816 120158
rect 180076 92138 180104 153274
rect 180156 116000 180208 116006
rect 180156 115942 180208 115948
rect 180064 92132 180116 92138
rect 180064 92074 180116 92080
rect 180168 86766 180196 115942
rect 180628 92478 180656 251194
rect 180720 248402 180748 697546
rect 182088 287088 182140 287094
rect 182088 287030 182140 287036
rect 181996 251320 182048 251326
rect 181996 251262 182048 251268
rect 180708 248396 180760 248402
rect 180708 248338 180760 248344
rect 182008 195294 182036 251262
rect 181996 195288 182048 195294
rect 181996 195230 182048 195236
rect 182100 178809 182128 287030
rect 183468 280220 183520 280226
rect 183468 280162 183520 280168
rect 182086 178800 182142 178809
rect 182086 178735 182142 178744
rect 183480 176050 183508 280162
rect 184756 274712 184808 274718
rect 184756 274654 184808 274660
rect 184664 256828 184716 256834
rect 184664 256770 184716 256776
rect 184676 188358 184704 256770
rect 184664 188352 184716 188358
rect 184664 188294 184716 188300
rect 184768 185706 184796 274654
rect 184860 255270 184888 700266
rect 195244 698964 195296 698970
rect 195244 698906 195296 698912
rect 188344 632732 188396 632738
rect 188344 632674 188396 632680
rect 186228 288448 186280 288454
rect 186228 288390 186280 288396
rect 186136 269136 186188 269142
rect 186136 269078 186188 269084
rect 184848 255264 184900 255270
rect 184848 255206 184900 255212
rect 184756 185700 184808 185706
rect 184756 185642 184808 185648
rect 186148 178673 186176 269078
rect 186240 185842 186268 288390
rect 187424 277432 187476 277438
rect 187424 277374 187476 277380
rect 187332 250504 187384 250510
rect 187332 250446 187384 250452
rect 186228 185836 186280 185842
rect 186228 185778 186280 185784
rect 187344 182986 187372 250446
rect 187332 182980 187384 182986
rect 187332 182922 187384 182928
rect 187436 180334 187464 277374
rect 187516 274780 187568 274786
rect 187516 274722 187568 274728
rect 187424 180328 187476 180334
rect 187424 180270 187476 180276
rect 186134 178664 186190 178673
rect 186134 178599 186190 178608
rect 187528 176118 187556 274722
rect 188356 267646 188384 632674
rect 193128 295452 193180 295458
rect 193128 295394 193180 295400
rect 188988 289876 189040 289882
rect 188988 289818 189040 289824
rect 188896 284368 188948 284374
rect 188896 284310 188948 284316
rect 188344 267640 188396 267646
rect 188344 267582 188396 267588
rect 187608 264988 187660 264994
rect 187608 264930 187660 264936
rect 187516 176112 187568 176118
rect 187516 176054 187568 176060
rect 183468 176044 183520 176050
rect 183468 175986 183520 175992
rect 184204 132592 184256 132598
rect 184204 132534 184256 132540
rect 180616 92472 180668 92478
rect 180616 92414 180668 92420
rect 184216 92070 184244 132534
rect 186964 131164 187016 131170
rect 186964 131106 187016 131112
rect 184296 100768 184348 100774
rect 184296 100710 184348 100716
rect 184204 92064 184256 92070
rect 184204 92006 184256 92012
rect 184308 88330 184336 100710
rect 186976 93906 187004 131106
rect 187056 113280 187108 113286
rect 187056 113222 187108 113228
rect 186964 93900 187016 93906
rect 186964 93842 187016 93848
rect 184296 88324 184348 88330
rect 184296 88266 184348 88272
rect 180156 86760 180208 86766
rect 180156 86702 180208 86708
rect 187068 85406 187096 113222
rect 187620 95198 187648 264930
rect 188712 263696 188764 263702
rect 188712 263638 188764 263644
rect 188724 233918 188752 263638
rect 188804 258120 188856 258126
rect 188804 258062 188856 258068
rect 188712 233912 188764 233918
rect 188712 233854 188764 233860
rect 188816 180198 188844 258062
rect 188908 193186 188936 284310
rect 188896 193180 188948 193186
rect 188896 193122 188948 193128
rect 189000 183054 189028 289818
rect 190368 287156 190420 287162
rect 190368 287098 190420 287104
rect 190092 277500 190144 277506
rect 190092 277442 190144 277448
rect 190104 228478 190132 277442
rect 190276 276072 190328 276078
rect 190276 276014 190328 276020
rect 190184 241528 190236 241534
rect 190184 241470 190236 241476
rect 190092 228472 190144 228478
rect 190092 228414 190144 228420
rect 188988 183048 189040 183054
rect 188988 182990 189040 182996
rect 190196 180402 190224 241470
rect 190288 185910 190316 276014
rect 190276 185904 190328 185910
rect 190276 185846 190328 185852
rect 190184 180396 190236 180402
rect 190184 180338 190236 180344
rect 188804 180192 188856 180198
rect 188804 180134 188856 180140
rect 190380 177313 190408 287098
rect 192852 270564 192904 270570
rect 192852 270506 192904 270512
rect 191656 262268 191708 262274
rect 191656 262210 191708 262216
rect 191564 249824 191616 249830
rect 191564 249766 191616 249772
rect 191104 244928 191156 244934
rect 191104 244870 191156 244876
rect 190550 240136 190606 240145
rect 190550 240071 190606 240080
rect 190564 239902 190592 240071
rect 190552 239896 190604 239902
rect 190552 239838 190604 239844
rect 191116 238678 191144 244870
rect 191104 238672 191156 238678
rect 191104 238614 191156 238620
rect 191104 232620 191156 232626
rect 191104 232562 191156 232568
rect 190366 177304 190422 177313
rect 190366 177239 190422 177248
rect 188344 142180 188396 142186
rect 188344 142122 188396 142128
rect 187608 95192 187660 95198
rect 187608 95134 187660 95140
rect 188356 92274 188384 142122
rect 188436 125724 188488 125730
rect 188436 125666 188488 125672
rect 188344 92268 188396 92274
rect 188344 92210 188396 92216
rect 188448 90982 188476 125666
rect 188436 90976 188488 90982
rect 188436 90918 188488 90924
rect 188344 90364 188396 90370
rect 188344 90306 188396 90312
rect 187056 85400 187108 85406
rect 187056 85342 187108 85348
rect 178776 83904 178828 83910
rect 178776 83846 178828 83852
rect 177488 78532 177540 78538
rect 177488 78474 177540 78480
rect 174636 78464 174688 78470
rect 174636 78406 174688 78412
rect 173164 77172 173216 77178
rect 173164 77114 173216 77120
rect 125600 75336 125652 75342
rect 125600 75278 125652 75284
rect 117964 74520 118016 74526
rect 117964 74462 118016 74468
rect 99380 73908 99432 73914
rect 99380 73850 99432 73856
rect 96620 72480 96672 72486
rect 96620 72422 96672 72428
rect 96632 16574 96660 72422
rect 98000 54596 98052 54602
rect 98000 54538 98052 54544
rect 98012 16574 98040 54538
rect 99392 16574 99420 73850
rect 100760 69692 100812 69698
rect 100760 69634 100812 69640
rect 93872 16546 93992 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93964 480 93992 16546
rect 95148 3528 95200 3534
rect 95148 3470 95200 3476
rect 95160 480 95188 3470
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 69634
rect 107660 68400 107712 68406
rect 107660 68342 107712 68348
rect 103520 66972 103572 66978
rect 103520 66914 103572 66920
rect 102140 38004 102192 38010
rect 102140 37946 102192 37952
rect 102152 16574 102180 37946
rect 103532 16574 103560 66914
rect 104900 42152 104952 42158
rect 104900 42094 104952 42100
rect 104912 16574 104940 42094
rect 106924 33788 106976 33794
rect 106924 33730 106976 33736
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 102244 480 102272 16546
rect 103334 10432 103390 10441
rect 103334 10367 103390 10376
rect 103348 480 103376 10367
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 106464 11756 106516 11762
rect 106464 11698 106516 11704
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 11698
rect 106936 3466 106964 33730
rect 107672 16574 107700 68342
rect 110420 65612 110472 65618
rect 110420 65554 110472 65560
rect 109040 53168 109092 53174
rect 109040 53110 109092 53116
rect 107672 16546 108160 16574
rect 106924 3460 106976 3466
rect 106924 3402 106976 3408
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 53110
rect 110432 6914 110460 65554
rect 121460 64252 121512 64258
rect 121460 64194 121512 64200
rect 118700 55888 118752 55894
rect 118700 55830 118752 55836
rect 115940 46232 115992 46238
rect 115940 46174 115992 46180
rect 111800 44872 111852 44878
rect 111800 44814 111852 44820
rect 110512 24200 110564 24206
rect 110512 24142 110564 24148
rect 110524 16574 110552 24142
rect 111812 16574 111840 44814
rect 114560 25628 114612 25634
rect 114560 25570 114612 25576
rect 114572 16574 114600 25570
rect 115952 16574 115980 46174
rect 118712 16574 118740 55830
rect 121472 16574 121500 64194
rect 124218 62792 124274 62801
rect 124218 62727 124274 62736
rect 122840 58744 122892 58750
rect 122840 58686 122892 58692
rect 122852 16574 122880 58686
rect 124232 16574 124260 62727
rect 110524 16546 111656 16574
rect 111812 16546 112392 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 118712 16546 118832 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 110432 6886 110552 6914
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114008 13184 114060 13190
rect 114008 13126 114060 13132
rect 114020 480 114048 13126
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 117320 14544 117372 14550
rect 117320 14486 117372 14492
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 14486
rect 118804 480 118832 16546
rect 120632 15972 120684 15978
rect 120632 15914 120684 15920
rect 119896 3460 119948 3466
rect 119896 3402 119948 3408
rect 119908 480 119936 3402
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 15914
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 75278
rect 188356 3534 188384 90306
rect 191116 75342 191144 232562
rect 191576 178838 191604 249766
rect 191668 183122 191696 262210
rect 191748 258324 191800 258330
rect 191748 258266 191800 258272
rect 191656 183116 191708 183122
rect 191656 183058 191708 183064
rect 191564 178832 191616 178838
rect 191564 178774 191616 178780
rect 191760 175953 191788 258266
rect 192864 242894 192892 270506
rect 192944 269204 192996 269210
rect 192944 269146 192996 269152
rect 192852 242888 192904 242894
rect 192852 242830 192904 242836
rect 191840 240168 191892 240174
rect 191840 240110 191892 240116
rect 191852 238542 191880 240110
rect 192956 239601 192984 269146
rect 193036 253972 193088 253978
rect 193036 253914 193088 253920
rect 192942 239592 192998 239601
rect 192942 239527 192998 239536
rect 191840 238536 191892 238542
rect 191840 238478 191892 238484
rect 193048 182889 193076 253914
rect 193034 182880 193090 182889
rect 193034 182815 193090 182824
rect 191746 175944 191802 175953
rect 191746 175879 191802 175888
rect 191196 117428 191248 117434
rect 191196 117370 191248 117376
rect 191208 93226 191236 117370
rect 193140 96626 193168 295394
rect 193864 294092 193916 294098
rect 193864 294034 193916 294040
rect 193876 185638 193904 294034
rect 195256 289814 195284 698906
rect 200028 510672 200080 510678
rect 200028 510614 200080 510620
rect 198648 315308 198700 315314
rect 198648 315250 198700 315256
rect 198556 301504 198608 301510
rect 198556 301446 198608 301452
rect 197268 298172 197320 298178
rect 197268 298114 197320 298120
rect 196624 294296 196676 294302
rect 196624 294238 196676 294244
rect 195796 292596 195848 292602
rect 195796 292538 195848 292544
rect 195244 289808 195296 289814
rect 195244 289750 195296 289756
rect 195704 260976 195756 260982
rect 195704 260918 195756 260924
rect 194508 248736 194560 248742
rect 194508 248678 194560 248684
rect 194416 247104 194468 247110
rect 194416 247046 194468 247052
rect 193864 185632 193916 185638
rect 193864 185574 193916 185580
rect 194428 177410 194456 247046
rect 194416 177404 194468 177410
rect 194416 177346 194468 177352
rect 194520 176186 194548 248678
rect 195612 244316 195664 244322
rect 195612 244258 195664 244264
rect 195624 177342 195652 244258
rect 195716 204950 195744 260918
rect 195808 239834 195836 292538
rect 196636 284986 196664 294238
rect 197084 294024 197136 294030
rect 197084 293966 197136 293972
rect 196624 284980 196676 284986
rect 196624 284922 196676 284928
rect 195888 276140 195940 276146
rect 195888 276082 195940 276088
rect 195796 239828 195848 239834
rect 195796 239770 195848 239776
rect 195704 204944 195756 204950
rect 195704 204886 195756 204892
rect 195900 185609 195928 276082
rect 196990 272912 197046 272921
rect 196990 272847 197046 272856
rect 197004 225622 197032 272847
rect 197096 239737 197124 293966
rect 197280 284481 197308 298114
rect 197358 291272 197414 291281
rect 197358 291207 197360 291216
rect 197412 291207 197414 291216
rect 197360 291178 197412 291184
rect 197358 290592 197414 290601
rect 197358 290527 197414 290536
rect 197372 289882 197400 290527
rect 197360 289876 197412 289882
rect 197360 289818 197412 289824
rect 197728 289808 197780 289814
rect 197728 289750 197780 289756
rect 197358 289232 197414 289241
rect 197358 289167 197414 289176
rect 197372 288454 197400 289167
rect 197740 288561 197768 289750
rect 197726 288552 197782 288561
rect 197726 288487 197782 288496
rect 197360 288448 197412 288454
rect 197360 288390 197412 288396
rect 197450 287872 197506 287881
rect 197450 287807 197506 287816
rect 197358 287192 197414 287201
rect 197358 287127 197360 287136
rect 197412 287127 197414 287136
rect 197360 287098 197412 287104
rect 197464 287094 197492 287807
rect 197452 287088 197504 287094
rect 197452 287030 197504 287036
rect 197360 287020 197412 287026
rect 197360 286962 197412 286968
rect 197372 286521 197400 286962
rect 197358 286512 197414 286521
rect 197358 286447 197414 286456
rect 198002 285832 198058 285841
rect 198002 285767 198058 285776
rect 197358 285152 197414 285161
rect 197358 285087 197414 285096
rect 197266 284472 197322 284481
rect 197266 284407 197322 284416
rect 197372 284374 197400 285087
rect 197360 284368 197412 284374
rect 197360 284310 197412 284316
rect 197358 280392 197414 280401
rect 197358 280327 197414 280336
rect 197372 280226 197400 280327
rect 197360 280220 197412 280226
rect 197360 280162 197412 280168
rect 197358 279712 197414 279721
rect 197358 279647 197414 279656
rect 197372 278798 197400 279647
rect 197360 278792 197412 278798
rect 197360 278734 197412 278740
rect 197450 278352 197506 278361
rect 197450 278287 197506 278296
rect 197358 277672 197414 277681
rect 197358 277607 197414 277616
rect 197372 277438 197400 277607
rect 197464 277506 197492 278287
rect 197452 277500 197504 277506
rect 197452 277442 197504 277448
rect 197360 277432 197412 277438
rect 197360 277374 197412 277380
rect 197358 276992 197414 277001
rect 197358 276927 197414 276936
rect 197372 276078 197400 276927
rect 197726 276312 197782 276321
rect 197726 276247 197782 276256
rect 197740 276146 197768 276247
rect 197728 276140 197780 276146
rect 197728 276082 197780 276088
rect 197360 276072 197412 276078
rect 197360 276014 197412 276020
rect 197450 275632 197506 275641
rect 197450 275567 197506 275576
rect 197358 274952 197414 274961
rect 197358 274887 197414 274896
rect 197372 274786 197400 274887
rect 197360 274780 197412 274786
rect 197360 274722 197412 274728
rect 197464 274718 197492 275567
rect 197452 274712 197504 274718
rect 197452 274654 197504 274660
rect 197360 274644 197412 274650
rect 197360 274586 197412 274592
rect 197372 274281 197400 274586
rect 197358 274272 197414 274281
rect 197358 274207 197414 274216
rect 197266 272232 197322 272241
rect 197266 272167 197322 272176
rect 197174 248432 197230 248441
rect 197174 248367 197230 248376
rect 197082 239728 197138 239737
rect 197082 239663 197138 239672
rect 196992 225616 197044 225622
rect 196992 225558 197044 225564
rect 195886 185600 195942 185609
rect 195886 185535 195942 185544
rect 197188 177449 197216 248367
rect 197280 184346 197308 272167
rect 197360 271856 197412 271862
rect 197360 271798 197412 271804
rect 197372 270881 197400 271798
rect 197450 271552 197506 271561
rect 197450 271487 197506 271496
rect 197358 270872 197414 270881
rect 197358 270807 197414 270816
rect 197464 270570 197492 271487
rect 197452 270564 197504 270570
rect 197452 270506 197504 270512
rect 197450 270192 197506 270201
rect 197450 270127 197506 270136
rect 197358 269512 197414 269521
rect 197358 269447 197414 269456
rect 197372 269142 197400 269447
rect 197464 269210 197492 270127
rect 197452 269204 197504 269210
rect 197452 269146 197504 269152
rect 197360 269136 197412 269142
rect 197360 269078 197412 269084
rect 197358 268152 197414 268161
rect 197358 268087 197414 268096
rect 197372 267782 197400 268087
rect 197360 267776 197412 267782
rect 197360 267718 197412 267724
rect 197452 267708 197504 267714
rect 197452 267650 197504 267656
rect 197360 267640 197412 267646
rect 197360 267582 197412 267588
rect 197372 266801 197400 267582
rect 197464 267481 197492 267650
rect 197450 267472 197506 267481
rect 197450 267407 197506 267416
rect 197358 266792 197414 266801
rect 197358 266727 197414 266736
rect 197360 266348 197412 266354
rect 197360 266290 197412 266296
rect 197372 265441 197400 266290
rect 197450 266112 197506 266121
rect 197450 266047 197506 266056
rect 197358 265432 197414 265441
rect 197358 265367 197414 265376
rect 197464 264994 197492 266047
rect 197452 264988 197504 264994
rect 197452 264930 197504 264936
rect 197450 264752 197506 264761
rect 197450 264687 197506 264696
rect 197358 264072 197414 264081
rect 197358 264007 197414 264016
rect 197372 263702 197400 264007
rect 197360 263696 197412 263702
rect 197360 263638 197412 263644
rect 197464 263634 197492 264687
rect 197452 263628 197504 263634
rect 197452 263570 197504 263576
rect 197360 263560 197412 263566
rect 197360 263502 197412 263508
rect 197372 263401 197400 263502
rect 197358 263392 197414 263401
rect 197358 263327 197414 263336
rect 197358 262712 197414 262721
rect 197358 262647 197414 262656
rect 197372 262274 197400 262647
rect 197360 262268 197412 262274
rect 197360 262210 197412 262216
rect 197450 262032 197506 262041
rect 197450 261967 197506 261976
rect 197464 260914 197492 261967
rect 197542 261352 197598 261361
rect 197542 261287 197598 261296
rect 197556 260982 197584 261287
rect 197544 260976 197596 260982
rect 197544 260918 197596 260924
rect 197452 260908 197504 260914
rect 197452 260850 197504 260856
rect 197360 260840 197412 260846
rect 197360 260782 197412 260788
rect 197372 260681 197400 260782
rect 197358 260672 197414 260681
rect 197358 260607 197414 260616
rect 197358 259992 197414 260001
rect 197358 259927 197414 259936
rect 197372 259486 197400 259927
rect 197360 259480 197412 259486
rect 197360 259422 197412 259428
rect 197358 259312 197414 259321
rect 197358 259247 197414 259256
rect 197372 258126 197400 259247
rect 197450 258632 197506 258641
rect 197450 258567 197506 258576
rect 197464 258330 197492 258567
rect 197452 258324 197504 258330
rect 197452 258266 197504 258272
rect 197360 258120 197412 258126
rect 197360 258062 197412 258068
rect 197450 257952 197506 257961
rect 197450 257887 197506 257896
rect 197358 257272 197414 257281
rect 197358 257207 197414 257216
rect 197372 256834 197400 257207
rect 197360 256828 197412 256834
rect 197360 256770 197412 256776
rect 197464 256766 197492 257887
rect 197452 256760 197504 256766
rect 197452 256702 197504 256708
rect 197450 255912 197506 255921
rect 197450 255847 197506 255856
rect 197464 255338 197492 255847
rect 197452 255332 197504 255338
rect 197452 255274 197504 255280
rect 197360 255264 197412 255270
rect 197358 255232 197360 255241
rect 197412 255232 197414 255241
rect 197358 255167 197414 255176
rect 197358 254552 197414 254561
rect 197358 254487 197414 254496
rect 197372 253978 197400 254487
rect 197360 253972 197412 253978
rect 197360 253914 197412 253920
rect 197358 253872 197414 253881
rect 197358 253807 197414 253816
rect 197372 252618 197400 253807
rect 197360 252612 197412 252618
rect 197360 252554 197412 252560
rect 197450 252512 197506 252521
rect 197450 252447 197506 252456
rect 197358 251832 197414 251841
rect 197358 251767 197414 251776
rect 197372 251258 197400 251767
rect 197464 251326 197492 252447
rect 198016 252385 198044 285767
rect 198568 283121 198596 301446
rect 198554 283112 198610 283121
rect 198554 283047 198610 283056
rect 198660 281761 198688 315250
rect 198646 281752 198702 281761
rect 198646 281687 198702 281696
rect 198646 281072 198702 281081
rect 198646 281007 198702 281016
rect 198094 273592 198150 273601
rect 198094 273527 198150 273536
rect 198002 252376 198058 252385
rect 198002 252311 198058 252320
rect 197452 251320 197504 251326
rect 197452 251262 197504 251268
rect 197360 251252 197412 251258
rect 197360 251194 197412 251200
rect 198108 250510 198136 273527
rect 198554 251152 198610 251161
rect 198554 251087 198610 251096
rect 198096 250504 198148 250510
rect 197450 250472 197506 250481
rect 198096 250446 198148 250452
rect 197450 250407 197506 250416
rect 197464 249830 197492 250407
rect 197452 249824 197504 249830
rect 197358 249792 197414 249801
rect 197452 249766 197504 249772
rect 197358 249727 197360 249736
rect 197412 249727 197414 249736
rect 197360 249698 197412 249704
rect 197358 249112 197414 249121
rect 197358 249047 197414 249056
rect 197372 248742 197400 249047
rect 197360 248736 197412 248742
rect 197360 248678 197412 248684
rect 197452 248396 197504 248402
rect 197452 248338 197504 248344
rect 197464 247081 197492 248338
rect 197542 247752 197598 247761
rect 197542 247687 197598 247696
rect 197556 247110 197584 247687
rect 197544 247104 197596 247110
rect 197450 247072 197506 247081
rect 197360 247036 197412 247042
rect 197544 247046 197596 247052
rect 197450 247007 197506 247016
rect 197360 246978 197412 246984
rect 197372 245721 197400 246978
rect 197358 245712 197414 245721
rect 197358 245647 197414 245656
rect 197450 244352 197506 244361
rect 197450 244287 197452 244296
rect 197504 244287 197506 244296
rect 197452 244258 197504 244264
rect 197360 244248 197412 244254
rect 197360 244190 197412 244196
rect 197372 243681 197400 244190
rect 197358 243672 197414 243681
rect 197358 243607 197414 243616
rect 197358 242312 197414 242321
rect 197358 242247 197414 242256
rect 197372 241534 197400 242247
rect 197360 241528 197412 241534
rect 197360 241470 197412 241476
rect 198568 206310 198596 251087
rect 198556 206304 198608 206310
rect 198556 206246 198608 206252
rect 198660 193905 198688 281007
rect 200040 279041 200068 510614
rect 201512 312594 201540 702986
rect 218992 700398 219020 703520
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 235184 699718 235212 703520
rect 267660 699718 267688 703520
rect 268384 700392 268436 700398
rect 268384 700334 268436 700340
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 240784 699712 240836 699718
rect 240784 699654 240836 699660
rect 258724 699712 258776 699718
rect 258724 699654 258776 699660
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 237564 694816 237616 694822
rect 237564 694758 237616 694764
rect 215668 693456 215720 693462
rect 215668 693398 215720 693404
rect 206284 404388 206336 404394
rect 206284 404330 206336 404336
rect 204904 351960 204956 351966
rect 204904 351902 204956 351908
rect 201500 312588 201552 312594
rect 201500 312530 201552 312536
rect 203432 300960 203484 300966
rect 203432 300902 203484 300908
rect 202144 299600 202196 299606
rect 202144 299542 202196 299548
rect 201500 295996 201552 296002
rect 201500 295938 201552 295944
rect 200854 295488 200910 295497
rect 200854 295423 200910 295432
rect 200868 292145 200896 295423
rect 201408 292528 201460 292534
rect 201406 292496 201408 292505
rect 201460 292496 201462 292505
rect 201406 292431 201462 292440
rect 201512 292145 201540 295938
rect 202156 292145 202184 299542
rect 202788 298784 202840 298790
rect 202788 298726 202840 298732
rect 202800 292145 202828 298726
rect 203444 292145 203472 300902
rect 204916 295526 204944 351902
rect 206008 303680 206060 303686
rect 206008 303622 206060 303628
rect 204996 300892 205048 300898
rect 204996 300834 205048 300840
rect 204076 295520 204128 295526
rect 204076 295462 204128 295468
rect 204904 295520 204956 295526
rect 204904 295462 204956 295468
rect 204088 292145 204116 295462
rect 204720 294024 204772 294030
rect 204720 293966 204772 293972
rect 204732 292145 204760 293966
rect 205008 292534 205036 300834
rect 205364 292596 205416 292602
rect 205364 292538 205416 292544
rect 204996 292528 205048 292534
rect 204996 292470 205048 292476
rect 205376 292145 205404 292538
rect 206020 292145 206048 303622
rect 206296 301510 206324 404330
rect 213184 357468 213236 357474
rect 213184 357410 213236 357416
rect 208584 307080 208636 307086
rect 208584 307022 208636 307028
rect 206284 301504 206336 301510
rect 206284 301446 206336 301452
rect 207940 301504 207992 301510
rect 207940 301446 207992 301452
rect 206652 298240 206704 298246
rect 206652 298182 206704 298188
rect 206664 292145 206692 298182
rect 207296 292596 207348 292602
rect 207296 292538 207348 292544
rect 207308 292145 207336 292538
rect 207952 292145 207980 301446
rect 208596 292145 208624 307022
rect 211158 296984 211214 296993
rect 211158 296919 211214 296928
rect 210516 296744 210568 296750
rect 210516 296686 210568 296692
rect 209226 293992 209282 294001
rect 209226 293927 209282 293936
rect 209240 292145 209268 293927
rect 210528 292145 210556 296686
rect 211172 292145 211200 296919
rect 213196 296002 213224 357410
rect 215024 320884 215076 320890
rect 215024 320826 215076 320832
rect 213736 296812 213788 296818
rect 213736 296754 213788 296760
rect 213184 295996 213236 296002
rect 213184 295938 213236 295944
rect 213092 295588 213144 295594
rect 213092 295530 213144 295536
rect 211804 294636 211856 294642
rect 211804 294578 211856 294584
rect 211816 292145 211844 294578
rect 212448 292664 212500 292670
rect 212448 292606 212500 292612
rect 212460 292145 212488 292606
rect 213104 292145 213132 295530
rect 213748 292145 213776 296754
rect 214380 295384 214432 295390
rect 214380 295326 214432 295332
rect 214392 292145 214420 295326
rect 215036 292145 215064 320826
rect 215680 292145 215708 693398
rect 222844 670744 222896 670750
rect 222844 670686 222896 670692
rect 218888 302252 218940 302258
rect 218888 302194 218940 302200
rect 216312 298376 216364 298382
rect 216312 298318 216364 298324
rect 216324 292145 216352 298318
rect 216954 298208 217010 298217
rect 216954 298143 217010 298152
rect 216968 292145 216996 298143
rect 218244 294228 218296 294234
rect 218244 294170 218296 294176
rect 217600 292732 217652 292738
rect 217600 292674 217652 292680
rect 217612 292145 217640 292674
rect 218256 292145 218284 294170
rect 218900 292145 218928 302194
rect 220174 299568 220230 299577
rect 219532 299532 219584 299538
rect 220174 299503 220230 299512
rect 219532 299474 219584 299480
rect 219544 292145 219572 299474
rect 220188 292145 220216 299503
rect 222856 299470 222884 670686
rect 232504 563100 232556 563106
rect 232504 563042 232556 563048
rect 226984 418192 227036 418198
rect 226984 418134 227036 418140
rect 224224 345092 224276 345098
rect 224224 345034 224276 345040
rect 224236 304298 224264 345034
rect 225328 309800 225380 309806
rect 225328 309742 225380 309748
rect 224684 304360 224736 304366
rect 224684 304302 224736 304308
rect 224224 304292 224276 304298
rect 224224 304234 224276 304240
rect 221464 299464 221516 299470
rect 221464 299406 221516 299412
rect 222844 299464 222896 299470
rect 222844 299406 222896 299412
rect 220820 292800 220872 292806
rect 220820 292742 220872 292748
rect 220832 292145 220860 292742
rect 221476 292145 221504 299406
rect 223396 298444 223448 298450
rect 223396 298386 223448 298392
rect 222752 294296 222804 294302
rect 222752 294238 222804 294244
rect 222108 294160 222160 294166
rect 222108 294102 222160 294108
rect 222120 292145 222148 294102
rect 222764 292145 222792 294238
rect 223408 292145 223436 298386
rect 224040 295656 224092 295662
rect 224040 295598 224092 295604
rect 224052 292145 224080 295598
rect 224696 292145 224724 304302
rect 225340 292145 225368 309742
rect 226996 307086 227024 418134
rect 232516 309806 232544 563042
rect 234988 318096 235040 318102
rect 234988 318038 235040 318044
rect 232504 309800 232556 309806
rect 232504 309742 232556 309748
rect 226984 307080 227036 307086
rect 226984 307022 227036 307028
rect 233700 301028 233752 301034
rect 233700 300970 233752 300976
rect 231124 298512 231176 298518
rect 231124 298454 231176 298460
rect 227904 298308 227956 298314
rect 227904 298250 227956 298256
rect 226616 295452 226668 295458
rect 226616 295394 226668 295400
rect 225972 294296 226024 294302
rect 225972 294238 226024 294244
rect 225984 292145 226012 294238
rect 226628 292145 226656 295394
rect 227260 294364 227312 294370
rect 227260 294306 227312 294312
rect 227272 292145 227300 294306
rect 227916 292145 227944 298250
rect 228548 295996 228600 296002
rect 228548 295938 228600 295944
rect 228560 292145 228588 295938
rect 229192 295384 229244 295390
rect 229192 295326 229244 295332
rect 229204 292145 229232 295326
rect 229834 294264 229890 294273
rect 229834 294199 229890 294208
rect 229848 292145 229876 294199
rect 231136 292145 231164 298454
rect 232412 296880 232464 296886
rect 232412 296822 232464 296828
rect 231768 294092 231820 294098
rect 231768 294034 231820 294040
rect 231780 292145 231808 294034
rect 232424 292145 232452 296822
rect 233056 295724 233108 295730
rect 233056 295666 233108 295672
rect 233068 292145 233096 295666
rect 233712 292145 233740 300970
rect 234344 294364 234396 294370
rect 234344 294306 234396 294312
rect 234356 292145 234384 294306
rect 235000 292145 235028 318038
rect 236920 302320 236972 302326
rect 236920 302262 236972 302268
rect 236274 293992 236330 294001
rect 236274 293927 236330 293936
rect 235630 292768 235686 292777
rect 235630 292703 235686 292712
rect 235644 292145 235672 292703
rect 236288 292145 236316 293927
rect 236932 292145 236960 302262
rect 237576 292145 237604 694758
rect 238852 309800 238904 309806
rect 238852 309742 238904 309748
rect 238206 296848 238262 296857
rect 238206 296783 238262 296792
rect 238220 292145 238248 296783
rect 238864 292145 238892 309742
rect 239496 299668 239548 299674
rect 239496 299610 239548 299616
rect 239508 292145 239536 299610
rect 240140 296948 240192 296954
rect 240140 296890 240192 296896
rect 240152 294642 240180 296890
rect 240796 294710 240824 699654
rect 249064 656940 249116 656946
rect 249064 656882 249116 656888
rect 245292 316736 245344 316742
rect 245292 316678 245344 316684
rect 241428 295452 241480 295458
rect 241428 295394 241480 295400
rect 240784 294704 240836 294710
rect 240784 294646 240836 294652
rect 240140 294636 240192 294642
rect 240140 294578 240192 294584
rect 240140 294092 240192 294098
rect 240140 294034 240192 294040
rect 240152 292145 240180 294034
rect 241440 292145 241468 295394
rect 243358 295352 243414 295361
rect 243358 295287 243414 295296
rect 242716 292868 242768 292874
rect 242716 292810 242768 292816
rect 242346 292224 242402 292233
rect 242346 292159 242402 292168
rect 242098 292131 242388 292159
rect 242728 292145 242756 292810
rect 243372 292145 243400 295287
rect 244280 294228 244332 294234
rect 244280 294170 244332 294176
rect 244292 293282 244320 294170
rect 244646 294128 244702 294137
rect 244646 294063 244702 294072
rect 244280 293276 244332 293282
rect 244280 293218 244332 293224
rect 244002 292632 244058 292641
rect 244002 292567 244058 292576
rect 244016 292145 244044 292567
rect 244660 292145 244688 294063
rect 245304 292145 245332 316678
rect 246580 302932 246632 302938
rect 246580 302874 246632 302880
rect 245936 294024 245988 294030
rect 245936 293966 245988 293972
rect 245948 292145 245976 293966
rect 246592 292145 246620 302874
rect 249076 302666 249104 656882
rect 253204 579692 253256 579698
rect 253204 579634 253256 579640
rect 251824 501016 251876 501022
rect 251824 500958 251876 500964
rect 249984 312588 250036 312594
rect 249984 312530 250036 312536
rect 249892 304292 249944 304298
rect 249892 304234 249944 304240
rect 249064 302660 249116 302666
rect 249064 302602 249116 302608
rect 247868 297016 247920 297022
rect 247868 296958 247920 296964
rect 247224 295520 247276 295526
rect 247224 295462 247276 295468
rect 247236 292145 247264 295462
rect 247880 292145 247908 296958
rect 248510 292904 248566 292913
rect 248510 292839 248566 292848
rect 248524 292145 248552 292839
rect 249154 292360 249210 292369
rect 249154 292295 249210 292304
rect 249168 292145 249196 292295
rect 210240 292120 210292 292126
rect 209906 292068 210240 292074
rect 241152 292120 241204 292126
rect 209906 292062 210292 292068
rect 240818 292068 241152 292074
rect 249904 292074 249932 304234
rect 240818 292062 241204 292068
rect 209906 292046 210280 292062
rect 240818 292046 241192 292062
rect 249826 292046 249932 292074
rect 200118 291544 200174 291553
rect 200174 291502 200238 291530
rect 200118 291479 200174 291488
rect 249996 287609 250024 312530
rect 251272 305040 251324 305046
rect 251272 304982 251324 304988
rect 251180 300144 251232 300150
rect 251180 300086 251232 300092
rect 250536 294092 250588 294098
rect 250536 294034 250588 294040
rect 250444 294024 250496 294030
rect 250444 293966 250496 293972
rect 250168 292800 250220 292806
rect 250168 292742 250220 292748
rect 249982 287600 250038 287609
rect 249982 287535 250038 287544
rect 200026 279032 200082 279041
rect 200026 278967 200082 278976
rect 249982 269784 250038 269793
rect 249982 269719 250038 269728
rect 200026 268832 200082 268841
rect 200026 268767 200082 268776
rect 199934 256592 199990 256601
rect 199934 256527 199990 256536
rect 199842 253192 199898 253201
rect 199842 253127 199898 253136
rect 199750 245032 199806 245041
rect 199750 244967 199806 244976
rect 198740 242888 198792 242894
rect 198740 242830 198792 242836
rect 198752 239426 198780 242830
rect 199764 239465 199792 244967
rect 199750 239456 199806 239465
rect 198740 239420 198792 239426
rect 199750 239391 199806 239400
rect 198740 239362 198792 239368
rect 199856 236706 199884 253127
rect 199844 236700 199896 236706
rect 199844 236642 199896 236648
rect 199948 222902 199976 256527
rect 200040 224262 200068 268767
rect 200224 237454 200252 240244
rect 200762 240136 200818 240145
rect 200762 240071 200818 240080
rect 200776 239970 200804 240071
rect 200764 239964 200816 239970
rect 200764 239906 200816 239912
rect 200212 237448 200264 237454
rect 200212 237390 200264 237396
rect 200868 231130 200896 240219
rect 200856 231124 200908 231130
rect 200856 231066 200908 231072
rect 200028 224256 200080 224262
rect 200028 224198 200080 224204
rect 199936 222896 199988 222902
rect 199936 222838 199988 222844
rect 198646 193896 198702 193905
rect 198646 193831 198702 193840
rect 201512 185774 201540 240219
rect 202156 196654 202184 240219
rect 202800 237862 202828 240219
rect 202788 237856 202840 237862
rect 202788 237798 202840 237804
rect 202144 196648 202196 196654
rect 202144 196590 202196 196596
rect 201500 185768 201552 185774
rect 201500 185710 201552 185716
rect 197268 184340 197320 184346
rect 197268 184282 197320 184288
rect 203444 182850 203472 240219
rect 203432 182844 203484 182850
rect 203432 182786 203484 182792
rect 204088 178702 204116 240219
rect 204732 191049 204760 240219
rect 204718 191040 204774 191049
rect 204718 190975 204774 190984
rect 205376 186969 205404 240219
rect 206028 240106 206056 240219
rect 206016 240100 206068 240106
rect 206016 240042 206068 240048
rect 206376 239964 206428 239970
rect 206376 239906 206428 239912
rect 205548 237856 205600 237862
rect 205548 237798 205600 237804
rect 205560 235958 205588 237798
rect 206284 237448 206336 237454
rect 206284 237390 206336 237396
rect 205548 235952 205600 235958
rect 205548 235894 205600 235900
rect 205362 186960 205418 186969
rect 205362 186895 205418 186904
rect 204904 182232 204956 182238
rect 204904 182174 204956 182180
rect 204076 178696 204128 178702
rect 204076 178638 204128 178644
rect 197174 177440 197230 177449
rect 197174 177375 197230 177384
rect 195612 177336 195664 177342
rect 195612 177278 195664 177284
rect 198004 176792 198056 176798
rect 198004 176734 198056 176740
rect 194508 176180 194560 176186
rect 194508 176122 194560 176128
rect 198016 171018 198044 176734
rect 204916 173806 204944 182174
rect 206296 178770 206324 237390
rect 206388 181393 206416 239906
rect 206664 232558 206692 240219
rect 206652 232552 206704 232558
rect 206652 232494 206704 232500
rect 207308 197985 207336 240219
rect 207294 197976 207350 197985
rect 207294 197911 207350 197920
rect 207952 184249 207980 240219
rect 207938 184240 207994 184249
rect 207938 184175 207994 184184
rect 206374 181384 206430 181393
rect 206374 181319 206430 181328
rect 208596 178906 208624 240219
rect 209044 183592 209096 183598
rect 209044 183534 209096 183540
rect 208584 178900 208636 178906
rect 208584 178842 208636 178848
rect 206284 178764 206336 178770
rect 206284 178706 206336 178712
rect 204904 173800 204956 173806
rect 204904 173742 204956 173748
rect 198004 171012 198056 171018
rect 198004 170954 198056 170960
rect 209056 157350 209084 183534
rect 209240 180169 209268 240219
rect 209226 180160 209282 180169
rect 209226 180095 209282 180104
rect 209884 180033 209912 240219
rect 210528 188426 210556 240219
rect 211172 211818 211200 240219
rect 211816 238746 211844 240219
rect 212460 239902 212488 240219
rect 212448 239896 212500 239902
rect 212448 239838 212500 239844
rect 211804 238740 211856 238746
rect 211804 238682 211856 238688
rect 213104 228313 213132 240219
rect 213748 228410 213776 240219
rect 213736 228404 213788 228410
rect 213736 228346 213788 228352
rect 213090 228304 213146 228313
rect 213090 228239 213146 228248
rect 211160 211812 211212 211818
rect 211160 211754 211212 211760
rect 210516 188420 210568 188426
rect 210516 188362 210568 188368
rect 214392 182918 214420 240219
rect 215036 200802 215064 240219
rect 215024 200796 215076 200802
rect 215024 200738 215076 200744
rect 214380 182912 214432 182918
rect 214380 182854 214432 182860
rect 215680 181490 215708 240219
rect 215944 239420 215996 239426
rect 215944 239362 215996 239368
rect 215668 181484 215720 181490
rect 215668 181426 215720 181432
rect 213276 180872 213328 180878
rect 213276 180814 213328 180820
rect 209870 180024 209926 180033
rect 209870 179959 209926 179968
rect 211804 179444 211856 179450
rect 211804 179386 211856 179392
rect 211816 164150 211844 179386
rect 213184 178084 213236 178090
rect 213184 178026 213236 178032
rect 211896 175976 211948 175982
rect 211896 175918 211948 175924
rect 211908 165510 211936 175918
rect 211896 165504 211948 165510
rect 211896 165446 211948 165452
rect 211804 164144 211856 164150
rect 211804 164086 211856 164092
rect 213196 162081 213224 178026
rect 213288 166977 213316 180814
rect 214196 179512 214248 179518
rect 214196 179454 214248 179460
rect 214012 178152 214064 178158
rect 214012 178094 214064 178100
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175817 213960 176598
rect 213918 175808 213974 175817
rect 213918 175743 213974 175752
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175137 213960 175170
rect 213918 175128 213974 175137
rect 213918 175063 213974 175072
rect 214024 174729 214052 178094
rect 214104 177064 214156 177070
rect 214104 177006 214156 177012
rect 214010 174720 214066 174729
rect 214010 174655 214066 174664
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173777 213960 173810
rect 214012 173800 214064 173806
rect 213918 173768 213974 173777
rect 214012 173742 214064 173748
rect 213918 173703 213974 173712
rect 214024 173369 214052 173742
rect 214010 173360 214066 173369
rect 214010 173295 214066 173304
rect 214116 172009 214144 177006
rect 214208 172417 214236 179454
rect 214564 176928 214616 176934
rect 214564 176870 214616 176876
rect 214194 172408 214250 172417
rect 214194 172343 214250 172352
rect 214102 172000 214158 172009
rect 214102 171935 214158 171944
rect 213920 171080 213972 171086
rect 213920 171022 213972 171028
rect 213932 170785 213960 171022
rect 214012 171012 214064 171018
rect 214012 170954 214064 170960
rect 213918 170776 213974 170785
rect 213918 170711 213974 170720
rect 214024 170649 214052 170954
rect 214010 170640 214066 170649
rect 214010 170575 214066 170584
rect 213920 169720 213972 169726
rect 213920 169662 213972 169668
rect 213932 169425 213960 169662
rect 214012 169652 214064 169658
rect 214012 169594 214064 169600
rect 213918 169416 213974 169425
rect 213918 169351 213974 169360
rect 214024 169289 214052 169594
rect 214010 169280 214066 169289
rect 214010 169215 214066 169224
rect 213920 168360 213972 168366
rect 213920 168302 213972 168308
rect 213932 168065 213960 168302
rect 214012 168292 214064 168298
rect 214012 168234 214064 168240
rect 213918 168056 213974 168065
rect 213918 167991 213974 168000
rect 214024 167929 214052 168234
rect 214010 167920 214066 167929
rect 214010 167855 214066 167864
rect 213274 166968 213330 166977
rect 213274 166903 213330 166912
rect 214012 166932 214064 166938
rect 214012 166874 214064 166880
rect 213920 166864 213972 166870
rect 213920 166806 213972 166812
rect 213932 166705 213960 166806
rect 213918 166696 213974 166705
rect 213918 166631 213974 166640
rect 214024 166161 214052 166874
rect 214010 166152 214066 166161
rect 214010 166087 214066 166096
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 164801 213960 165514
rect 213918 164792 213974 164801
rect 213918 164727 213974 164736
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163441 213960 164154
rect 214472 164144 214524 164150
rect 214470 164112 214472 164121
rect 214524 164112 214526 164121
rect 214470 164047 214526 164056
rect 213918 163432 213974 163441
rect 213918 163367 213974 163376
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162625 213960 162794
rect 213918 162616 213974 162625
rect 213918 162551 213974 162560
rect 213182 162072 213238 162081
rect 213182 162007 213238 162016
rect 213920 161424 213972 161430
rect 213918 161392 213920 161401
rect 213972 161392 213974 161401
rect 213918 161327 213974 161336
rect 214104 160744 214156 160750
rect 214104 160686 214156 160692
rect 213920 160064 213972 160070
rect 213918 160032 213920 160041
rect 213972 160032 213974 160041
rect 213918 159967 213974 159976
rect 214012 159996 214064 160002
rect 214012 159938 214064 159944
rect 214024 159497 214052 159938
rect 214010 159488 214066 159497
rect 214010 159423 214066 159432
rect 213920 158704 213972 158710
rect 213918 158672 213920 158681
rect 213972 158672 213974 158681
rect 213918 158607 213974 158616
rect 214116 158137 214144 160686
rect 214102 158128 214158 158137
rect 214102 158063 214158 158072
rect 209044 157344 209096 157350
rect 209044 157286 209096 157292
rect 213920 157344 213972 157350
rect 213920 157286 213972 157292
rect 213932 156913 213960 157286
rect 213918 156904 213974 156913
rect 213918 156839 213974 156848
rect 213920 155916 213972 155922
rect 213920 155858 213972 155864
rect 213932 155553 213960 155858
rect 213918 155544 213974 155553
rect 213918 155479 213974 155488
rect 214010 153912 214066 153921
rect 214010 153847 214066 153856
rect 213918 153368 213974 153377
rect 213918 153303 213920 153312
rect 213972 153303 213974 153312
rect 213920 153274 213972 153280
rect 214024 153270 214052 153847
rect 214012 153264 214064 153270
rect 214012 153206 214064 153212
rect 214010 152688 214066 152697
rect 214010 152623 214066 152632
rect 213918 152008 213974 152017
rect 213918 151943 213974 151952
rect 213932 151910 213960 151943
rect 196624 151904 196676 151910
rect 196624 151846 196676 151852
rect 213920 151904 213972 151910
rect 213920 151846 213972 151852
rect 193128 96620 193180 96626
rect 193128 96562 193180 96568
rect 191196 93220 191248 93226
rect 191196 93162 191248 93168
rect 196636 85270 196664 151846
rect 214024 151842 214052 152623
rect 214012 151836 214064 151842
rect 214012 151778 214064 151784
rect 214010 150784 214066 150793
rect 214010 150719 214066 150728
rect 213918 150648 213974 150657
rect 213918 150583 213974 150592
rect 213932 150550 213960 150583
rect 198096 150544 198148 150550
rect 198096 150486 198148 150492
rect 213920 150544 213972 150550
rect 213920 150486 213972 150492
rect 198108 122126 198136 150486
rect 214024 150482 214052 150719
rect 214012 150476 214064 150482
rect 214012 150418 214064 150424
rect 213920 150408 213972 150414
rect 213920 150350 213972 150356
rect 213932 149569 213960 150350
rect 214576 150249 214604 176870
rect 214656 174548 214708 174554
rect 214656 174490 214708 174496
rect 214668 171134 214696 174490
rect 214668 171106 214788 171134
rect 214656 165504 214708 165510
rect 214654 165472 214656 165481
rect 214708 165472 214710 165481
rect 214654 165407 214710 165416
rect 214562 150240 214618 150249
rect 214562 150175 214618 150184
rect 213918 149560 213974 149569
rect 213918 149495 213974 149504
rect 214760 148889 214788 171106
rect 215022 151872 215078 151881
rect 215022 151807 215078 151816
rect 214746 148880 214802 148889
rect 214746 148815 214802 148824
rect 213918 148064 213974 148073
rect 213918 147999 213974 148008
rect 213932 147694 213960 147999
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 213918 146704 213974 146713
rect 213918 146639 213974 146648
rect 213932 146334 213960 146639
rect 214562 146432 214618 146441
rect 214562 146367 214618 146376
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 213918 145344 213974 145353
rect 213918 145279 213974 145288
rect 213932 144974 213960 145279
rect 213920 144968 213972 144974
rect 213920 144910 213972 144916
rect 214010 143984 214066 143993
rect 214010 143919 214066 143928
rect 214024 143682 214052 143919
rect 214012 143676 214064 143682
rect 214012 143618 214064 143624
rect 213920 143608 213972 143614
rect 213918 143576 213920 143585
rect 213972 143576 213974 143585
rect 213918 143511 213974 143520
rect 213918 142760 213974 142769
rect 213918 142695 213974 142704
rect 213932 142186 213960 142695
rect 213920 142180 213972 142186
rect 213920 142122 213972 142128
rect 214010 141400 214066 141409
rect 214010 141335 214066 141344
rect 213918 140992 213974 141001
rect 213918 140927 213974 140936
rect 213932 140894 213960 140927
rect 213920 140888 213972 140894
rect 213920 140830 213972 140836
rect 214024 140826 214052 141335
rect 214012 140820 214064 140826
rect 214012 140762 214064 140768
rect 213918 139496 213974 139505
rect 210424 139460 210476 139466
rect 213918 139431 213920 139440
rect 210424 139402 210476 139408
rect 213972 139431 213974 139440
rect 213920 139402 213972 139408
rect 202144 138100 202196 138106
rect 202144 138042 202196 138048
rect 199384 124296 199436 124302
rect 199384 124238 199436 124244
rect 198096 122120 198148 122126
rect 198096 122062 198148 122068
rect 198004 121508 198056 121514
rect 198004 121450 198056 121456
rect 196716 110560 196768 110566
rect 196716 110502 196768 110508
rect 196728 92410 196756 110502
rect 196716 92404 196768 92410
rect 196716 92346 196768 92352
rect 198016 89554 198044 121450
rect 198004 89548 198056 89554
rect 198004 89490 198056 89496
rect 196624 85264 196676 85270
rect 196624 85206 196676 85212
rect 199396 79898 199424 124238
rect 202156 92342 202184 138042
rect 206376 136672 206428 136678
rect 206376 136614 206428 136620
rect 204904 133952 204956 133958
rect 204904 133894 204956 133900
rect 202236 107704 202288 107710
rect 202236 107646 202288 107652
rect 202144 92336 202196 92342
rect 202144 92278 202196 92284
rect 202248 81394 202276 107646
rect 202236 81388 202288 81394
rect 202236 81330 202288 81336
rect 199384 79892 199436 79898
rect 199384 79834 199436 79840
rect 204916 78606 204944 133894
rect 206284 131232 206336 131238
rect 206284 131174 206336 131180
rect 204996 104984 205048 104990
rect 204996 104926 205048 104932
rect 205008 94897 205036 104926
rect 205088 103556 205140 103562
rect 205088 103498 205140 103504
rect 205100 95062 205128 103498
rect 205088 95056 205140 95062
rect 205088 94998 205140 95004
rect 204994 94888 205050 94897
rect 204994 94823 205050 94832
rect 204904 78600 204956 78606
rect 204904 78542 204956 78548
rect 191104 75336 191156 75342
rect 191104 75278 191156 75284
rect 206296 74526 206324 131174
rect 206388 79966 206416 136614
rect 209136 114640 209188 114646
rect 209136 114582 209188 114588
rect 209044 107772 209096 107778
rect 209044 107714 209096 107720
rect 207756 100836 207808 100842
rect 207756 100778 207808 100784
rect 207664 96688 207716 96694
rect 207664 96630 207716 96636
rect 207676 85542 207704 96630
rect 207768 89690 207796 100778
rect 207756 89684 207808 89690
rect 207756 89626 207808 89632
rect 207664 85536 207716 85542
rect 207664 85478 207716 85484
rect 206376 79960 206428 79966
rect 206376 79902 206428 79908
rect 209056 78674 209084 107714
rect 209148 93158 209176 114582
rect 209228 98116 209280 98122
rect 209228 98058 209280 98064
rect 209136 93152 209188 93158
rect 209136 93094 209188 93100
rect 209240 86902 209268 98058
rect 209228 86896 209280 86902
rect 209228 86838 209280 86844
rect 210436 84114 210464 139402
rect 214010 138816 214066 138825
rect 214010 138751 214066 138760
rect 213918 138136 213974 138145
rect 213918 138071 213920 138080
rect 213972 138071 213974 138080
rect 213920 138042 213972 138048
rect 214024 138038 214052 138751
rect 214012 138032 214064 138038
rect 214012 137974 214064 137980
rect 213918 137456 213974 137465
rect 213918 137391 213974 137400
rect 213932 136678 213960 137391
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 213182 136096 213238 136105
rect 213182 136031 213238 136040
rect 211804 121576 211856 121582
rect 211804 121518 211856 121524
rect 210516 106412 210568 106418
rect 210516 106354 210568 106360
rect 210424 84108 210476 84114
rect 210424 84050 210476 84056
rect 210528 80034 210556 106354
rect 211816 81326 211844 121518
rect 211896 111920 211948 111926
rect 211896 111862 211948 111868
rect 211908 86970 211936 111862
rect 211896 86964 211948 86970
rect 211896 86906 211948 86912
rect 213196 85474 213224 136031
rect 213918 134056 213974 134065
rect 213918 133991 213974 134000
rect 213932 133958 213960 133991
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 214010 132832 214066 132841
rect 214010 132767 214066 132776
rect 213920 132592 213972 132598
rect 213918 132560 213920 132569
rect 213972 132560 213974 132569
rect 214024 132530 214052 132767
rect 213918 132495 213974 132504
rect 214012 132524 214064 132530
rect 214012 132466 214064 132472
rect 214010 131472 214066 131481
rect 214010 131407 214066 131416
rect 213920 131232 213972 131238
rect 213918 131200 213920 131209
rect 213972 131200 213974 131209
rect 214024 131170 214052 131407
rect 213918 131135 213974 131144
rect 214012 131164 214064 131170
rect 214012 131106 214064 131112
rect 214010 130112 214066 130121
rect 214010 130047 214066 130056
rect 214024 129878 214052 130047
rect 214012 129872 214064 129878
rect 213918 129840 213974 129849
rect 214012 129814 214064 129820
rect 213918 129775 213920 129784
rect 213972 129775 213974 129784
rect 213920 129746 213972 129752
rect 213918 128480 213974 128489
rect 213918 128415 213974 128424
rect 213932 128382 213960 128415
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 213918 127120 213974 127129
rect 213918 127055 213974 127064
rect 213932 127022 213960 127055
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 214010 126168 214066 126177
rect 214010 126103 214066 126112
rect 213918 125760 213974 125769
rect 214024 125730 214052 126103
rect 213918 125695 213974 125704
rect 214012 125724 214064 125730
rect 213932 125662 213960 125695
rect 214012 125666 214064 125672
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214010 124808 214066 124817
rect 214010 124743 214066 124752
rect 213918 124400 213974 124409
rect 213918 124335 213974 124344
rect 213932 124302 213960 124335
rect 213920 124296 213972 124302
rect 213920 124238 213972 124244
rect 214024 124234 214052 124743
rect 214012 124228 214064 124234
rect 214012 124170 214064 124176
rect 214010 123584 214066 123593
rect 214010 123519 214066 123528
rect 213918 123176 213974 123185
rect 213918 123111 213974 123120
rect 213932 122942 213960 123111
rect 213920 122936 213972 122942
rect 213920 122878 213972 122884
rect 214024 122874 214052 123519
rect 214012 122868 214064 122874
rect 214012 122810 214064 122816
rect 213918 122224 213974 122233
rect 213918 122159 213974 122168
rect 213932 121514 213960 122159
rect 214470 121680 214526 121689
rect 214470 121615 214526 121624
rect 214484 121582 214512 121615
rect 214472 121576 214524 121582
rect 214472 121518 214524 121524
rect 213920 121508 213972 121514
rect 213920 121450 213972 121456
rect 214010 120864 214066 120873
rect 214010 120799 214066 120808
rect 213918 120456 213974 120465
rect 213918 120391 213974 120400
rect 213932 120222 213960 120391
rect 213920 120216 213972 120222
rect 213920 120158 213972 120164
rect 214024 120154 214052 120799
rect 214012 120148 214064 120154
rect 214012 120090 214064 120096
rect 214010 119640 214066 119649
rect 214010 119575 214066 119584
rect 213274 119096 213330 119105
rect 213274 119031 213330 119040
rect 213184 85468 213236 85474
rect 213184 85410 213236 85416
rect 213288 82754 213316 119031
rect 213918 118960 213974 118969
rect 213918 118895 213974 118904
rect 213932 118794 213960 118895
rect 214024 118862 214052 119575
rect 214012 118856 214064 118862
rect 214012 118798 214064 118804
rect 213920 118788 213972 118794
rect 213920 118730 213972 118736
rect 214010 117600 214066 117609
rect 214010 117535 214066 117544
rect 214024 117434 214052 117535
rect 214012 117428 214064 117434
rect 214012 117370 214064 117376
rect 213920 117360 213972 117366
rect 213918 117328 213920 117337
rect 213972 117328 213974 117337
rect 213918 117263 213974 117272
rect 213918 116240 213974 116249
rect 213918 116175 213974 116184
rect 213932 116006 213960 116175
rect 213920 116000 213972 116006
rect 213366 115968 213422 115977
rect 213920 115942 213972 115948
rect 213366 115903 213422 115912
rect 213380 84182 213408 115903
rect 214010 115016 214066 115025
rect 214010 114951 214066 114960
rect 214024 114646 214052 114951
rect 214012 114640 214064 114646
rect 213918 114608 213974 114617
rect 214012 114582 214064 114588
rect 213918 114543 213920 114552
rect 213972 114543 213974 114552
rect 213920 114514 213972 114520
rect 214010 113656 214066 113665
rect 214010 113591 214066 113600
rect 213920 113280 213972 113286
rect 213918 113248 213920 113257
rect 213972 113248 213974 113257
rect 214024 113218 214052 113591
rect 213918 113183 213974 113192
rect 214012 113212 214064 113218
rect 214012 113154 214064 113160
rect 214010 112296 214066 112305
rect 214010 112231 214066 112240
rect 214024 111926 214052 112231
rect 214012 111920 214064 111926
rect 213918 111888 213974 111897
rect 214012 111862 214064 111868
rect 213918 111823 213920 111832
rect 213972 111823 213974 111832
rect 213920 111794 213972 111800
rect 214010 110936 214066 110945
rect 214010 110871 214066 110880
rect 213920 110560 213972 110566
rect 213918 110528 213920 110537
rect 213972 110528 213974 110537
rect 214024 110498 214052 110871
rect 213918 110463 213974 110472
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 214010 109712 214066 109721
rect 214010 109647 214066 109656
rect 213918 109168 213974 109177
rect 213918 109103 213920 109112
rect 213972 109103 213974 109112
rect 213920 109074 213972 109080
rect 214024 109070 214052 109647
rect 214012 109064 214064 109070
rect 214012 109006 214064 109012
rect 214010 108352 214066 108361
rect 214010 108287 214066 108296
rect 213918 107944 213974 107953
rect 213918 107879 213974 107888
rect 213932 107710 213960 107879
rect 214024 107778 214052 108287
rect 214012 107772 214064 107778
rect 214012 107714 214064 107720
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 214010 106992 214066 107001
rect 214010 106927 214066 106936
rect 213918 106584 213974 106593
rect 213918 106519 213974 106528
rect 213932 106350 213960 106519
rect 214024 106418 214052 106927
rect 214012 106412 214064 106418
rect 214012 106354 214064 106360
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 214010 105768 214066 105777
rect 214010 105703 214066 105712
rect 213918 105360 213974 105369
rect 213918 105295 213974 105304
rect 213458 105224 213514 105233
rect 213458 105159 213514 105168
rect 213472 93809 213500 105159
rect 213932 104990 213960 105295
rect 214024 105058 214052 105703
rect 214012 105052 214064 105058
rect 214012 104994 214064 105000
rect 213920 104984 213972 104990
rect 213920 104926 213972 104932
rect 213918 103728 213974 103737
rect 213918 103663 213974 103672
rect 213932 103562 213960 103663
rect 213920 103556 213972 103562
rect 213920 103498 213972 103504
rect 214576 101454 214604 146367
rect 215036 142154 215064 151807
rect 214852 142126 215064 142154
rect 214746 135552 214802 135561
rect 214746 135487 214802 135496
rect 214654 134192 214710 134201
rect 214654 134127 214710 134136
rect 214564 101448 214616 101454
rect 214564 101390 214616 101396
rect 214010 101280 214066 101289
rect 214010 101215 214066 101224
rect 213918 101144 213974 101153
rect 213918 101079 213974 101088
rect 213932 100774 213960 101079
rect 214024 100842 214052 101215
rect 214012 100836 214064 100842
rect 214012 100778 214064 100784
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 213918 99784 213974 99793
rect 213918 99719 213974 99728
rect 213932 99414 213960 99719
rect 214102 99512 214158 99521
rect 214102 99447 214158 99456
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214010 98424 214066 98433
rect 214010 98359 214066 98368
rect 213920 98116 213972 98122
rect 213920 98058 213972 98064
rect 213932 98025 213960 98058
rect 214024 98054 214052 98359
rect 214012 98048 214064 98054
rect 213918 98016 213974 98025
rect 214012 97990 214064 97996
rect 213918 97951 213974 97960
rect 213918 97064 213974 97073
rect 213918 96999 213974 97008
rect 213932 96694 213960 96999
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 214116 95849 214144 99447
rect 214102 95840 214158 95849
rect 214102 95775 214158 95784
rect 214562 95840 214618 95849
rect 214562 95775 214618 95784
rect 213458 93800 213514 93809
rect 213458 93735 213514 93744
rect 213368 84176 213420 84182
rect 213368 84118 213420 84124
rect 214576 82822 214604 95775
rect 214668 94518 214696 134127
rect 214760 108497 214788 135487
rect 214852 134570 214880 142126
rect 214840 134564 214892 134570
rect 214840 134506 214892 134512
rect 214746 108488 214802 108497
rect 214746 108423 214802 108432
rect 214746 102504 214802 102513
rect 214746 102439 214802 102448
rect 214656 94512 214708 94518
rect 214656 94454 214708 94460
rect 214564 82816 214616 82822
rect 214564 82758 214616 82764
rect 213276 82748 213328 82754
rect 213276 82690 213328 82696
rect 211804 81320 211856 81326
rect 211804 81262 211856 81268
rect 210516 80028 210568 80034
rect 210516 79970 210568 79976
rect 209044 78668 209096 78674
rect 209044 78610 209096 78616
rect 214760 77246 214788 102439
rect 214838 96656 214894 96665
rect 214838 96591 214894 96600
rect 214852 88233 214880 96591
rect 215956 95130 215984 239362
rect 215944 95124 215996 95130
rect 215944 95066 215996 95072
rect 216324 92614 216352 240219
rect 216968 238678 216996 240219
rect 216956 238672 217008 238678
rect 216956 238614 217008 238620
rect 217612 191146 217640 240219
rect 217600 191140 217652 191146
rect 217600 191082 217652 191088
rect 218256 178974 218284 240219
rect 218900 238066 218928 240219
rect 219544 238513 219572 240219
rect 219530 238504 219586 238513
rect 219530 238439 219586 238448
rect 218888 238060 218940 238066
rect 218888 238002 218940 238008
rect 220188 183190 220216 240219
rect 220176 183184 220228 183190
rect 220176 183126 220228 183132
rect 218244 178968 218296 178974
rect 218244 178910 218296 178916
rect 220832 177478 220860 240219
rect 221476 238678 221504 240219
rect 222120 238746 222148 240219
rect 222108 238740 222160 238746
rect 222108 238682 222160 238688
rect 221464 238672 221516 238678
rect 221464 238614 221516 238620
rect 222764 177546 222792 240219
rect 223408 185638 223436 240219
rect 224052 191214 224080 240219
rect 224040 191208 224092 191214
rect 224040 191150 224092 191156
rect 223396 185632 223448 185638
rect 223396 185574 223448 185580
rect 224696 180130 224724 240219
rect 225340 184210 225368 240219
rect 225984 238649 226012 240219
rect 225970 238640 226026 238649
rect 225970 238575 226026 238584
rect 225328 184204 225380 184210
rect 225328 184146 225380 184152
rect 226628 180266 226656 240219
rect 226616 180260 226668 180266
rect 226616 180202 226668 180208
rect 224684 180124 224736 180130
rect 224684 180066 224736 180072
rect 227272 178022 227300 240219
rect 227916 184278 227944 240219
rect 228560 238610 228588 240219
rect 228548 238604 228600 238610
rect 228548 238546 228600 238552
rect 229204 238474 229232 240219
rect 229192 238468 229244 238474
rect 229192 238410 229244 238416
rect 229848 202162 229876 240219
rect 230492 225758 230520 240219
rect 231136 233238 231164 240219
rect 231124 233232 231176 233238
rect 231124 233174 231176 233180
rect 230480 225752 230532 225758
rect 230480 225694 230532 225700
rect 230480 225616 230532 225622
rect 230480 225558 230532 225564
rect 229836 202156 229888 202162
rect 229836 202098 229888 202104
rect 227904 184272 227956 184278
rect 227904 184214 227956 184220
rect 227628 180464 227680 180470
rect 227628 180406 227680 180412
rect 227260 178016 227312 178022
rect 227260 177958 227312 177964
rect 222752 177540 222804 177546
rect 222752 177482 222804 177488
rect 220820 177472 220872 177478
rect 220820 177414 220872 177420
rect 227640 175817 227668 180406
rect 229100 178968 229152 178974
rect 229100 178910 229152 178916
rect 227626 175808 227682 175817
rect 227626 175743 227682 175752
rect 229112 154329 229140 178910
rect 229192 178016 229244 178022
rect 229192 177958 229244 177964
rect 229204 169017 229232 177958
rect 229190 169008 229246 169017
rect 229190 168943 229246 168952
rect 229098 154320 229154 154329
rect 229098 154255 229154 154264
rect 230492 147801 230520 225558
rect 230572 224256 230624 224262
rect 230572 224198 230624 224204
rect 230584 161474 230612 224198
rect 231780 223582 231808 240219
rect 231860 225752 231912 225758
rect 231860 225694 231912 225700
rect 231768 223576 231820 223582
rect 231768 223518 231820 223524
rect 230664 222896 230716 222902
rect 230664 222838 230716 222844
rect 230676 166274 230704 222838
rect 230756 184340 230808 184346
rect 230756 184282 230808 184288
rect 230768 171134 230796 184282
rect 231766 175264 231822 175273
rect 231124 175228 231176 175234
rect 231766 175199 231822 175208
rect 231124 175170 231176 175176
rect 231136 174729 231164 175170
rect 231780 175166 231808 175199
rect 231768 175160 231820 175166
rect 231768 175102 231820 175108
rect 231122 174720 231178 174729
rect 231122 174655 231178 174664
rect 231216 173868 231268 173874
rect 231216 173810 231268 173816
rect 231228 173369 231256 173810
rect 231768 173800 231820 173806
rect 231674 173768 231730 173777
rect 231768 173742 231820 173748
rect 231674 173703 231676 173712
rect 231728 173703 231730 173712
rect 231676 173674 231728 173680
rect 231214 173360 231270 173369
rect 231214 173295 231270 173304
rect 231780 172825 231808 173742
rect 231766 172816 231822 172825
rect 231766 172751 231822 172760
rect 231768 172508 231820 172514
rect 231768 172450 231820 172456
rect 231676 172440 231728 172446
rect 231780 172417 231808 172450
rect 231676 172382 231728 172388
rect 231766 172408 231822 172417
rect 231688 171873 231716 172382
rect 231766 172343 231822 172352
rect 231674 171864 231730 171873
rect 231674 171799 231730 171808
rect 231676 171760 231728 171766
rect 231676 171702 231728 171708
rect 231688 171465 231716 171702
rect 231674 171456 231730 171465
rect 231674 171391 231730 171400
rect 230768 171106 230980 171134
rect 230676 166246 230796 166274
rect 230664 164620 230716 164626
rect 230664 164562 230716 164568
rect 230676 164393 230704 164562
rect 230662 164384 230718 164393
rect 230662 164319 230718 164328
rect 230584 161446 230704 161474
rect 230676 158681 230704 161446
rect 230662 158672 230718 158681
rect 230662 158607 230718 158616
rect 230768 157729 230796 166246
rect 230754 157720 230810 157729
rect 230754 157655 230810 157664
rect 230952 156233 230980 171106
rect 231768 171080 231820 171086
rect 231768 171022 231820 171028
rect 231780 170921 231808 171022
rect 231766 170912 231822 170921
rect 231766 170847 231822 170856
rect 231308 170604 231360 170610
rect 231308 170546 231360 170552
rect 231320 169969 231348 170546
rect 231768 170536 231820 170542
rect 231766 170504 231768 170513
rect 231820 170504 231822 170513
rect 231766 170439 231822 170448
rect 231306 169960 231362 169969
rect 231306 169895 231362 169904
rect 231768 169720 231820 169726
rect 231768 169662 231820 169668
rect 231676 169584 231728 169590
rect 231674 169552 231676 169561
rect 231728 169552 231730 169561
rect 231674 169487 231730 169496
rect 231780 168609 231808 169662
rect 231766 168600 231822 168609
rect 231766 168535 231822 168544
rect 231768 168360 231820 168366
rect 231768 168302 231820 168308
rect 231676 168292 231728 168298
rect 231676 168234 231728 168240
rect 231584 168224 231636 168230
rect 231584 168166 231636 168172
rect 231596 167113 231624 168166
rect 231688 167657 231716 168234
rect 231780 168065 231808 168302
rect 231766 168056 231822 168065
rect 231766 167991 231822 168000
rect 231674 167648 231730 167657
rect 231674 167583 231730 167592
rect 231582 167104 231638 167113
rect 231582 167039 231638 167048
rect 231768 167000 231820 167006
rect 231768 166942 231820 166948
rect 231124 166932 231176 166938
rect 231124 166874 231176 166880
rect 231136 166161 231164 166874
rect 231780 166705 231808 166942
rect 231766 166696 231822 166705
rect 231766 166631 231822 166640
rect 231122 166152 231178 166161
rect 231122 166087 231178 166096
rect 231492 166116 231544 166122
rect 231492 166058 231544 166064
rect 231504 165753 231532 166058
rect 231490 165744 231546 165753
rect 231490 165679 231546 165688
rect 231768 165572 231820 165578
rect 231768 165514 231820 165520
rect 231308 165504 231360 165510
rect 231308 165446 231360 165452
rect 231320 164801 231348 165446
rect 231780 165209 231808 165514
rect 231766 165200 231822 165209
rect 231766 165135 231822 165144
rect 231306 164792 231362 164801
rect 231306 164727 231362 164736
rect 231676 164212 231728 164218
rect 231676 164154 231728 164160
rect 231688 162897 231716 164154
rect 231674 162888 231730 162897
rect 231674 162823 231730 162832
rect 231768 162852 231820 162858
rect 231768 162794 231820 162800
rect 231676 162784 231728 162790
rect 231676 162726 231728 162732
rect 231688 161537 231716 162726
rect 231780 162489 231808 162794
rect 231766 162480 231822 162489
rect 231766 162415 231822 162424
rect 231768 162036 231820 162042
rect 231768 161978 231820 161984
rect 231780 161945 231808 161978
rect 231766 161936 231822 161945
rect 231766 161871 231822 161880
rect 231674 161528 231730 161537
rect 231674 161463 231730 161472
rect 231768 161424 231820 161430
rect 231768 161366 231820 161372
rect 231400 161356 231452 161362
rect 231400 161298 231452 161304
rect 231412 160585 231440 161298
rect 231780 160993 231808 161366
rect 231766 160984 231822 160993
rect 231766 160919 231822 160928
rect 231398 160576 231454 160585
rect 231398 160511 231454 160520
rect 231492 160064 231544 160070
rect 231492 160006 231544 160012
rect 231504 159089 231532 160006
rect 231768 159996 231820 160002
rect 231768 159938 231820 159944
rect 231780 159633 231808 159938
rect 231766 159624 231822 159633
rect 231766 159559 231822 159568
rect 231490 159080 231546 159089
rect 231490 159015 231546 159024
rect 231768 158704 231820 158710
rect 231768 158646 231820 158652
rect 231780 158137 231808 158646
rect 231766 158128 231822 158137
rect 231766 158063 231822 158072
rect 231768 157344 231820 157350
rect 231768 157286 231820 157292
rect 231676 157276 231728 157282
rect 231676 157218 231728 157224
rect 231688 156777 231716 157218
rect 231780 157185 231808 157286
rect 231766 157176 231822 157185
rect 231766 157111 231822 157120
rect 231674 156768 231730 156777
rect 231674 156703 231730 156712
rect 230938 156224 230994 156233
rect 230938 156159 230994 156168
rect 231124 155848 231176 155854
rect 231122 155816 231124 155825
rect 231176 155816 231178 155825
rect 231122 155751 231178 155760
rect 231768 155780 231820 155786
rect 231768 155722 231820 155728
rect 230572 155440 230624 155446
rect 230572 155382 230624 155388
rect 230584 155281 230612 155382
rect 230570 155272 230626 155281
rect 230570 155207 230626 155216
rect 231582 155272 231638 155281
rect 231582 155207 231638 155216
rect 231596 152017 231624 155207
rect 231780 154873 231808 155722
rect 231766 154864 231822 154873
rect 231766 154799 231822 154808
rect 231768 153196 231820 153202
rect 231768 153138 231820 153144
rect 231676 153128 231728 153134
rect 231676 153070 231728 153076
rect 231688 152561 231716 153070
rect 231780 152969 231808 153138
rect 231766 152960 231822 152969
rect 231766 152895 231822 152904
rect 231674 152552 231730 152561
rect 231674 152487 231730 152496
rect 231582 152008 231638 152017
rect 231582 151943 231638 151952
rect 231676 151700 231728 151706
rect 231676 151642 231728 151648
rect 231688 151609 231716 151642
rect 231768 151632 231820 151638
rect 231674 151600 231730 151609
rect 231768 151574 231820 151580
rect 231674 151535 231730 151544
rect 231780 151065 231808 151574
rect 231766 151056 231822 151065
rect 231766 150991 231822 151000
rect 231766 150648 231822 150657
rect 231872 150634 231900 225694
rect 232424 185774 232452 240219
rect 233068 237454 233096 240219
rect 233712 238542 233740 240219
rect 233700 238536 233752 238542
rect 233700 238478 233752 238484
rect 233056 237448 233108 237454
rect 233056 237390 233108 237396
rect 233240 233232 233292 233238
rect 233240 233174 233292 233180
rect 231952 185768 232004 185774
rect 231952 185710 232004 185716
rect 232412 185768 232464 185774
rect 232412 185710 232464 185716
rect 231964 153377 231992 185710
rect 232136 183184 232188 183190
rect 232136 183126 232188 183132
rect 232044 181484 232096 181490
rect 232044 181426 232096 181432
rect 232056 155446 232084 181426
rect 232148 164626 232176 183126
rect 232136 164620 232188 164626
rect 232136 164562 232188 164568
rect 232504 157412 232556 157418
rect 232504 157354 232556 157360
rect 232044 155440 232096 155446
rect 232044 155382 232096 155388
rect 231950 153368 232006 153377
rect 231950 153303 232006 153312
rect 231822 150606 231900 150634
rect 231766 150583 231822 150592
rect 231676 150340 231728 150346
rect 231676 150282 231728 150288
rect 230940 150068 230992 150074
rect 230940 150010 230992 150016
rect 230952 149705 230980 150010
rect 231216 149728 231268 149734
rect 230938 149696 230994 149705
rect 231216 149670 231268 149676
rect 230938 149631 230994 149640
rect 230478 147792 230534 147801
rect 230478 147727 230534 147736
rect 230940 147076 230992 147082
rect 230940 147018 230992 147024
rect 230952 146849 230980 147018
rect 230938 146840 230994 146849
rect 230938 146775 230994 146784
rect 231032 146124 231084 146130
rect 231032 146066 231084 146072
rect 231044 145353 231072 146066
rect 231030 145344 231086 145353
rect 231030 145279 231086 145288
rect 229928 143608 229980 143614
rect 229928 143550 229980 143556
rect 229744 138032 229796 138038
rect 229744 137974 229796 137980
rect 229008 96620 229060 96626
rect 229008 96562 229060 96568
rect 229020 95946 229048 96562
rect 229008 95940 229060 95946
rect 229008 95882 229060 95888
rect 228364 95260 228416 95266
rect 228364 95202 228416 95208
rect 216312 92608 216364 92614
rect 216312 92550 216364 92556
rect 220084 92608 220136 92614
rect 220084 92550 220136 92556
rect 215944 89004 215996 89010
rect 215944 88946 215996 88952
rect 214838 88224 214894 88233
rect 214838 88159 214894 88168
rect 214748 77240 214800 77246
rect 214748 77182 214800 77188
rect 206284 74520 206336 74526
rect 206284 74462 206336 74468
rect 188344 3528 188396 3534
rect 188344 3470 188396 3476
rect 215956 3466 215984 88946
rect 220096 6866 220124 92550
rect 228376 19990 228404 95202
rect 228364 19984 228416 19990
rect 228364 19926 228416 19932
rect 229756 14550 229784 137974
rect 229836 133952 229888 133958
rect 229836 133894 229888 133900
rect 229848 69766 229876 133894
rect 229940 101833 229968 143550
rect 231124 143404 231176 143410
rect 231124 143346 231176 143352
rect 231136 142497 231164 143346
rect 231122 142488 231178 142497
rect 231122 142423 231178 142432
rect 231228 142154 231256 149670
rect 231688 149161 231716 150282
rect 231768 150272 231820 150278
rect 231768 150214 231820 150220
rect 231780 150113 231808 150214
rect 231766 150104 231822 150113
rect 231766 150039 231822 150048
rect 231674 149152 231730 149161
rect 231674 149087 231730 149096
rect 231768 149048 231820 149054
rect 231768 148990 231820 148996
rect 231780 148209 231808 148990
rect 231766 148200 231822 148209
rect 231766 148135 231822 148144
rect 231768 147620 231820 147626
rect 231768 147562 231820 147568
rect 231780 147257 231808 147562
rect 231766 147248 231822 147257
rect 231766 147183 231822 147192
rect 231766 146296 231822 146305
rect 231766 146231 231768 146240
rect 231820 146231 231822 146240
rect 231768 146202 231820 146208
rect 231676 146192 231728 146198
rect 231676 146134 231728 146140
rect 231688 145897 231716 146134
rect 231674 145888 231730 145897
rect 231674 145823 231730 145832
rect 231766 145616 231822 145625
rect 231766 145551 231822 145560
rect 231584 144900 231636 144906
rect 231584 144842 231636 144848
rect 231596 143993 231624 144842
rect 231780 144401 231808 145551
rect 231766 144392 231822 144401
rect 231766 144327 231822 144336
rect 231582 143984 231638 143993
rect 231582 143919 231638 143928
rect 231676 143540 231728 143546
rect 231676 143482 231728 143488
rect 231688 143041 231716 143482
rect 231768 143472 231820 143478
rect 231766 143440 231768 143449
rect 231820 143440 231822 143449
rect 231766 143375 231822 143384
rect 231674 143032 231730 143041
rect 231674 142967 231730 142976
rect 231136 142126 231256 142154
rect 231032 135108 231084 135114
rect 231032 135050 231084 135056
rect 231044 134065 231072 135050
rect 231030 134056 231086 134065
rect 231030 133991 231086 134000
rect 230940 133816 230992 133822
rect 230940 133758 230992 133764
rect 230952 133113 230980 133758
rect 230938 133104 230994 133113
rect 230938 133039 230994 133048
rect 231136 132494 231164 142126
rect 231768 142112 231820 142118
rect 231768 142054 231820 142060
rect 231308 141500 231360 141506
rect 231308 141442 231360 141448
rect 231216 138712 231268 138718
rect 231216 138654 231268 138660
rect 231044 132466 231164 132494
rect 231044 126041 231072 132466
rect 231124 126948 231176 126954
rect 231124 126890 231176 126896
rect 231136 126449 231164 126890
rect 231122 126440 231178 126449
rect 231122 126375 231178 126384
rect 231030 126032 231086 126041
rect 231030 125967 231086 125976
rect 230848 124908 230900 124914
rect 230848 124850 230900 124856
rect 230756 123548 230808 123554
rect 230756 123490 230808 123496
rect 230664 118652 230716 118658
rect 230664 118594 230716 118600
rect 230676 118425 230704 118594
rect 230662 118416 230718 118425
rect 230662 118351 230718 118360
rect 230664 117292 230716 117298
rect 230664 117234 230716 117240
rect 230676 117065 230704 117234
rect 230662 117056 230718 117065
rect 230662 116991 230718 117000
rect 230572 116544 230624 116550
rect 230570 116512 230572 116521
rect 230624 116512 230626 116521
rect 230570 116447 230626 116456
rect 230768 116113 230796 123490
rect 230860 121689 230888 124850
rect 231228 122834 231256 138654
rect 231320 131617 231348 141442
rect 231780 141137 231808 142054
rect 231766 141128 231822 141137
rect 231766 141063 231822 141072
rect 231676 140752 231728 140758
rect 231676 140694 231728 140700
rect 231766 140720 231822 140729
rect 231688 140185 231716 140694
rect 231766 140655 231768 140664
rect 231820 140655 231822 140664
rect 231768 140626 231820 140632
rect 231674 140176 231730 140185
rect 231674 140111 231730 140120
rect 231400 137964 231452 137970
rect 231400 137906 231452 137912
rect 231412 137329 231440 137906
rect 231768 137896 231820 137902
rect 231768 137838 231820 137844
rect 231398 137320 231454 137329
rect 231398 137255 231454 137264
rect 231584 137284 231636 137290
rect 231584 137226 231636 137232
rect 231400 136604 231452 136610
rect 231400 136546 231452 136552
rect 231412 135969 231440 136546
rect 231398 135960 231454 135969
rect 231398 135895 231454 135904
rect 231492 135244 231544 135250
rect 231492 135186 231544 135192
rect 231504 134473 231532 135186
rect 231490 134464 231546 134473
rect 231490 134399 231546 134408
rect 231596 133521 231624 137226
rect 231780 136921 231808 137838
rect 231766 136912 231822 136921
rect 231766 136847 231822 136856
rect 231768 136536 231820 136542
rect 231768 136478 231820 136484
rect 231780 135425 231808 136478
rect 231766 135416 231822 135425
rect 231766 135351 231822 135360
rect 231676 133884 231728 133890
rect 231676 133826 231728 133832
rect 231582 133512 231638 133521
rect 231582 133447 231638 133456
rect 231688 132569 231716 133826
rect 231674 132560 231730 132569
rect 231674 132495 231730 132504
rect 231768 132456 231820 132462
rect 231768 132398 231820 132404
rect 231676 132388 231728 132394
rect 231676 132330 231728 132336
rect 231306 131608 231362 131617
rect 231306 131543 231362 131552
rect 231688 131209 231716 132330
rect 231780 132161 231808 132398
rect 231766 132152 231822 132161
rect 231766 132087 231822 132096
rect 231674 131200 231730 131209
rect 231492 131164 231544 131170
rect 231674 131135 231730 131144
rect 231492 131106 231544 131112
rect 231400 131028 231452 131034
rect 231400 130970 231452 130976
rect 231412 130257 231440 130970
rect 231398 130248 231454 130257
rect 231398 130183 231454 130192
rect 231308 129736 231360 129742
rect 231308 129678 231360 129684
rect 231320 129305 231348 129678
rect 231306 129296 231362 129305
rect 231306 129231 231362 129240
rect 231504 128897 231532 131106
rect 231768 131096 231820 131102
rect 231768 131038 231820 131044
rect 231676 130960 231728 130966
rect 231676 130902 231728 130908
rect 231688 129849 231716 130902
rect 231780 130665 231808 131038
rect 231766 130656 231822 130665
rect 231766 130591 231822 130600
rect 231674 129840 231730 129849
rect 231674 129775 231730 129784
rect 231584 129056 231636 129062
rect 231584 128998 231636 129004
rect 231490 128888 231546 128897
rect 231490 128823 231546 128832
rect 231492 126268 231544 126274
rect 231492 126210 231544 126216
rect 231308 124976 231360 124982
rect 231308 124918 231360 124924
rect 231320 124545 231348 124918
rect 231306 124536 231362 124545
rect 231306 124471 231362 124480
rect 231136 122806 231256 122834
rect 230846 121680 230902 121689
rect 230846 121615 230902 121624
rect 230940 121372 230992 121378
rect 230940 121314 230992 121320
rect 230952 120737 230980 121314
rect 230938 120728 230994 120737
rect 230938 120663 230994 120672
rect 231136 120329 231164 122806
rect 231308 122800 231360 122806
rect 231308 122742 231360 122748
rect 231320 122233 231348 122742
rect 231504 122641 231532 126210
rect 231596 124137 231624 128998
rect 231766 128344 231822 128353
rect 231676 128308 231728 128314
rect 231766 128279 231822 128288
rect 231676 128250 231728 128256
rect 231688 127945 231716 128250
rect 231780 128246 231808 128279
rect 231768 128240 231820 128246
rect 231768 128182 231820 128188
rect 231674 127936 231730 127945
rect 231674 127871 231730 127880
rect 231676 127832 231728 127838
rect 231676 127774 231728 127780
rect 231688 127401 231716 127774
rect 231674 127392 231730 127401
rect 231674 127327 231730 127336
rect 231766 126984 231822 126993
rect 231766 126919 231822 126928
rect 231780 126886 231808 126919
rect 231768 126880 231820 126886
rect 231768 126822 231820 126828
rect 231768 125588 231820 125594
rect 231768 125530 231820 125536
rect 231780 125089 231808 125530
rect 231766 125080 231822 125089
rect 231766 125015 231822 125024
rect 231768 124160 231820 124166
rect 231582 124128 231638 124137
rect 231768 124102 231820 124108
rect 231582 124063 231638 124072
rect 231584 123616 231636 123622
rect 231582 123584 231584 123593
rect 231636 123584 231638 123593
rect 231582 123519 231638 123528
rect 231780 123185 231808 124102
rect 231766 123176 231822 123185
rect 231766 123111 231822 123120
rect 231490 122632 231546 122641
rect 231490 122567 231546 122576
rect 231306 122224 231362 122233
rect 231306 122159 231362 122168
rect 231676 122120 231728 122126
rect 231676 122062 231728 122068
rect 231216 120760 231268 120766
rect 231216 120702 231268 120708
rect 231122 120320 231178 120329
rect 231122 120255 231178 120264
rect 230940 120080 230992 120086
rect 230940 120022 230992 120028
rect 230952 119785 230980 120022
rect 230938 119776 230994 119785
rect 230938 119711 230994 119720
rect 230940 117564 230992 117570
rect 230940 117506 230992 117512
rect 230952 117473 230980 117506
rect 230938 117464 230994 117473
rect 230938 117399 230994 117408
rect 231228 116906 231256 120702
rect 231492 120012 231544 120018
rect 231492 119954 231544 119960
rect 231504 118969 231532 119954
rect 231490 118960 231546 118969
rect 231490 118895 231546 118904
rect 231136 116878 231256 116906
rect 230754 116104 230810 116113
rect 230754 116039 230810 116048
rect 230572 114504 230624 114510
rect 230572 114446 230624 114452
rect 230584 113257 230612 114446
rect 230664 114436 230716 114442
rect 230664 114378 230716 114384
rect 230676 114209 230704 114378
rect 230662 114200 230718 114209
rect 230662 114135 230718 114144
rect 230570 113248 230626 113257
rect 230570 113183 230626 113192
rect 231136 113174 231164 116878
rect 231216 116612 231268 116618
rect 231216 116554 231268 116560
rect 230940 113144 230992 113150
rect 230940 113086 230992 113092
rect 231044 113146 231164 113174
rect 231228 113174 231256 116554
rect 231584 115252 231636 115258
rect 231584 115194 231636 115200
rect 231492 114368 231544 114374
rect 231492 114310 231544 114316
rect 231504 113665 231532 114310
rect 231490 113656 231546 113665
rect 231490 113591 231546 113600
rect 231228 113146 231348 113174
rect 230952 112713 230980 113086
rect 230938 112704 230994 112713
rect 230938 112639 230994 112648
rect 230848 108180 230900 108186
rect 230848 108122 230900 108128
rect 230572 107568 230624 107574
rect 230572 107510 230624 107516
rect 230584 106593 230612 107510
rect 230570 106584 230626 106593
rect 230570 106519 230626 106528
rect 230480 105596 230532 105602
rect 230480 105538 230532 105544
rect 229926 101824 229982 101833
rect 229926 101759 229982 101768
rect 230492 97617 230520 105538
rect 230860 105233 230888 108122
rect 230846 105224 230902 105233
rect 230846 105159 230902 105168
rect 230664 103828 230716 103834
rect 230664 103770 230716 103776
rect 230572 102128 230624 102134
rect 230572 102070 230624 102076
rect 230584 100881 230612 102070
rect 230570 100872 230626 100881
rect 230570 100807 230626 100816
rect 230676 98977 230704 103770
rect 231044 103737 231072 113146
rect 231124 110356 231176 110362
rect 231124 110298 231176 110304
rect 231136 109857 231164 110298
rect 231122 109848 231178 109857
rect 231122 109783 231178 109792
rect 231124 108996 231176 109002
rect 231124 108938 231176 108944
rect 231136 108497 231164 108938
rect 231122 108488 231178 108497
rect 231122 108423 231178 108432
rect 231030 103728 231086 103737
rect 231030 103663 231086 103672
rect 231320 102377 231348 113146
rect 231492 112464 231544 112470
rect 231492 112406 231544 112412
rect 231504 109449 231532 112406
rect 231596 110809 231624 115194
rect 231688 114617 231716 122062
rect 231768 121440 231820 121446
rect 231768 121382 231820 121388
rect 231780 121281 231808 121382
rect 231766 121272 231822 121281
rect 231766 121207 231822 121216
rect 231768 119944 231820 119950
rect 231768 119886 231820 119892
rect 231780 119377 231808 119886
rect 231766 119368 231822 119377
rect 231766 119303 231822 119312
rect 231768 118584 231820 118590
rect 231768 118526 231820 118532
rect 231780 118017 231808 118526
rect 231766 118008 231822 118017
rect 231766 117943 231822 117952
rect 232516 116550 232544 157354
rect 233252 155854 233280 233174
rect 233332 223576 233384 223582
rect 233332 223518 233384 223524
rect 233240 155848 233292 155854
rect 233240 155790 233292 155796
rect 232780 148368 232832 148374
rect 232780 148310 232832 148316
rect 232596 146940 232648 146946
rect 232596 146882 232648 146888
rect 232504 116544 232556 116550
rect 232504 116486 232556 116492
rect 231768 115932 231820 115938
rect 231768 115874 231820 115880
rect 231780 115569 231808 115874
rect 231766 115560 231822 115569
rect 231766 115495 231822 115504
rect 231768 115184 231820 115190
rect 231766 115152 231768 115161
rect 231820 115152 231822 115161
rect 231766 115087 231822 115096
rect 231674 114608 231730 114617
rect 231674 114543 231730 114552
rect 231676 112736 231728 112742
rect 231676 112678 231728 112684
rect 231688 112305 231716 112678
rect 231674 112296 231730 112305
rect 231674 112231 231730 112240
rect 231768 111784 231820 111790
rect 231766 111752 231768 111761
rect 231820 111752 231822 111761
rect 231676 111716 231728 111722
rect 231766 111687 231822 111696
rect 231676 111658 231728 111664
rect 231688 111353 231716 111658
rect 231674 111344 231730 111353
rect 231674 111279 231730 111288
rect 231676 111104 231728 111110
rect 231676 111046 231728 111052
rect 231582 110800 231638 110809
rect 231582 110735 231638 110744
rect 231490 109440 231546 109449
rect 231490 109375 231546 109384
rect 231584 109132 231636 109138
rect 231584 109074 231636 109080
rect 231596 107137 231624 109074
rect 231688 107953 231716 111046
rect 231768 110424 231820 110430
rect 231766 110392 231768 110401
rect 231820 110392 231822 110401
rect 231766 110327 231822 110336
rect 231768 108928 231820 108934
rect 231766 108896 231768 108905
rect 231820 108896 231822 108905
rect 231766 108831 231822 108840
rect 231674 107944 231730 107953
rect 231674 107879 231730 107888
rect 231768 107636 231820 107642
rect 231768 107578 231820 107584
rect 231780 107545 231808 107578
rect 232608 107574 232636 146882
rect 232688 146328 232740 146334
rect 232688 146270 232740 146276
rect 232700 108186 232728 146270
rect 232792 114510 232820 148310
rect 233344 147082 233372 223518
rect 234356 193866 234384 240219
rect 234344 193860 234396 193866
rect 234344 193802 234396 193808
rect 233424 191208 233476 191214
rect 233424 191150 233476 191156
rect 233436 150074 233464 191150
rect 234620 183116 234672 183122
rect 234620 183058 234672 183064
rect 234632 166938 234660 183058
rect 235000 181529 235028 240219
rect 235644 238134 235672 240219
rect 235632 238128 235684 238134
rect 235632 238070 235684 238076
rect 235264 225616 235316 225622
rect 235264 225558 235316 225564
rect 234986 181520 235042 181529
rect 234986 181455 235042 181464
rect 234712 180328 234764 180334
rect 234712 180270 234764 180276
rect 234620 166932 234672 166938
rect 234620 166874 234672 166880
rect 234724 165510 234752 180270
rect 235276 171766 235304 225558
rect 236288 187066 236316 240219
rect 236932 239970 236960 240219
rect 236920 239964 236972 239970
rect 236920 239906 236972 239912
rect 237380 237448 237432 237454
rect 237380 237390 237432 237396
rect 236276 187060 236328 187066
rect 236276 187002 236328 187008
rect 236000 185904 236052 185910
rect 236000 185846 236052 185852
rect 235356 175296 235408 175302
rect 235356 175238 235408 175244
rect 235264 171760 235316 171766
rect 235264 171702 235316 171708
rect 234712 165504 234764 165510
rect 234712 165446 234764 165452
rect 235264 162920 235316 162926
rect 235264 162862 235316 162868
rect 234160 153264 234212 153270
rect 234160 153206 234212 153212
rect 233790 151056 233846 151065
rect 233790 150991 233846 151000
rect 233424 150068 233476 150074
rect 233424 150010 233476 150016
rect 233332 147076 233384 147082
rect 233332 147018 233384 147024
rect 233804 143410 233832 150991
rect 234068 146396 234120 146402
rect 234068 146338 234120 146344
rect 233976 145104 234028 145110
rect 233976 145046 234028 145052
rect 233792 143404 233844 143410
rect 233792 143346 233844 143352
rect 233884 142860 233936 142866
rect 233884 142802 233936 142808
rect 233896 124982 233924 142802
rect 233884 124976 233936 124982
rect 233884 124918 233936 124924
rect 233884 121508 233936 121514
rect 233884 121450 233936 121456
rect 232780 114504 232832 114510
rect 232780 114446 232832 114452
rect 232688 108180 232740 108186
rect 232688 108122 232740 108128
rect 232596 107568 232648 107574
rect 231766 107536 231822 107545
rect 232596 107510 232648 107516
rect 231766 107471 231822 107480
rect 231582 107128 231638 107137
rect 231582 107063 231638 107072
rect 231400 106956 231452 106962
rect 231400 106898 231452 106904
rect 231306 102368 231362 102377
rect 231306 102303 231362 102312
rect 231124 102060 231176 102066
rect 231124 102002 231176 102008
rect 231136 101425 231164 102002
rect 231122 101416 231178 101425
rect 231122 101351 231178 101360
rect 231412 99521 231440 106898
rect 231768 106276 231820 106282
rect 231768 106218 231820 106224
rect 231676 106208 231728 106214
rect 231674 106176 231676 106185
rect 231728 106176 231730 106185
rect 231674 106111 231730 106120
rect 231780 105641 231808 106218
rect 231766 105632 231822 105641
rect 231766 105567 231822 105576
rect 231768 104848 231820 104854
rect 231768 104790 231820 104796
rect 231584 104712 231636 104718
rect 231582 104680 231584 104689
rect 231636 104680 231638 104689
rect 231582 104615 231638 104624
rect 231780 104281 231808 104790
rect 231766 104272 231822 104281
rect 231766 104207 231822 104216
rect 231768 103488 231820 103494
rect 231768 103430 231820 103436
rect 231584 103352 231636 103358
rect 231582 103320 231584 103329
rect 231636 103320 231638 103329
rect 231582 103255 231638 103264
rect 231780 102785 231808 103430
rect 231766 102776 231822 102785
rect 231766 102711 231822 102720
rect 232504 102196 232556 102202
rect 232504 102138 232556 102144
rect 231676 100700 231728 100706
rect 231676 100642 231728 100648
rect 231688 99929 231716 100642
rect 231768 100632 231820 100638
rect 231768 100574 231820 100580
rect 231780 100473 231808 100574
rect 231766 100464 231822 100473
rect 231766 100399 231822 100408
rect 231674 99920 231730 99929
rect 231674 99855 231730 99864
rect 231398 99512 231454 99521
rect 231398 99447 231454 99456
rect 231492 99340 231544 99346
rect 231492 99282 231544 99288
rect 230662 98968 230718 98977
rect 230662 98903 230718 98912
rect 231504 98569 231532 99282
rect 231490 98560 231546 98569
rect 231490 98495 231546 98504
rect 230478 97608 230534 97617
rect 230478 97543 230534 97552
rect 230478 97064 230534 97073
rect 230478 96999 230534 97008
rect 230492 95946 230520 96999
rect 231122 96656 231178 96665
rect 231122 96591 231178 96600
rect 230480 95940 230532 95946
rect 230480 95882 230532 95888
rect 230478 95704 230534 95713
rect 230478 95639 230534 95648
rect 230492 93226 230520 95639
rect 231136 93838 231164 96591
rect 231124 93832 231176 93838
rect 231124 93774 231176 93780
rect 230480 93220 230532 93226
rect 230480 93162 230532 93168
rect 229836 69760 229888 69766
rect 229836 69702 229888 69708
rect 231136 58682 231164 93774
rect 231124 58676 231176 58682
rect 231124 58618 231176 58624
rect 229744 14544 229796 14550
rect 229744 14486 229796 14492
rect 220084 6860 220136 6866
rect 220084 6802 220136 6808
rect 232516 6186 232544 102138
rect 233896 17270 233924 121450
rect 233988 103358 234016 145046
rect 234080 104718 234108 146338
rect 234172 112742 234200 153206
rect 234528 152516 234580 152522
rect 234528 152458 234580 152464
rect 234540 151706 234568 152458
rect 234528 151700 234580 151706
rect 234528 151642 234580 151648
rect 235276 123622 235304 162862
rect 235264 123616 235316 123622
rect 235264 123558 235316 123564
rect 235264 113212 235316 113218
rect 235264 113154 235316 113160
rect 234160 112736 234212 112742
rect 234160 112678 234212 112684
rect 234068 104712 234120 104718
rect 234068 104654 234120 104660
rect 233976 103352 234028 103358
rect 233976 103294 234028 103300
rect 234068 96688 234120 96694
rect 234068 96630 234120 96636
rect 233976 93220 234028 93226
rect 233976 93162 234028 93168
rect 233884 17264 233936 17270
rect 233884 17206 233936 17212
rect 232504 6180 232556 6186
rect 232504 6122 232556 6128
rect 233988 3534 234016 93162
rect 234080 49026 234108 96630
rect 234068 49020 234120 49026
rect 234068 48962 234120 48968
rect 235276 35222 235304 113154
rect 235368 103834 235396 175238
rect 236012 173738 236040 185846
rect 236092 177540 236144 177546
rect 236092 177482 236144 177488
rect 236000 173732 236052 173738
rect 236000 173674 236052 173680
rect 235540 168428 235592 168434
rect 235540 168370 235592 168376
rect 235448 147688 235500 147694
rect 235448 147630 235500 147636
rect 235460 109138 235488 147630
rect 235552 131170 235580 168370
rect 236104 166122 236132 177482
rect 236276 177404 236328 177410
rect 236276 177346 236328 177352
rect 236184 176112 236236 176118
rect 236184 176054 236236 176060
rect 236196 170610 236224 176054
rect 236184 170604 236236 170610
rect 236184 170546 236236 170552
rect 236288 170542 236316 177346
rect 236828 172576 236880 172582
rect 236828 172518 236880 172524
rect 236276 170536 236328 170542
rect 236276 170478 236328 170484
rect 236644 170400 236696 170406
rect 236644 170342 236696 170348
rect 236092 166116 236144 166122
rect 236092 166058 236144 166064
rect 236656 135114 236684 170342
rect 236736 157480 236788 157486
rect 236736 157422 236788 157428
rect 236644 135108 236696 135114
rect 236644 135050 236696 135056
rect 236644 132524 236696 132530
rect 236644 132466 236696 132472
rect 235540 131164 235592 131170
rect 235540 131106 235592 131112
rect 235448 109132 235500 109138
rect 235448 109074 235500 109080
rect 235908 104168 235960 104174
rect 235908 104110 235960 104116
rect 235356 103828 235408 103834
rect 235356 103770 235408 103776
rect 235920 102066 235948 104110
rect 235908 102060 235960 102066
rect 235908 102002 235960 102008
rect 235356 98048 235408 98054
rect 235356 97990 235408 97996
rect 235368 50386 235396 97990
rect 235356 50380 235408 50386
rect 235356 50322 235408 50328
rect 236656 40730 236684 132466
rect 236748 117570 236776 157422
rect 236840 133822 236868 172518
rect 237392 169590 237420 237390
rect 237576 234598 237604 240219
rect 237564 234592 237616 234598
rect 237564 234534 237616 234540
rect 237472 180396 237524 180402
rect 237472 180338 237524 180344
rect 237380 169584 237432 169590
rect 237380 169526 237432 169532
rect 236920 164892 236972 164898
rect 236920 164834 236972 164840
rect 236828 133816 236880 133822
rect 236828 133758 236880 133764
rect 236932 127838 236960 164834
rect 237484 146130 237512 180338
rect 237564 176044 237616 176050
rect 237564 175986 237616 175992
rect 237576 162042 237604 175986
rect 238220 175982 238248 240219
rect 238760 239828 238812 239834
rect 238760 239770 238812 239776
rect 238772 239737 238800 239770
rect 238758 239728 238814 239737
rect 238758 239663 238814 239672
rect 238864 186998 238892 240219
rect 240152 218754 240180 240219
rect 240796 220114 240824 240219
rect 240784 220108 240836 220114
rect 240784 220050 240836 220056
rect 240140 218748 240192 218754
rect 240140 218690 240192 218696
rect 238852 186992 238904 186998
rect 238852 186934 238904 186940
rect 240232 185836 240284 185842
rect 240232 185778 240284 185784
rect 238852 178900 238904 178906
rect 238852 178842 238904 178848
rect 238760 177472 238812 177478
rect 238760 177414 238812 177420
rect 238208 175976 238260 175982
rect 238208 175918 238260 175924
rect 238024 173936 238076 173942
rect 238024 173878 238076 173884
rect 237564 162036 237616 162042
rect 237564 161978 237616 161984
rect 237472 146124 237524 146130
rect 237472 146066 237524 146072
rect 238036 135289 238064 173878
rect 238300 161492 238352 161498
rect 238300 161434 238352 161440
rect 238208 155984 238260 155990
rect 238208 155926 238260 155932
rect 238116 135312 238168 135318
rect 238022 135280 238078 135289
rect 238116 135254 238168 135260
rect 238022 135215 238078 135224
rect 236920 127832 236972 127838
rect 236920 127774 236972 127780
rect 238024 120148 238076 120154
rect 238024 120090 238076 120096
rect 236736 117564 236788 117570
rect 236736 117506 236788 117512
rect 236644 40724 236696 40730
rect 236644 40666 236696 40672
rect 235264 35216 235316 35222
rect 235264 35158 235316 35164
rect 238036 4826 238064 120090
rect 238128 32502 238156 135254
rect 238220 115190 238248 155926
rect 238312 121378 238340 161434
rect 238772 151638 238800 177414
rect 238864 162790 238892 178842
rect 239680 167068 239732 167074
rect 239680 167010 239732 167016
rect 238852 162784 238904 162790
rect 238852 162726 238904 162732
rect 239496 160132 239548 160138
rect 239496 160074 239548 160080
rect 238760 151632 238812 151638
rect 238760 151574 238812 151580
rect 238392 145580 238444 145586
rect 238392 145522 238444 145528
rect 238300 121372 238352 121378
rect 238300 121314 238352 121320
rect 238208 115184 238260 115190
rect 238208 115126 238260 115132
rect 238404 106214 238432 145522
rect 239404 136672 239456 136678
rect 239404 136614 239456 136620
rect 238392 106208 238444 106214
rect 238392 106150 238444 106156
rect 238208 100768 238260 100774
rect 238208 100710 238260 100716
rect 238116 32496 238168 32502
rect 238116 32438 238168 32444
rect 238220 25566 238248 100710
rect 238208 25560 238260 25566
rect 238208 25502 238260 25508
rect 239416 11762 239444 136614
rect 239508 119950 239536 160074
rect 239588 154624 239640 154630
rect 239588 154566 239640 154572
rect 239496 119944 239548 119950
rect 239496 119886 239548 119892
rect 239496 117360 239548 117366
rect 239496 117302 239548 117308
rect 239508 31142 239536 117302
rect 239600 114442 239628 154566
rect 239692 126886 239720 167010
rect 240244 160002 240272 185778
rect 240876 168564 240928 168570
rect 240876 168506 240928 168512
rect 240784 166320 240836 166326
rect 240784 166262 240836 166268
rect 240232 159996 240284 160002
rect 240232 159938 240284 159944
rect 240796 129742 240824 166262
rect 240784 129736 240836 129742
rect 240784 129678 240836 129684
rect 240888 128246 240916 168506
rect 241152 153332 241204 153338
rect 241152 153274 241204 153280
rect 241060 151972 241112 151978
rect 241060 151914 241112 151920
rect 240876 128240 240928 128246
rect 240876 128182 240928 128188
rect 240784 127016 240836 127022
rect 240784 126958 240836 126964
rect 239680 126880 239732 126886
rect 239680 126822 239732 126828
rect 239588 114436 239640 114442
rect 239588 114378 239640 114384
rect 239496 31136 239548 31142
rect 239496 31078 239548 31084
rect 240796 21418 240824 126958
rect 240876 124228 240928 124234
rect 240876 124170 240928 124176
rect 240888 46238 240916 124170
rect 240968 111852 241020 111858
rect 240968 111794 241020 111800
rect 240980 55894 241008 111794
rect 241072 111722 241100 151914
rect 241164 113150 241192 153274
rect 241440 153241 241468 240219
rect 241426 153232 241482 153241
rect 241426 153167 241482 153176
rect 242084 152522 242112 240219
rect 242728 240038 242756 240219
rect 242716 240032 242768 240038
rect 242716 239974 242768 239980
rect 242164 235408 242216 235414
rect 242164 235350 242216 235356
rect 242176 164218 242204 235350
rect 243372 181490 243400 240219
rect 244024 240038 244052 240219
rect 244012 240032 244064 240038
rect 244012 239974 244064 239980
rect 244660 235890 244688 240219
rect 245016 239420 245068 239426
rect 245016 239362 245068 239368
rect 244924 236768 244976 236774
rect 244924 236710 244976 236716
rect 244648 235884 244700 235890
rect 244648 235826 244700 235832
rect 243544 235340 243596 235346
rect 243544 235282 243596 235288
rect 243360 181484 243412 181490
rect 243360 181426 243412 181432
rect 242992 180192 243044 180198
rect 242992 180134 243044 180140
rect 242900 176180 242952 176186
rect 242900 176122 242952 176128
rect 242256 164280 242308 164286
rect 242256 164222 242308 164228
rect 242164 164212 242216 164218
rect 242164 164154 242216 164160
rect 242164 158772 242216 158778
rect 242164 158714 242216 158720
rect 242072 152516 242124 152522
rect 242072 152458 242124 152464
rect 242176 118590 242204 158714
rect 242268 125594 242296 164222
rect 242348 162988 242400 162994
rect 242348 162930 242400 162936
rect 242360 126274 242388 162930
rect 242912 137902 242940 176122
rect 243004 146198 243032 180134
rect 243556 149054 243584 235282
rect 244372 183048 244424 183054
rect 244372 182990 244424 182996
rect 244280 178832 244332 178838
rect 244280 178774 244332 178780
rect 243636 172644 243688 172650
rect 243636 172586 243688 172592
rect 243544 149048 243596 149054
rect 243544 148990 243596 148996
rect 242992 146192 243044 146198
rect 242992 146134 243044 146140
rect 243544 138100 243596 138106
rect 243544 138042 243596 138048
rect 242900 137896 242952 137902
rect 242900 137838 242952 137844
rect 242348 126268 242400 126274
rect 242348 126210 242400 126216
rect 242532 126268 242584 126274
rect 242532 126210 242584 126216
rect 242256 125588 242308 125594
rect 242256 125530 242308 125536
rect 242256 123480 242308 123486
rect 242256 123422 242308 123428
rect 242164 118584 242216 118590
rect 242164 118526 242216 118532
rect 241152 113144 241204 113150
rect 241152 113086 241204 113092
rect 242164 111920 242216 111926
rect 242164 111862 242216 111868
rect 241060 111716 241112 111722
rect 241060 111658 241112 111664
rect 241060 107908 241112 107914
rect 241060 107850 241112 107856
rect 241072 60110 241100 107850
rect 241060 60104 241112 60110
rect 241060 60046 241112 60052
rect 240968 55888 241020 55894
rect 240968 55830 241020 55836
rect 240876 46232 240928 46238
rect 240876 46174 240928 46180
rect 242176 28286 242204 111862
rect 242268 102134 242296 123422
rect 242256 102128 242308 102134
rect 242256 102070 242308 102076
rect 242440 100836 242492 100842
rect 242440 100778 242492 100784
rect 242348 98116 242400 98122
rect 242348 98058 242400 98064
rect 242256 96756 242308 96762
rect 242256 96698 242308 96704
rect 242268 47598 242296 96698
rect 242360 53106 242388 98058
rect 242452 61402 242480 100778
rect 242544 99346 242572 126210
rect 242532 99340 242584 99346
rect 242532 99282 242584 99288
rect 242440 61396 242492 61402
rect 242440 61338 242492 61344
rect 242348 53100 242400 53106
rect 242348 53042 242400 53048
rect 242256 47592 242308 47598
rect 242256 47534 242308 47540
rect 242164 28280 242216 28286
rect 242164 28222 242216 28228
rect 240784 21412 240836 21418
rect 240784 21354 240836 21360
rect 243556 13190 243584 138042
rect 243648 137290 243676 172586
rect 244292 146266 244320 178774
rect 244384 153134 244412 182990
rect 244936 167006 244964 236710
rect 245028 175166 245056 239362
rect 245304 237386 245332 240219
rect 245292 237380 245344 237386
rect 245292 237322 245344 237328
rect 245948 188494 245976 240219
rect 246304 238808 246356 238814
rect 246304 238750 246356 238756
rect 245936 188488 245988 188494
rect 245936 188430 245988 188436
rect 245016 175160 245068 175166
rect 245016 175102 245068 175108
rect 245016 168496 245068 168502
rect 245016 168438 245068 168444
rect 244924 167000 244976 167006
rect 244924 166942 244976 166948
rect 245028 161362 245056 168438
rect 245108 165640 245160 165646
rect 245108 165582 245160 165588
rect 245016 161356 245068 161362
rect 245016 161298 245068 161304
rect 244924 160200 244976 160206
rect 244924 160142 244976 160148
rect 244372 153128 244424 153134
rect 244372 153070 244424 153076
rect 244280 146260 244332 146266
rect 244280 146202 244332 146208
rect 243728 142316 243780 142322
rect 243728 142258 243780 142264
rect 243636 137284 243688 137290
rect 243636 137226 243688 137232
rect 243740 100638 243768 142258
rect 244936 138718 244964 160142
rect 245120 149734 245148 165582
rect 246316 155786 246344 238750
rect 246396 169788 246448 169794
rect 246396 169730 246448 169736
rect 246304 155780 246356 155786
rect 246304 155722 246356 155728
rect 245200 152516 245252 152522
rect 245200 152458 245252 152464
rect 245108 149728 245160 149734
rect 245108 149670 245160 149676
rect 245016 149116 245068 149122
rect 245016 149058 245068 149064
rect 244924 138712 244976 138718
rect 244924 138654 244976 138660
rect 244924 128376 244976 128382
rect 244924 128318 244976 128324
rect 243728 100632 243780 100638
rect 243728 100574 243780 100580
rect 243636 99408 243688 99414
rect 243636 99350 243688 99356
rect 243648 15910 243676 99350
rect 244936 18630 244964 128318
rect 245028 111110 245056 149058
rect 245212 114374 245240 152458
rect 245292 141432 245344 141438
rect 245292 141374 245344 141380
rect 245200 114368 245252 114374
rect 245200 114310 245252 114316
rect 245108 113280 245160 113286
rect 245108 113222 245160 113228
rect 245016 111104 245068 111110
rect 245016 111046 245068 111052
rect 245016 103556 245068 103562
rect 245016 103498 245068 103504
rect 244924 18624 244976 18630
rect 244924 18566 244976 18572
rect 243636 15904 243688 15910
rect 243636 15846 243688 15852
rect 243544 13184 243596 13190
rect 243544 13126 243596 13132
rect 239404 11756 239456 11762
rect 239404 11698 239456 11704
rect 245028 8974 245056 103498
rect 245120 39370 245148 113222
rect 245200 110492 245252 110498
rect 245200 110434 245252 110440
rect 245212 68406 245240 110434
rect 245304 104854 245332 141374
rect 246408 132394 246436 169730
rect 246592 168502 246620 240219
rect 247236 238542 247264 240219
rect 247224 238536 247276 238542
rect 247224 238478 247276 238484
rect 247880 235278 247908 240219
rect 248532 240009 248560 240219
rect 249064 240168 249116 240174
rect 249064 240110 249116 240116
rect 248518 240000 248574 240009
rect 248518 239935 248574 239944
rect 247868 235272 247920 235278
rect 247868 235214 247920 235220
rect 247040 182980 247092 182986
rect 247040 182922 247092 182928
rect 246580 168496 246632 168502
rect 246580 168438 246632 168444
rect 246488 167680 246540 167686
rect 246488 167622 246540 167628
rect 246396 132388 246448 132394
rect 246396 132330 246448 132336
rect 246304 131164 246356 131170
rect 246304 131106 246356 131112
rect 245292 104848 245344 104854
rect 245292 104790 245344 104796
rect 245200 68400 245252 68406
rect 245200 68342 245252 68348
rect 245108 39364 245160 39370
rect 245108 39306 245160 39312
rect 246316 37942 246344 131106
rect 246500 130966 246528 167622
rect 246672 156052 246724 156058
rect 246672 155994 246724 156000
rect 246580 150476 246632 150482
rect 246580 150418 246632 150424
rect 246488 130960 246540 130966
rect 246488 130902 246540 130908
rect 246396 116000 246448 116006
rect 246396 115942 246448 115948
rect 246304 37936 246356 37942
rect 246304 37878 246356 37884
rect 246408 29646 246436 115942
rect 246488 114572 246540 114578
rect 246488 114514 246540 114520
rect 246500 64190 246528 114514
rect 246592 108934 246620 150418
rect 246684 115938 246712 155994
rect 247052 140690 247080 182922
rect 247868 174004 247920 174010
rect 247868 173946 247920 173952
rect 247684 171148 247736 171154
rect 247684 171090 247736 171096
rect 247040 140684 247092 140690
rect 247040 140626 247092 140632
rect 247696 132462 247724 171090
rect 247776 138168 247828 138174
rect 247776 138110 247828 138116
rect 247684 132456 247736 132462
rect 247684 132398 247736 132404
rect 247684 125656 247736 125662
rect 247684 125598 247736 125604
rect 246672 115932 246724 115938
rect 246672 115874 246724 115880
rect 246580 108928 246632 108934
rect 246580 108870 246632 108876
rect 246580 104916 246632 104922
rect 246580 104858 246632 104864
rect 246488 64184 246540 64190
rect 246488 64126 246540 64132
rect 246592 61470 246620 104858
rect 246580 61464 246632 61470
rect 246580 61406 246632 61412
rect 246396 29640 246448 29646
rect 246396 29582 246448 29588
rect 247696 24138 247724 125598
rect 247788 65618 247816 138110
rect 247880 136542 247908 173946
rect 249076 150346 249104 240110
rect 249168 238649 249196 240219
rect 249248 239828 249300 239834
rect 249248 239770 249300 239776
rect 249154 238640 249210 238649
rect 249154 238575 249210 238584
rect 249260 160070 249288 239770
rect 249812 232694 249840 240244
rect 249800 232688 249852 232694
rect 249800 232630 249852 232636
rect 249996 162858 250024 269719
rect 250074 253464 250130 253473
rect 250074 253399 250130 253408
rect 250088 168230 250116 253399
rect 250180 238814 250208 292742
rect 250456 282198 250484 293966
rect 250444 282192 250496 282198
rect 250444 282134 250496 282140
rect 250442 282024 250498 282033
rect 250442 281959 250498 281968
rect 250350 258904 250406 258913
rect 250350 258839 250406 258848
rect 250364 258058 250392 258839
rect 250352 258052 250404 258058
rect 250352 257994 250404 258000
rect 250258 240408 250314 240417
rect 250258 240343 250314 240352
rect 250272 240174 250300 240343
rect 250260 240168 250312 240174
rect 250260 240110 250312 240116
rect 250168 238808 250220 238814
rect 250168 238750 250220 238756
rect 250456 175234 250484 281959
rect 250548 271182 250576 294034
rect 250536 271176 250588 271182
rect 250536 271118 250588 271124
rect 251192 261361 251220 300086
rect 251284 286521 251312 304982
rect 251270 286512 251326 286521
rect 251270 286447 251326 286456
rect 251270 273592 251326 273601
rect 251270 273527 251326 273536
rect 251178 261352 251234 261361
rect 251178 261287 251234 261296
rect 251178 257952 251234 257961
rect 251178 257887 251234 257896
rect 251086 240544 251142 240553
rect 251086 240479 251142 240488
rect 251100 236774 251128 240479
rect 251088 236768 251140 236774
rect 251088 236710 251140 236716
rect 250444 175228 250496 175234
rect 250444 175170 250496 175176
rect 250076 168224 250128 168230
rect 250076 168166 250128 168172
rect 250628 163056 250680 163062
rect 250628 162998 250680 163004
rect 249984 162852 250036 162858
rect 249984 162794 250036 162800
rect 249524 161560 249576 161566
rect 249524 161502 249576 161508
rect 249248 160064 249300 160070
rect 249248 160006 249300 160012
rect 249432 158840 249484 158846
rect 249432 158782 249484 158788
rect 249064 150340 249116 150346
rect 249064 150282 249116 150288
rect 249340 149184 249392 149190
rect 249340 149126 249392 149132
rect 249248 136740 249300 136746
rect 249248 136682 249300 136688
rect 247868 136536 247920 136542
rect 247868 136478 247920 136484
rect 247868 131232 247920 131238
rect 247868 131174 247920 131180
rect 247880 68338 247908 131174
rect 249156 124296 249208 124302
rect 249156 124238 249208 124244
rect 249064 106344 249116 106350
rect 249064 106286 249116 106292
rect 247868 68332 247920 68338
rect 247868 68274 247920 68280
rect 247776 65612 247828 65618
rect 247776 65554 247828 65560
rect 247684 24132 247736 24138
rect 247684 24074 247736 24080
rect 245016 8968 245068 8974
rect 245016 8910 245068 8916
rect 249076 6254 249104 106286
rect 249168 44878 249196 124238
rect 249260 73914 249288 136682
rect 249352 107642 249380 149126
rect 249444 120018 249472 158782
rect 249536 124914 249564 161502
rect 250444 131300 250496 131306
rect 250444 131242 250496 131248
rect 249524 124908 249576 124914
rect 249524 124850 249576 124856
rect 249432 120012 249484 120018
rect 249432 119954 249484 119960
rect 249340 107636 249392 107642
rect 249340 107578 249392 107584
rect 249340 102264 249392 102270
rect 249340 102206 249392 102212
rect 249248 73908 249300 73914
rect 249248 73850 249300 73856
rect 249352 51746 249380 102206
rect 249340 51740 249392 51746
rect 249340 51682 249392 51688
rect 249156 44872 249208 44878
rect 249156 44814 249208 44820
rect 250456 43450 250484 131242
rect 250640 124166 250668 162998
rect 250720 154692 250772 154698
rect 250720 154634 250772 154640
rect 250628 124160 250680 124166
rect 250628 124102 250680 124108
rect 250536 123004 250588 123010
rect 250536 122946 250588 122952
rect 250548 54602 250576 122946
rect 250732 122126 250760 154634
rect 250812 143676 250864 143682
rect 250812 143618 250864 143624
rect 250720 122120 250772 122126
rect 250720 122062 250772 122068
rect 250824 116618 250852 143618
rect 251192 143478 251220 257887
rect 251284 172514 251312 273527
rect 251836 271930 251864 500958
rect 251916 474768 251968 474774
rect 251916 474710 251968 474716
rect 251928 277030 251956 474710
rect 252560 302660 252612 302666
rect 252560 302602 252612 302608
rect 252572 291961 252600 302602
rect 252558 291952 252614 291961
rect 252558 291887 252614 291896
rect 252926 289232 252982 289241
rect 252926 289167 252982 289176
rect 252940 288454 252968 289167
rect 252928 288448 252980 288454
rect 252928 288390 252980 288396
rect 252558 280392 252614 280401
rect 252558 280327 252560 280336
rect 252612 280327 252614 280336
rect 252560 280298 252612 280304
rect 252006 279032 252062 279041
rect 252006 278967 252062 278976
rect 251916 277024 251968 277030
rect 251916 276966 251968 276972
rect 251824 271924 251876 271930
rect 251824 271866 251876 271872
rect 251362 271552 251418 271561
rect 251362 271487 251418 271496
rect 251272 172508 251324 172514
rect 251272 172450 251324 172456
rect 251376 172446 251404 271487
rect 252020 173806 252048 278967
rect 252560 277024 252612 277030
rect 252560 276966 252612 276972
rect 252572 263401 252600 276966
rect 252652 274304 252704 274310
rect 252650 274272 252652 274281
rect 252704 274272 252706 274281
rect 252650 274207 252706 274216
rect 253216 272921 253244 579634
rect 257436 324352 257488 324358
rect 257436 324294 257488 324300
rect 254584 311908 254636 311914
rect 254584 311850 254636 311856
rect 253296 300144 253348 300150
rect 253296 300086 253348 300092
rect 253308 283801 253336 300086
rect 254032 294160 254084 294166
rect 254032 294102 254084 294108
rect 253388 292732 253440 292738
rect 253388 292674 253440 292680
rect 253294 283792 253350 283801
rect 253294 283727 253350 283736
rect 253400 278050 253428 292674
rect 253940 292664 253992 292670
rect 253940 292606 253992 292612
rect 253756 291372 253808 291378
rect 253756 291314 253808 291320
rect 253768 291281 253796 291314
rect 253754 291272 253810 291281
rect 253754 291207 253810 291216
rect 253756 291168 253808 291174
rect 253756 291110 253808 291116
rect 253768 289921 253796 291110
rect 253754 289912 253810 289921
rect 253754 289847 253810 289856
rect 253754 288552 253810 288561
rect 253754 288487 253756 288496
rect 253808 288487 253810 288496
rect 253756 288458 253808 288464
rect 253754 287872 253810 287881
rect 253754 287807 253810 287816
rect 253768 287094 253796 287807
rect 253756 287088 253808 287094
rect 253756 287030 253808 287036
rect 253754 285832 253810 285841
rect 253754 285767 253810 285776
rect 253768 285734 253796 285767
rect 253756 285728 253808 285734
rect 253756 285670 253808 285676
rect 253848 285660 253900 285666
rect 253848 285602 253900 285608
rect 253860 284481 253888 285602
rect 253846 284472 253902 284481
rect 253846 284407 253902 284416
rect 253754 283112 253810 283121
rect 253754 283047 253810 283056
rect 253768 282946 253796 283047
rect 253756 282940 253808 282946
rect 253756 282882 253808 282888
rect 253754 281072 253810 281081
rect 253754 281007 253810 281016
rect 253768 280226 253796 281007
rect 253756 280220 253808 280226
rect 253756 280162 253808 280168
rect 253754 278352 253810 278361
rect 253754 278287 253810 278296
rect 253388 278044 253440 278050
rect 253388 277986 253440 277992
rect 253294 276992 253350 277001
rect 253294 276927 253350 276936
rect 253308 276078 253336 276927
rect 253478 276312 253534 276321
rect 253478 276247 253534 276256
rect 253296 276072 253348 276078
rect 253296 276014 253348 276020
rect 253294 275632 253350 275641
rect 253294 275567 253350 275576
rect 253308 274718 253336 275567
rect 253296 274712 253348 274718
rect 253296 274654 253348 274660
rect 253202 272912 253258 272921
rect 253202 272847 253258 272856
rect 253492 272542 253520 276247
rect 253768 273970 253796 278287
rect 253846 277672 253902 277681
rect 253846 277607 253902 277616
rect 253860 277438 253888 277607
rect 253848 277432 253900 277438
rect 253848 277374 253900 277380
rect 253756 273964 253808 273970
rect 253756 273906 253808 273912
rect 253480 272536 253532 272542
rect 253480 272478 253532 272484
rect 252650 272232 252706 272241
rect 252650 272167 252652 272176
rect 252704 272167 252706 272176
rect 252652 272138 252704 272144
rect 252652 271924 252704 271930
rect 252652 271866 252704 271872
rect 252664 268841 252692 271866
rect 252650 268832 252706 268841
rect 252650 268767 252706 268776
rect 253202 268152 253258 268161
rect 253202 268087 253258 268096
rect 253216 267782 253244 268087
rect 253204 267776 253256 267782
rect 253204 267718 253256 267724
rect 253294 267472 253350 267481
rect 253294 267407 253350 267416
rect 253308 266422 253336 267407
rect 253754 266792 253810 266801
rect 253754 266727 253810 266736
rect 253768 266490 253796 266727
rect 253756 266484 253808 266490
rect 253756 266426 253808 266432
rect 253296 266416 253348 266422
rect 253296 266358 253348 266364
rect 253846 266112 253902 266121
rect 253846 266047 253902 266056
rect 253754 265432 253810 265441
rect 253754 265367 253810 265376
rect 253768 265062 253796 265367
rect 253756 265056 253808 265062
rect 253756 264998 253808 265004
rect 253860 264994 253888 266047
rect 253848 264988 253900 264994
rect 253848 264930 253900 264936
rect 253756 264920 253808 264926
rect 253756 264862 253808 264868
rect 253768 264761 253796 264862
rect 253754 264752 253810 264761
rect 253754 264687 253810 264696
rect 252742 264072 252798 264081
rect 252742 264007 252798 264016
rect 252558 263392 252614 263401
rect 252558 263327 252614 263336
rect 252560 259072 252612 259078
rect 252560 259014 252612 259020
rect 252572 258641 252600 259014
rect 252558 258632 252614 258641
rect 252558 258567 252614 258576
rect 252756 258074 252784 264007
rect 253754 262712 253810 262721
rect 253754 262647 253810 262656
rect 253768 262274 253796 262647
rect 253756 262268 253808 262274
rect 253756 262210 253808 262216
rect 253386 262032 253442 262041
rect 253386 261967 253442 261976
rect 253400 260914 253428 261967
rect 253388 260908 253440 260914
rect 253388 260850 253440 260856
rect 252834 260672 252890 260681
rect 252834 260607 252890 260616
rect 252848 259486 252876 260607
rect 253202 259992 253258 260001
rect 253202 259927 253258 259936
rect 253216 259554 253244 259927
rect 253204 259548 253256 259554
rect 253204 259490 253256 259496
rect 252836 259480 252888 259486
rect 252836 259422 252888 259428
rect 253848 258120 253900 258126
rect 252756 258046 252876 258074
rect 253768 258068 253848 258074
rect 253768 258062 253900 258068
rect 253768 258058 253888 258062
rect 252742 250472 252798 250481
rect 252742 250407 252798 250416
rect 252650 248432 252706 248441
rect 252650 248367 252706 248376
rect 252558 241632 252614 241641
rect 252558 241567 252560 241576
rect 252612 241567 252614 241576
rect 252560 241538 252612 241544
rect 252664 225622 252692 248367
rect 252756 239426 252784 250407
rect 252744 239420 252796 239426
rect 252744 239362 252796 239368
rect 252848 235414 252876 258046
rect 253756 258052 253888 258058
rect 253808 258046 253888 258052
rect 253756 257994 253808 258000
rect 253020 257576 253072 257582
rect 253020 257518 253072 257524
rect 253032 257281 253060 257518
rect 253018 257272 253074 257281
rect 253018 257207 253074 257216
rect 253112 256692 253164 256698
rect 253112 256634 253164 256640
rect 253124 255921 253152 256634
rect 253756 256624 253808 256630
rect 253754 256592 253756 256601
rect 253808 256592 253810 256601
rect 253754 256527 253810 256536
rect 253110 255912 253166 255921
rect 253110 255847 253166 255856
rect 253754 255232 253810 255241
rect 253754 255167 253810 255176
rect 253018 254552 253074 254561
rect 253018 254487 253074 254496
rect 253032 254046 253060 254487
rect 253020 254040 253072 254046
rect 253020 253982 253072 253988
rect 253768 253978 253796 255167
rect 253756 253972 253808 253978
rect 253756 253914 253808 253920
rect 253846 253192 253902 253201
rect 253846 253127 253902 253136
rect 253860 252618 253888 253127
rect 253848 252612 253900 252618
rect 253848 252554 253900 252560
rect 253756 252544 253808 252550
rect 253754 252512 253756 252521
rect 253808 252512 253810 252521
rect 253754 252447 253810 252456
rect 253478 251832 253534 251841
rect 253478 251767 253534 251776
rect 253386 251152 253442 251161
rect 253386 251087 253442 251096
rect 253400 250034 253428 251087
rect 253492 250510 253520 251767
rect 253480 250504 253532 250510
rect 253480 250446 253532 250452
rect 253388 250028 253440 250034
rect 253388 249970 253440 249976
rect 253754 249792 253810 249801
rect 253754 249727 253756 249736
rect 253808 249727 253810 249736
rect 253756 249698 253808 249704
rect 253754 249112 253810 249121
rect 253754 249047 253810 249056
rect 253768 248470 253796 249047
rect 253756 248464 253808 248470
rect 253756 248406 253808 248412
rect 253848 248396 253900 248402
rect 253848 248338 253900 248344
rect 253860 247761 253888 248338
rect 253846 247752 253902 247761
rect 253846 247687 253902 247696
rect 253756 247104 253808 247110
rect 253754 247072 253756 247081
rect 253808 247072 253810 247081
rect 253754 247007 253810 247016
rect 253754 245712 253810 245721
rect 253754 245647 253756 245656
rect 253808 245647 253810 245656
rect 253756 245618 253808 245624
rect 253848 245608 253900 245614
rect 253848 245550 253900 245556
rect 253860 245041 253888 245550
rect 253846 245032 253902 245041
rect 253846 244967 253902 244976
rect 253754 244352 253810 244361
rect 253754 244287 253756 244296
rect 253808 244287 253810 244296
rect 253756 244258 253808 244264
rect 253388 244248 253440 244254
rect 253388 244190 253440 244196
rect 253400 243001 253428 244190
rect 253754 243672 253810 243681
rect 253754 243607 253810 243616
rect 253768 243030 253796 243607
rect 253756 243024 253808 243030
rect 253386 242992 253442 243001
rect 253756 242966 253808 242972
rect 253386 242927 253442 242936
rect 253756 242888 253808 242894
rect 253756 242830 253808 242836
rect 253768 242321 253796 242830
rect 253754 242312 253810 242321
rect 253754 242247 253810 242256
rect 253754 240272 253810 240281
rect 253754 240207 253810 240216
rect 253768 240174 253796 240207
rect 253756 240168 253808 240174
rect 253756 240110 253808 240116
rect 252836 235408 252888 235414
rect 252836 235350 252888 235356
rect 253848 233980 253900 233986
rect 253848 233922 253900 233928
rect 252652 225616 252704 225622
rect 252652 225558 252704 225564
rect 252008 173800 252060 173806
rect 252008 173742 252060 173748
rect 251364 172440 251416 172446
rect 251364 172382 251416 172388
rect 251824 171216 251876 171222
rect 251824 171158 251876 171164
rect 251180 143472 251232 143478
rect 251180 143414 251232 143420
rect 251836 141506 251864 171158
rect 253204 156120 253256 156126
rect 253204 156062 253256 156068
rect 252192 153876 252244 153882
rect 252192 153818 252244 153824
rect 252100 145036 252152 145042
rect 252100 144978 252152 144984
rect 251824 141500 251876 141506
rect 251824 141442 251876 141448
rect 252008 127084 252060 127090
rect 252008 127026 252060 127032
rect 251916 124364 251968 124370
rect 251916 124306 251968 124312
rect 250812 116612 250864 116618
rect 250812 116554 250864 116560
rect 251824 116068 251876 116074
rect 251824 116010 251876 116016
rect 250628 109064 250680 109070
rect 250628 109006 250680 109012
rect 250640 72486 250668 109006
rect 250628 72480 250680 72486
rect 250628 72422 250680 72428
rect 250536 54596 250588 54602
rect 250536 54538 250588 54544
rect 250444 43444 250496 43450
rect 250444 43386 250496 43392
rect 251836 20058 251864 116010
rect 251928 53174 251956 124306
rect 252020 76566 252048 127026
rect 252112 103494 252140 144978
rect 252204 117298 252232 153818
rect 253216 123554 253244 156062
rect 253388 135380 253440 135386
rect 253388 135322 253440 135328
rect 253296 134020 253348 134026
rect 253296 133962 253348 133968
rect 253204 123548 253256 123554
rect 253204 123490 253256 123496
rect 253204 121576 253256 121582
rect 253204 121518 253256 121524
rect 252192 117292 252244 117298
rect 252192 117234 252244 117240
rect 252100 103488 252152 103494
rect 252100 103430 252152 103436
rect 252100 99476 252152 99482
rect 252100 99418 252152 99424
rect 252008 76560 252060 76566
rect 252008 76502 252060 76508
rect 252112 62830 252140 99418
rect 252100 62824 252152 62830
rect 252100 62766 252152 62772
rect 251916 53168 251968 53174
rect 251916 53110 251968 53116
rect 253216 21486 253244 121518
rect 253308 36582 253336 133962
rect 253400 75274 253428 135322
rect 253860 93838 253888 233922
rect 253952 150278 253980 292606
rect 254044 168298 254072 294102
rect 254122 290592 254178 290601
rect 254122 290527 254178 290536
rect 254136 239834 254164 290527
rect 254596 274310 254624 311850
rect 255504 294704 255556 294710
rect 255504 294646 255556 294652
rect 255412 291304 255464 291310
rect 255412 291246 255464 291252
rect 254584 274304 254636 274310
rect 254584 274246 254636 274252
rect 254216 272196 254268 272202
rect 254216 272138 254268 272144
rect 254124 239828 254176 239834
rect 254124 239770 254176 239776
rect 254228 232626 254256 272138
rect 254216 232620 254268 232626
rect 254216 232562 254268 232568
rect 254676 173188 254728 173194
rect 254676 173130 254728 173136
rect 254032 168292 254084 168298
rect 254032 168234 254084 168240
rect 253940 150272 253992 150278
rect 253940 150214 253992 150220
rect 254688 135250 254716 173130
rect 255424 165578 255452 291246
rect 255516 259078 255544 294646
rect 257342 292768 257398 292777
rect 257342 292703 257398 292712
rect 256700 291236 256752 291242
rect 256700 291178 256752 291184
rect 255596 280356 255648 280362
rect 255596 280298 255648 280304
rect 255504 259072 255556 259078
rect 255504 259014 255556 259020
rect 255504 241596 255556 241602
rect 255504 241538 255556 241544
rect 255516 233986 255544 241538
rect 255504 233980 255556 233986
rect 255504 233922 255556 233928
rect 255412 165572 255464 165578
rect 255412 165514 255464 165520
rect 254768 158024 254820 158030
rect 254768 157966 254820 157972
rect 254676 135244 254728 135250
rect 254676 135186 254728 135192
rect 254584 134088 254636 134094
rect 254584 134030 254636 134036
rect 253848 93832 253900 93838
rect 253848 93774 253900 93780
rect 253388 75268 253440 75274
rect 253388 75210 253440 75216
rect 253296 36576 253348 36582
rect 253296 36518 253348 36524
rect 253204 21480 253256 21486
rect 253204 21422 253256 21428
rect 251824 20052 251876 20058
rect 251824 19994 251876 20000
rect 254596 9042 254624 134030
rect 254780 126954 254808 157966
rect 254860 150544 254912 150550
rect 254860 150486 254912 150492
rect 254768 126948 254820 126954
rect 254768 126890 254820 126896
rect 254676 122936 254728 122942
rect 254676 122878 254728 122884
rect 254688 38010 254716 122878
rect 254768 118720 254820 118726
rect 254768 118662 254820 118668
rect 254780 49094 254808 118662
rect 254872 110362 254900 150486
rect 255608 142118 255636 280298
rect 256056 174072 256108 174078
rect 256056 174014 256108 174020
rect 255964 160268 256016 160274
rect 255964 160210 256016 160216
rect 255596 142112 255648 142118
rect 255596 142054 255648 142060
rect 255976 120086 256004 160210
rect 256068 136610 256096 174014
rect 256332 140820 256384 140826
rect 256332 140762 256384 140768
rect 256056 136604 256108 136610
rect 256056 136546 256108 136552
rect 255964 120080 256016 120086
rect 255964 120022 256016 120028
rect 256148 118788 256200 118794
rect 256148 118730 256200 118736
rect 256056 113348 256108 113354
rect 256056 113290 256108 113296
rect 254860 110356 254912 110362
rect 254860 110298 254912 110304
rect 255964 104984 256016 104990
rect 255964 104926 256016 104932
rect 254860 100904 254912 100910
rect 254860 100846 254912 100852
rect 254872 60042 254900 100846
rect 254860 60036 254912 60042
rect 254860 59978 254912 59984
rect 254768 49088 254820 49094
rect 254768 49030 254820 49036
rect 254676 38004 254728 38010
rect 254676 37946 254728 37952
rect 255976 14482 256004 104926
rect 256068 26926 256096 113290
rect 256160 50454 256188 118730
rect 256240 116136 256292 116142
rect 256240 116078 256292 116084
rect 256252 66910 256280 116078
rect 256344 105602 256372 140762
rect 256712 140758 256740 291178
rect 256792 259548 256844 259554
rect 256792 259490 256844 259496
rect 256804 157282 256832 259490
rect 256884 254040 256936 254046
rect 256884 253982 256936 253988
rect 256896 240417 256924 253982
rect 256882 240408 256938 240417
rect 256882 240343 256938 240352
rect 257356 206990 257384 292703
rect 257448 257582 257476 324294
rect 258172 295724 258224 295730
rect 258172 295666 258224 295672
rect 258080 293276 258132 293282
rect 258080 293218 258132 293224
rect 257436 257576 257488 257582
rect 257436 257518 257488 257524
rect 257344 206984 257396 206990
rect 257344 206926 257396 206932
rect 258092 169726 258120 293218
rect 258184 235249 258212 295666
rect 258736 239970 258764 699654
rect 260104 698964 260156 698970
rect 260104 698906 260156 698912
rect 259552 298512 259604 298518
rect 259552 298454 259604 298460
rect 259460 291372 259512 291378
rect 259460 291314 259512 291320
rect 258724 239964 258776 239970
rect 258724 239906 258776 239912
rect 258170 235240 258226 235249
rect 258170 235175 258226 235184
rect 258816 171556 258868 171562
rect 258816 171498 258868 171504
rect 258080 169720 258132 169726
rect 258080 169662 258132 169668
rect 257436 164348 257488 164354
rect 257436 164290 257488 164296
rect 256792 157276 256844 157282
rect 256792 157218 256844 157224
rect 256700 140752 256752 140758
rect 256700 140694 256752 140700
rect 257344 139460 257396 139466
rect 257344 139402 257396 139408
rect 256332 105596 256384 105602
rect 256332 105538 256384 105544
rect 256240 66904 256292 66910
rect 256240 66846 256292 66852
rect 256148 50448 256200 50454
rect 256148 50390 256200 50396
rect 256056 26920 256108 26926
rect 256056 26862 256108 26868
rect 257356 15978 257384 139402
rect 257448 129062 257476 164290
rect 258724 150612 258776 150618
rect 258724 150554 258776 150560
rect 257436 129056 257488 129062
rect 257436 128998 257488 129004
rect 257528 128444 257580 128450
rect 257528 128386 257580 128392
rect 257436 117428 257488 117434
rect 257436 117370 257488 117376
rect 257448 31074 257476 117370
rect 257540 42090 257568 128386
rect 257620 125724 257672 125730
rect 257620 125666 257672 125672
rect 257632 58750 257660 125666
rect 258736 112470 258764 150554
rect 258828 133890 258856 171498
rect 258908 155576 258960 155582
rect 258908 155518 258960 155524
rect 258816 133884 258868 133890
rect 258816 133826 258868 133832
rect 258920 121446 258948 155518
rect 259000 147756 259052 147762
rect 259000 147698 259052 147704
rect 258908 121440 258960 121446
rect 258908 121382 258960 121388
rect 258816 120216 258868 120222
rect 258816 120158 258868 120164
rect 258724 112464 258776 112470
rect 258724 112406 258776 112412
rect 258724 105052 258776 105058
rect 258724 104994 258776 105000
rect 257620 58744 257672 58750
rect 257620 58686 257672 58692
rect 257528 42084 257580 42090
rect 257528 42026 257580 42032
rect 257436 31068 257488 31074
rect 257436 31010 257488 31016
rect 257344 15972 257396 15978
rect 257344 15914 257396 15920
rect 255964 14476 256016 14482
rect 255964 14418 256016 14424
rect 258736 13122 258764 104994
rect 258828 29714 258856 120158
rect 258908 110628 258960 110634
rect 258908 110570 258960 110576
rect 258816 29708 258868 29714
rect 258816 29650 258868 29656
rect 258920 25634 258948 110570
rect 259012 106282 259040 147698
rect 259472 143546 259500 291314
rect 259564 157350 259592 298454
rect 259644 250028 259696 250034
rect 259644 249970 259696 249976
rect 259656 202842 259684 249970
rect 260116 243030 260144 698906
rect 264244 696244 264296 696250
rect 264244 696186 264296 696192
rect 262864 643136 262916 643142
rect 262864 643078 262916 643084
rect 260840 298444 260892 298450
rect 260840 298386 260892 298392
rect 260104 243024 260156 243030
rect 260104 242966 260156 242972
rect 259644 202836 259696 202842
rect 259644 202778 259696 202784
rect 260288 168564 260340 168570
rect 260288 168506 260340 168512
rect 260196 162172 260248 162178
rect 260196 162114 260248 162120
rect 259552 157344 259604 157350
rect 259552 157286 259604 157292
rect 259460 143540 259512 143546
rect 259460 143482 259512 143488
rect 260104 135516 260156 135522
rect 260104 135458 260156 135464
rect 259092 106480 259144 106486
rect 259092 106422 259144 106428
rect 259000 106276 259052 106282
rect 259000 106218 259052 106224
rect 259104 75206 259132 106422
rect 259092 75200 259144 75206
rect 259092 75142 259144 75148
rect 258908 25628 258960 25634
rect 258908 25570 258960 25576
rect 260116 22778 260144 135458
rect 260208 122806 260236 162114
rect 260300 131034 260328 168506
rect 260852 158710 260880 298386
rect 262312 296812 262364 296818
rect 262312 296754 262364 296760
rect 260932 295588 260984 295594
rect 260932 295530 260984 295536
rect 260944 168366 260972 295530
rect 262220 292868 262272 292874
rect 262220 292810 262272 292816
rect 260932 168360 260984 168366
rect 260932 168302 260984 168308
rect 261390 166832 261446 166841
rect 261390 166767 261446 166776
rect 261404 164898 261432 166767
rect 261484 165708 261536 165714
rect 261484 165650 261536 165656
rect 261392 164892 261444 164898
rect 261392 164834 261444 164840
rect 260840 158704 260892 158710
rect 260840 158646 260892 158652
rect 261496 144129 261524 165650
rect 261666 157312 261722 157321
rect 261666 157247 261722 157256
rect 261680 155582 261708 157247
rect 261668 155576 261720 155582
rect 261668 155518 261720 155524
rect 262232 153202 262260 292810
rect 262324 161430 262352 296754
rect 262402 268424 262458 268433
rect 262402 268359 262458 268368
rect 262312 161424 262364 161430
rect 262312 161366 262364 161372
rect 262220 153196 262272 153202
rect 262220 153138 262272 153144
rect 261760 151836 261812 151842
rect 261760 151778 261812 151784
rect 261574 146160 261630 146169
rect 261574 146095 261630 146104
rect 261588 145586 261616 146095
rect 261576 145580 261628 145586
rect 261576 145522 261628 145528
rect 261482 144120 261538 144129
rect 261482 144055 261538 144064
rect 260380 142384 260432 142390
rect 260380 142326 260432 142332
rect 260288 131028 260340 131034
rect 260288 130970 260340 130976
rect 260196 122800 260248 122806
rect 260196 122742 260248 122748
rect 260288 111988 260340 111994
rect 260288 111930 260340 111936
rect 260196 107772 260248 107778
rect 260196 107714 260248 107720
rect 260104 22772 260156 22778
rect 260104 22714 260156 22720
rect 258724 13116 258776 13122
rect 258724 13058 258776 13064
rect 254584 9036 254636 9042
rect 254584 8978 254636 8984
rect 260208 7614 260236 107714
rect 260300 64258 260328 111930
rect 260392 100706 260420 142326
rect 260470 140176 260526 140185
rect 260470 140111 260526 140120
rect 260484 139777 260512 140111
rect 260470 139768 260526 139777
rect 260470 139703 260526 139712
rect 261484 135448 261536 135454
rect 261484 135390 261536 135396
rect 260380 100700 260432 100706
rect 260380 100642 260432 100648
rect 260472 99544 260524 99550
rect 260472 99486 260524 99492
rect 260484 65550 260512 99486
rect 260472 65544 260524 65550
rect 260472 65486 260524 65492
rect 260288 64252 260340 64258
rect 260288 64194 260340 64200
rect 261496 28354 261524 135390
rect 261666 119912 261722 119921
rect 261666 119847 261722 119856
rect 261576 110560 261628 110566
rect 261576 110502 261628 110508
rect 261484 28348 261536 28354
rect 261484 28290 261536 28296
rect 261588 24206 261616 110502
rect 261680 35290 261708 119847
rect 261772 110430 261800 151778
rect 261852 144900 261904 144906
rect 261852 144842 261904 144848
rect 261864 111790 261892 144842
rect 262416 137970 262444 268359
rect 262876 240009 262904 643078
rect 263692 298376 263744 298382
rect 263692 298318 263744 298324
rect 263600 278044 263652 278050
rect 263600 277986 263652 277992
rect 262862 240000 262918 240009
rect 262862 239935 262918 239944
rect 262956 167136 263008 167142
rect 262956 167078 263008 167084
rect 262404 137964 262456 137970
rect 262404 137906 262456 137912
rect 262864 132660 262916 132666
rect 262864 132602 262916 132608
rect 261852 111784 261904 111790
rect 261852 111726 261904 111732
rect 261760 110424 261812 110430
rect 261760 110366 261812 110372
rect 261852 109132 261904 109138
rect 261852 109074 261904 109080
rect 261864 69698 261892 109074
rect 261852 69692 261904 69698
rect 261852 69634 261904 69640
rect 262876 39438 262904 132602
rect 262968 128314 262996 167078
rect 263048 158908 263100 158914
rect 263048 158850 263100 158856
rect 262956 128308 263008 128314
rect 262956 128250 263008 128256
rect 263060 118658 263088 158850
rect 263140 149252 263192 149258
rect 263140 149194 263192 149200
rect 263048 118652 263100 118658
rect 263048 118594 263100 118600
rect 262956 117496 263008 117502
rect 262956 117438 263008 117444
rect 262968 54534 262996 117438
rect 263152 109002 263180 149194
rect 263612 147626 263640 277986
rect 263704 171086 263732 298318
rect 263784 247104 263836 247110
rect 263784 247046 263836 247052
rect 263692 171080 263744 171086
rect 263692 171022 263744 171028
rect 263600 147620 263652 147626
rect 263600 147562 263652 147568
rect 263796 144838 263824 247046
rect 264256 245614 264284 696186
rect 267004 524476 267056 524482
rect 267004 524418 267056 524424
rect 265072 296880 265124 296886
rect 265072 296822 265124 296828
rect 264980 295656 265032 295662
rect 264980 295598 265032 295604
rect 264244 245608 264296 245614
rect 264244 245550 264296 245556
rect 264992 190454 265020 295598
rect 265084 235346 265112 296822
rect 267016 249762 267044 524418
rect 267096 297016 267148 297022
rect 267096 296958 267148 296964
rect 267004 249756 267056 249762
rect 267004 249698 267056 249704
rect 267004 238128 267056 238134
rect 267004 238070 267056 238076
rect 265072 235340 265124 235346
rect 265072 235282 265124 235288
rect 264992 190426 265388 190454
rect 265360 176654 265388 190426
rect 265268 176626 265388 176654
rect 265268 173874 265296 176626
rect 265806 175400 265862 175409
rect 265806 175335 265862 175344
rect 265820 175302 265848 175335
rect 265808 175296 265860 175302
rect 265808 175238 265860 175244
rect 265346 174992 265402 175001
rect 265346 174927 265402 174936
rect 265360 174078 265388 174927
rect 265806 174584 265862 174593
rect 265806 174519 265862 174528
rect 265622 174176 265678 174185
rect 265622 174111 265678 174120
rect 265348 174072 265400 174078
rect 265348 174014 265400 174020
rect 265636 173942 265664 174111
rect 265820 174010 265848 174519
rect 265898 174040 265954 174049
rect 265808 174004 265860 174010
rect 265898 173975 265954 173984
rect 265808 173946 265860 173952
rect 265624 173936 265676 173942
rect 265624 173878 265676 173884
rect 265256 173868 265308 173874
rect 265256 173810 265308 173816
rect 265714 173224 265770 173233
rect 265912 173194 265940 173975
rect 265714 173159 265770 173168
rect 265900 173188 265952 173194
rect 265346 172000 265402 172009
rect 265346 171935 265402 171944
rect 265360 171562 265388 171935
rect 265348 171556 265400 171562
rect 265348 171498 265400 171504
rect 265346 170640 265402 170649
rect 265346 170575 265402 170584
rect 264242 170232 264298 170241
rect 264242 170167 264298 170176
rect 263784 144832 263836 144838
rect 263784 144774 263836 144780
rect 264256 131102 264284 170167
rect 265360 169794 265388 170575
rect 265728 170406 265756 173159
rect 265900 173130 265952 173136
rect 265898 172816 265954 172825
rect 265898 172751 265954 172760
rect 265912 172650 265940 172751
rect 265900 172644 265952 172650
rect 265900 172586 265952 172592
rect 265808 172576 265860 172582
rect 265806 172544 265808 172553
rect 265860 172544 265862 172553
rect 265806 172479 265862 172488
rect 265806 171592 265862 171601
rect 265806 171527 265862 171536
rect 265820 171154 265848 171527
rect 265900 171216 265952 171222
rect 265898 171184 265900 171193
rect 265952 171184 265954 171193
rect 265808 171148 265860 171154
rect 265898 171119 265954 171128
rect 265808 171090 265860 171096
rect 265716 170400 265768 170406
rect 265716 170342 265768 170348
rect 265622 169824 265678 169833
rect 265348 169788 265400 169794
rect 265622 169759 265678 169768
rect 265348 169730 265400 169736
rect 265438 169416 265494 169425
rect 265438 169351 265494 169360
rect 265346 169008 265402 169017
rect 265346 168943 265402 168952
rect 264428 168428 264480 168434
rect 264428 168370 264480 168376
rect 264440 168201 264468 168370
rect 264426 168192 264482 168201
rect 264426 168127 264482 168136
rect 265162 167648 265218 167657
rect 265162 167583 265218 167592
rect 265176 167142 265204 167583
rect 265164 167136 265216 167142
rect 265164 167078 265216 167084
rect 265360 166326 265388 168943
rect 265452 167686 265480 169351
rect 265636 168570 265664 169759
rect 265806 168600 265862 168609
rect 265624 168564 265676 168570
rect 265806 168535 265862 168544
rect 265624 168506 265676 168512
rect 265820 168502 265848 168535
rect 265808 168496 265860 168502
rect 265808 168438 265860 168444
rect 265440 167680 265492 167686
rect 265440 167622 265492 167628
rect 265806 167240 265862 167249
rect 265806 167175 265862 167184
rect 265820 167074 265848 167175
rect 265808 167068 265860 167074
rect 265808 167010 265860 167016
rect 265990 166424 266046 166433
rect 265990 166359 266046 166368
rect 265348 166320 265400 166326
rect 265348 166262 265400 166268
rect 265714 166016 265770 166025
rect 265714 165951 265770 165960
rect 265728 165646 265756 165951
rect 265806 165744 265862 165753
rect 265806 165679 265808 165688
rect 265860 165679 265862 165688
rect 265808 165650 265860 165656
rect 265716 165640 265768 165646
rect 265716 165582 265768 165588
rect 265438 165064 265494 165073
rect 265438 164999 265494 165008
rect 265452 164286 265480 164999
rect 265714 164656 265770 164665
rect 265714 164591 265770 164600
rect 265440 164280 265492 164286
rect 265440 164222 265492 164228
rect 265530 163432 265586 163441
rect 265530 163367 265586 163376
rect 265544 163062 265572 163367
rect 265532 163056 265584 163062
rect 265346 163024 265402 163033
rect 265532 162998 265584 163004
rect 265346 162959 265348 162968
rect 265400 162959 265402 162968
rect 265348 162930 265400 162936
rect 265346 162072 265402 162081
rect 265346 162007 265402 162016
rect 265360 161566 265388 162007
rect 265348 161560 265400 161566
rect 265348 161502 265400 161508
rect 265346 160848 265402 160857
rect 265346 160783 265402 160792
rect 265360 160206 265388 160783
rect 265622 160440 265678 160449
rect 265622 160375 265678 160384
rect 265636 160274 265664 160375
rect 265624 160268 265676 160274
rect 265624 160210 265676 160216
rect 265348 160200 265400 160206
rect 265348 160142 265400 160148
rect 265346 159488 265402 159497
rect 265346 159423 265402 159432
rect 265360 158846 265388 159423
rect 265622 159080 265678 159089
rect 265622 159015 265678 159024
rect 265636 158914 265664 159015
rect 265624 158908 265676 158914
rect 265624 158850 265676 158856
rect 265348 158840 265400 158846
rect 265348 158782 265400 158788
rect 265622 158264 265678 158273
rect 265622 158199 265678 158208
rect 265254 157856 265310 157865
rect 265254 157791 265310 157800
rect 265268 153882 265296 157791
rect 265636 157486 265664 158199
rect 265624 157480 265676 157486
rect 265530 157448 265586 157457
rect 265624 157422 265676 157428
rect 265530 157383 265532 157392
rect 265584 157383 265586 157392
rect 265532 157354 265584 157360
rect 265728 157334 265756 164591
rect 265808 164348 265860 164354
rect 265808 164290 265860 164296
rect 265820 164257 265848 164290
rect 265806 164248 265862 164257
rect 265806 164183 265862 164192
rect 265898 163840 265954 163849
rect 265898 163775 265954 163784
rect 265912 162926 265940 163775
rect 265900 162920 265952 162926
rect 265806 162888 265862 162897
rect 265900 162862 265952 162868
rect 265806 162823 265862 162832
rect 265820 162178 265848 162823
rect 265808 162172 265860 162178
rect 265808 162114 265860 162120
rect 265806 161664 265862 161673
rect 265806 161599 265862 161608
rect 265820 161498 265848 161599
rect 265808 161492 265860 161498
rect 265808 161434 265860 161440
rect 265806 160168 265862 160177
rect 265806 160103 265808 160112
rect 265860 160103 265862 160112
rect 265808 160074 265860 160080
rect 265806 158808 265862 158817
rect 265806 158743 265808 158752
rect 265860 158743 265862 158752
rect 265808 158714 265860 158720
rect 266004 158030 266032 166359
rect 265992 158024 266044 158030
rect 265992 157966 266044 157972
rect 265636 157306 265756 157334
rect 265530 156496 265586 156505
rect 265530 156431 265586 156440
rect 265544 156058 265572 156431
rect 265532 156052 265584 156058
rect 265532 155994 265584 156000
rect 265256 153876 265308 153882
rect 265256 153818 265308 153824
rect 264426 152144 264482 152153
rect 264426 152079 264482 152088
rect 264336 142384 264388 142390
rect 264336 142326 264388 142332
rect 264348 141953 264376 142326
rect 264334 141944 264390 141953
rect 264334 141879 264390 141888
rect 264244 131096 264296 131102
rect 264244 131038 264296 131044
rect 264334 123856 264390 123865
rect 264334 123791 264390 123800
rect 263140 108996 263192 109002
rect 263140 108938 263192 108944
rect 263048 107704 263100 107710
rect 263048 107646 263100 107652
rect 263060 57254 263088 107646
rect 264242 107536 264298 107545
rect 264242 107471 264298 107480
rect 263140 106412 263192 106418
rect 263140 106354 263192 106360
rect 263152 73846 263180 106354
rect 263140 73840 263192 73846
rect 263140 73782 263192 73788
rect 263048 57248 263100 57254
rect 263048 57190 263100 57196
rect 262956 54528 263008 54534
rect 262956 54470 263008 54476
rect 262864 39432 262916 39438
rect 262864 39374 262916 39380
rect 261668 35284 261720 35290
rect 261668 35226 261720 35232
rect 261576 24200 261628 24206
rect 261576 24142 261628 24148
rect 264256 18698 264284 107471
rect 264348 42158 264376 123791
rect 264440 115258 264468 152079
rect 265346 150104 265402 150113
rect 265346 150039 265402 150048
rect 265360 149258 265388 150039
rect 265348 149252 265400 149258
rect 265348 149194 265400 149200
rect 265438 148744 265494 148753
rect 265438 148679 265494 148688
rect 265162 148336 265218 148345
rect 265162 148271 265218 148280
rect 265176 146946 265204 148271
rect 265452 147694 265480 148679
rect 265440 147688 265492 147694
rect 265440 147630 265492 147636
rect 265530 147112 265586 147121
rect 265530 147047 265586 147056
rect 265164 146940 265216 146946
rect 265164 146882 265216 146888
rect 265544 146334 265572 147047
rect 265532 146328 265584 146334
rect 265532 146270 265584 146276
rect 264518 145752 264574 145761
rect 264518 145687 264574 145696
rect 264532 120766 264560 145687
rect 265532 145036 265584 145042
rect 265532 144978 265584 144984
rect 265544 144945 265572 144978
rect 265530 144936 265586 144945
rect 265530 144871 265586 144880
rect 265438 144528 265494 144537
rect 265438 144463 265494 144472
rect 265452 143682 265480 144463
rect 265440 143676 265492 143682
rect 265440 143618 265492 143624
rect 265636 142866 265664 157306
rect 265898 156904 265954 156913
rect 265898 156839 265954 156848
rect 265912 156126 265940 156839
rect 265900 156120 265952 156126
rect 265806 156088 265862 156097
rect 265900 156062 265952 156068
rect 265806 156023 265862 156032
rect 265820 155990 265848 156023
rect 265808 155984 265860 155990
rect 265808 155926 265860 155932
rect 265806 155680 265862 155689
rect 265806 155615 265862 155624
rect 265714 155272 265770 155281
rect 265714 155207 265770 155216
rect 265728 154630 265756 155207
rect 265820 154698 265848 155615
rect 265990 154728 266046 154737
rect 265808 154692 265860 154698
rect 265990 154663 266046 154672
rect 265808 154634 265860 154640
rect 265716 154624 265768 154630
rect 265716 154566 265768 154572
rect 265898 153912 265954 153921
rect 265898 153847 265954 153856
rect 265806 153504 265862 153513
rect 265806 153439 265862 153448
rect 265820 153270 265848 153439
rect 265912 153338 265940 153847
rect 265900 153332 265952 153338
rect 265900 153274 265952 153280
rect 265808 153264 265860 153270
rect 265808 153206 265860 153212
rect 265898 153232 265954 153241
rect 265898 153167 265954 153176
rect 265714 152688 265770 152697
rect 265714 152623 265770 152632
rect 265728 151978 265756 152623
rect 265716 151972 265768 151978
rect 265716 151914 265768 151920
rect 265806 151872 265862 151881
rect 265806 151807 265808 151816
rect 265860 151807 265862 151816
rect 265808 151778 265860 151784
rect 265912 151042 265940 153167
rect 266004 152522 266032 154663
rect 266082 154592 266138 154601
rect 266082 154527 266138 154536
rect 265992 152516 266044 152522
rect 265992 152458 266044 152464
rect 265990 151328 266046 151337
rect 265990 151263 266046 151272
rect 265728 151014 265940 151042
rect 265728 144906 265756 151014
rect 265898 150920 265954 150929
rect 265898 150855 265954 150864
rect 265912 150618 265940 150855
rect 265900 150612 265952 150618
rect 265900 150554 265952 150560
rect 266004 150550 266032 151263
rect 265992 150544 266044 150550
rect 265806 150512 265862 150521
rect 265992 150486 266044 150492
rect 265806 150447 265808 150456
rect 265860 150447 265862 150456
rect 265808 150418 265860 150424
rect 265898 149696 265954 149705
rect 265898 149631 265954 149640
rect 265806 149288 265862 149297
rect 265806 149223 265862 149232
rect 265820 149190 265848 149223
rect 265808 149184 265860 149190
rect 265808 149126 265860 149132
rect 265912 149122 265940 149631
rect 265900 149116 265952 149122
rect 265900 149058 265952 149064
rect 266096 148374 266124 154527
rect 266084 148368 266136 148374
rect 266084 148310 266136 148316
rect 265806 147928 265862 147937
rect 265806 147863 265862 147872
rect 265820 147762 265848 147863
rect 265808 147756 265860 147762
rect 265808 147698 265860 147704
rect 265806 146704 265862 146713
rect 265806 146639 265862 146648
rect 265820 146402 265848 146639
rect 266082 146568 266138 146577
rect 266082 146503 266138 146512
rect 265808 146396 265860 146402
rect 265808 146338 265860 146344
rect 265806 145344 265862 145353
rect 265806 145279 265862 145288
rect 265820 145110 265848 145279
rect 265808 145104 265860 145110
rect 265808 145046 265860 145052
rect 265716 144900 265768 144906
rect 265716 144842 265768 144848
rect 265806 143984 265862 143993
rect 265806 143919 265862 143928
rect 265820 143614 265848 143919
rect 265808 143608 265860 143614
rect 265808 143550 265860 143556
rect 265898 143576 265954 143585
rect 265898 143511 265954 143520
rect 265714 143168 265770 143177
rect 265714 143103 265770 143112
rect 265624 142860 265676 142866
rect 265624 142802 265676 142808
rect 265346 142760 265402 142769
rect 265346 142695 265402 142704
rect 264610 142352 264666 142361
rect 265360 142322 265388 142695
rect 264610 142287 264666 142296
rect 265348 142316 265400 142322
rect 264520 120760 264572 120766
rect 264520 120702 264572 120708
rect 264520 116136 264572 116142
rect 264520 116078 264572 116084
rect 264532 115977 264560 116078
rect 264518 115968 264574 115977
rect 264518 115903 264574 115912
rect 264428 115252 264480 115258
rect 264428 115194 264480 115200
rect 264518 110120 264574 110129
rect 264518 110055 264574 110064
rect 264426 104544 264482 104553
rect 264426 104479 264482 104488
rect 264336 42152 264388 42158
rect 264336 42094 264388 42100
rect 264440 26994 264468 104479
rect 264532 66978 264560 110055
rect 264624 106962 264652 142287
rect 265348 142258 265400 142264
rect 265438 139496 265494 139505
rect 265438 139431 265440 139440
rect 265492 139431 265494 139440
rect 265440 139402 265492 139408
rect 265438 138816 265494 138825
rect 265438 138751 265494 138760
rect 265162 138408 265218 138417
rect 265162 138343 265218 138352
rect 265176 138106 265204 138343
rect 265164 138100 265216 138106
rect 265164 138042 265216 138048
rect 265452 138038 265480 138751
rect 265624 138168 265676 138174
rect 265622 138136 265624 138145
rect 265676 138136 265678 138145
rect 265622 138071 265678 138080
rect 265440 138032 265492 138038
rect 265440 137974 265492 137980
rect 265622 137592 265678 137601
rect 265622 137527 265678 137536
rect 265530 136776 265586 136785
rect 265530 136711 265532 136720
rect 265584 136711 265586 136720
rect 265532 136682 265584 136688
rect 265636 136678 265664 137527
rect 265624 136672 265676 136678
rect 265624 136614 265676 136620
rect 265622 136368 265678 136377
rect 265622 136303 265678 136312
rect 265346 135960 265402 135969
rect 265346 135895 265402 135904
rect 265360 135522 265388 135895
rect 265348 135516 265400 135522
rect 265348 135458 265400 135464
rect 265636 135386 265664 136303
rect 265624 135380 265676 135386
rect 265624 135322 265676 135328
rect 265530 134600 265586 134609
rect 265530 134535 265586 134544
rect 265544 134026 265572 134535
rect 265532 134020 265584 134026
rect 265532 133962 265584 133968
rect 265622 132832 265678 132841
rect 265622 132767 265678 132776
rect 265636 132666 265664 132767
rect 265624 132660 265676 132666
rect 265624 132602 265676 132608
rect 265162 131608 265218 131617
rect 265162 131543 265218 131552
rect 265176 131306 265204 131543
rect 265164 131300 265216 131306
rect 265164 131242 265216 131248
rect 265624 131232 265676 131238
rect 265622 131200 265624 131209
rect 265676 131200 265678 131209
rect 265622 131135 265678 131144
rect 265530 130656 265586 130665
rect 265530 130591 265586 130600
rect 265544 128354 265572 130591
rect 265622 129024 265678 129033
rect 265622 128959 265678 128968
rect 265636 128450 265664 128959
rect 265624 128444 265676 128450
rect 265624 128386 265676 128392
rect 265544 128326 265664 128354
rect 265346 127664 265402 127673
rect 265346 127599 265402 127608
rect 265360 127022 265388 127599
rect 265348 127016 265400 127022
rect 265348 126958 265400 126964
rect 265254 126032 265310 126041
rect 265254 125967 265310 125976
rect 265268 125730 265296 125967
rect 265256 125724 265308 125730
rect 265256 125666 265308 125672
rect 265530 124672 265586 124681
rect 265530 124607 265586 124616
rect 265544 124302 265572 124607
rect 265532 124296 265584 124302
rect 265532 124238 265584 124244
rect 265530 123448 265586 123457
rect 265530 123383 265586 123392
rect 265070 123040 265126 123049
rect 265070 122975 265072 122984
rect 265124 122975 265126 122984
rect 265072 122946 265124 122952
rect 265544 122942 265572 123383
rect 265532 122936 265584 122942
rect 265532 122878 265584 122884
rect 265254 119096 265310 119105
rect 265254 119031 265310 119040
rect 265268 118794 265296 119031
rect 265256 118788 265308 118794
rect 265256 118730 265308 118736
rect 265530 118280 265586 118289
rect 265530 118215 265586 118224
rect 265162 117872 265218 117881
rect 265162 117807 265218 117816
rect 265176 117502 265204 117807
rect 265164 117496 265216 117502
rect 265164 117438 265216 117444
rect 265544 117434 265572 118215
rect 265532 117428 265584 117434
rect 265532 117370 265584 117376
rect 265254 114880 265310 114889
rect 265254 114815 265310 114824
rect 265268 114578 265296 114815
rect 265256 114572 265308 114578
rect 265256 114514 265308 114520
rect 265254 113520 265310 113529
rect 265254 113455 265310 113464
rect 265268 113286 265296 113455
rect 265256 113280 265308 113286
rect 265256 113222 265308 113228
rect 265438 113248 265494 113257
rect 265438 113183 265440 113192
rect 265492 113183 265494 113192
rect 265440 113154 265492 113160
rect 265530 112704 265586 112713
rect 265530 112639 265586 112648
rect 265544 111926 265572 112639
rect 265532 111920 265584 111926
rect 265532 111862 265584 111868
rect 265530 111344 265586 111353
rect 265530 111279 265586 111288
rect 265162 110936 265218 110945
rect 265162 110871 265218 110880
rect 265176 110566 265204 110871
rect 265544 110634 265572 111279
rect 265532 110628 265584 110634
rect 265532 110570 265584 110576
rect 265164 110560 265216 110566
rect 265164 110502 265216 110508
rect 265530 109712 265586 109721
rect 265530 109647 265586 109656
rect 265544 109138 265572 109647
rect 265532 109132 265584 109138
rect 265532 109074 265584 109080
rect 265438 108352 265494 108361
rect 265438 108287 265494 108296
rect 265346 107944 265402 107953
rect 265346 107879 265348 107888
rect 265400 107879 265402 107888
rect 265348 107850 265400 107856
rect 265452 107778 265480 108287
rect 265440 107772 265492 107778
rect 265440 107714 265492 107720
rect 265530 107128 265586 107137
rect 265530 107063 265586 107072
rect 264612 106956 264664 106962
rect 264612 106898 264664 106904
rect 265440 106820 265492 106826
rect 265440 106762 265492 106768
rect 265452 104174 265480 106762
rect 265544 106418 265572 107063
rect 265532 106412 265584 106418
rect 265532 106354 265584 106360
rect 265440 104168 265492 104174
rect 265440 104110 265492 104116
rect 265530 101960 265586 101969
rect 265530 101895 265586 101904
rect 265544 100910 265572 101895
rect 265532 100904 265584 100910
rect 265532 100846 265584 100852
rect 265530 99512 265586 99521
rect 265530 99447 265586 99456
rect 265544 99414 265572 99447
rect 265532 99408 265584 99414
rect 265532 99350 265584 99356
rect 265440 98048 265492 98054
rect 265438 98016 265440 98025
rect 265492 98016 265494 98025
rect 265438 97951 265494 97960
rect 265162 97200 265218 97209
rect 265162 97135 265218 97144
rect 265176 96762 265204 97135
rect 265164 96756 265216 96762
rect 265164 96698 265216 96704
rect 264520 66972 264572 66978
rect 264520 66914 264572 66920
rect 265636 33794 265664 128326
rect 265728 123486 265756 143103
rect 265806 140992 265862 141001
rect 265806 140927 265862 140936
rect 265820 140826 265848 140927
rect 265808 140820 265860 140826
rect 265808 140762 265860 140768
rect 265912 138014 265940 143511
rect 266096 141438 266124 146503
rect 266084 141432 266136 141438
rect 265990 141400 266046 141409
rect 266084 141374 266136 141380
rect 265990 141335 266046 141344
rect 265820 137986 265940 138014
rect 265716 123480 265768 123486
rect 265716 123422 265768 123428
rect 265714 119504 265770 119513
rect 265714 119439 265770 119448
rect 265728 118726 265756 119439
rect 265716 118720 265768 118726
rect 265716 118662 265768 118668
rect 265714 117464 265770 117473
rect 265714 117399 265770 117408
rect 265728 117366 265756 117399
rect 265716 117360 265768 117366
rect 265716 117302 265768 117308
rect 265714 113928 265770 113937
rect 265714 113863 265770 113872
rect 265728 113354 265756 113863
rect 265716 113348 265768 113354
rect 265716 113290 265768 113296
rect 265714 112296 265770 112305
rect 265714 112231 265770 112240
rect 265728 111994 265756 112231
rect 265716 111988 265768 111994
rect 265716 111930 265768 111936
rect 265714 110528 265770 110537
rect 265714 110463 265716 110472
rect 265768 110463 265770 110472
rect 265716 110434 265768 110440
rect 265714 109304 265770 109313
rect 265714 109239 265770 109248
rect 265728 109070 265756 109239
rect 265716 109064 265768 109070
rect 265716 109006 265768 109012
rect 265714 108760 265770 108769
rect 265714 108695 265770 108704
rect 265728 107710 265756 108695
rect 265716 107704 265768 107710
rect 265716 107646 265768 107652
rect 265820 106826 265848 137986
rect 265898 135416 265954 135425
rect 265898 135351 265954 135360
rect 265912 135318 265940 135351
rect 265900 135312 265952 135318
rect 265900 135254 265952 135260
rect 265898 134192 265954 134201
rect 265898 134127 265954 134136
rect 265912 134094 265940 134127
rect 265900 134088 265952 134094
rect 265900 134030 265952 134036
rect 265900 133952 265952 133958
rect 265898 133920 265900 133929
rect 265952 133920 265954 133929
rect 265898 133855 265954 133864
rect 265898 132560 265954 132569
rect 265898 132495 265900 132504
rect 265952 132495 265954 132504
rect 265900 132466 265952 132472
rect 265898 132016 265954 132025
rect 265898 131951 265954 131960
rect 265912 131170 265940 131951
rect 265900 131164 265952 131170
rect 265900 131106 265952 131112
rect 265898 129432 265954 129441
rect 265898 129367 265954 129376
rect 265912 128382 265940 129367
rect 265900 128376 265952 128382
rect 265900 128318 265952 128324
rect 265898 127256 265954 127265
rect 265898 127191 265954 127200
rect 265912 127090 265940 127191
rect 265900 127084 265952 127090
rect 265900 127026 265952 127032
rect 265898 126440 265954 126449
rect 265898 126375 265954 126384
rect 265912 125662 265940 126375
rect 266004 126274 266032 141335
rect 266082 135824 266138 135833
rect 266082 135759 266138 135768
rect 266096 135454 266124 135759
rect 266084 135448 266136 135454
rect 266084 135390 266136 135396
rect 265992 126268 266044 126274
rect 265992 126210 266044 126216
rect 265900 125656 265952 125662
rect 265900 125598 265952 125604
rect 266174 125624 266230 125633
rect 266174 125559 266230 125568
rect 265898 125080 265954 125089
rect 265898 125015 265954 125024
rect 265912 124234 265940 125015
rect 265992 124364 266044 124370
rect 265992 124306 266044 124312
rect 266004 124273 266032 124306
rect 265990 124264 266046 124273
rect 265900 124228 265952 124234
rect 265990 124199 266046 124208
rect 265900 124170 265952 124176
rect 265990 122088 266046 122097
rect 265990 122023 266046 122032
rect 265898 121680 265954 121689
rect 265898 121615 265954 121624
rect 265912 121514 265940 121615
rect 266004 121582 266032 122023
rect 265992 121576 266044 121582
rect 265992 121518 266044 121524
rect 265900 121508 265952 121514
rect 265900 121450 265952 121456
rect 265990 120864 266046 120873
rect 265990 120799 266046 120808
rect 266004 120222 266032 120799
rect 265992 120216 266044 120222
rect 265898 120184 265954 120193
rect 265992 120158 266044 120164
rect 265898 120119 265900 120128
rect 265952 120119 265954 120128
rect 265900 120090 265952 120096
rect 266188 120034 266216 125559
rect 266266 122904 266322 122913
rect 266266 122839 266322 122848
rect 265912 120006 266216 120034
rect 265808 106820 265860 106826
rect 265808 106762 265860 106768
rect 265806 106720 265862 106729
rect 265806 106655 265862 106664
rect 265714 106584 265770 106593
rect 265714 106519 265770 106528
rect 265728 106350 265756 106519
rect 265820 106486 265848 106655
rect 265808 106480 265860 106486
rect 265808 106422 265860 106428
rect 265716 106344 265768 106350
rect 265716 106286 265768 106292
rect 265714 105768 265770 105777
rect 265714 105703 265770 105712
rect 265728 104990 265756 105703
rect 265806 105360 265862 105369
rect 265806 105295 265862 105304
rect 265716 104984 265768 104990
rect 265716 104926 265768 104932
rect 265820 104922 265848 105295
rect 265808 104916 265860 104922
rect 265808 104858 265860 104864
rect 265806 103592 265862 103601
rect 265806 103527 265808 103536
rect 265860 103527 265862 103536
rect 265808 103498 265860 103504
rect 265714 103184 265770 103193
rect 265714 103119 265770 103128
rect 265728 102202 265756 103119
rect 265806 102368 265862 102377
rect 265806 102303 265862 102312
rect 265820 102270 265848 102303
rect 265808 102264 265860 102270
rect 265808 102206 265860 102212
rect 265716 102196 265768 102202
rect 265716 102138 265768 102144
rect 265714 101552 265770 101561
rect 265714 101487 265770 101496
rect 265728 100842 265756 101487
rect 265806 101008 265862 101017
rect 265806 100943 265862 100952
rect 265716 100836 265768 100842
rect 265716 100778 265768 100784
rect 265820 100774 265848 100943
rect 265808 100768 265860 100774
rect 265808 100710 265860 100716
rect 265714 100192 265770 100201
rect 265714 100127 265770 100136
rect 265728 99482 265756 100127
rect 265806 99784 265862 99793
rect 265806 99719 265862 99728
rect 265820 99550 265848 99719
rect 265808 99544 265860 99550
rect 265808 99486 265860 99492
rect 265716 99476 265768 99482
rect 265716 99418 265768 99424
rect 265808 99408 265860 99414
rect 265728 99356 265808 99374
rect 265728 99350 265860 99356
rect 265728 99346 265848 99350
rect 265624 33788 265676 33794
rect 265624 33730 265676 33736
rect 265728 32434 265756 99346
rect 265806 98424 265862 98433
rect 265806 98359 265862 98368
rect 265820 98122 265848 98359
rect 265808 98116 265860 98122
rect 265808 98058 265860 98064
rect 265806 97608 265862 97617
rect 265806 97543 265862 97552
rect 265820 96694 265848 97543
rect 265808 96688 265860 96694
rect 265808 96630 265860 96636
rect 265806 96384 265862 96393
rect 265806 96319 265862 96328
rect 265820 95266 265848 96319
rect 265808 95260 265860 95266
rect 265808 95202 265860 95208
rect 265912 89010 265940 120006
rect 266280 118694 266308 122839
rect 266004 118666 266308 118694
rect 266004 90370 266032 118666
rect 266174 116920 266230 116929
rect 266174 116855 266230 116864
rect 266082 116512 266138 116521
rect 266082 116447 266138 116456
rect 266096 116074 266124 116447
rect 266084 116068 266136 116074
rect 266084 116010 266136 116016
rect 266188 116006 266216 116855
rect 266176 116000 266228 116006
rect 266176 115942 266228 115948
rect 266082 112160 266138 112169
rect 266082 112095 266138 112104
rect 266096 111858 266124 112095
rect 266084 111852 266136 111858
rect 266084 111794 266136 111800
rect 266084 105052 266136 105058
rect 266084 104994 266136 105000
rect 266096 104961 266124 104994
rect 266082 104952 266138 104961
rect 266082 104887 266138 104896
rect 266082 104000 266138 104009
rect 266082 103935 266138 103944
rect 266096 99414 266124 103935
rect 266084 99408 266136 99414
rect 266084 99350 266136 99356
rect 267016 96422 267044 238070
rect 267004 96416 267056 96422
rect 267004 96358 267056 96364
rect 267108 94994 267136 296958
rect 267188 294296 267240 294302
rect 267188 294238 267240 294244
rect 267200 95985 267228 294238
rect 267280 265056 267332 265062
rect 267280 264998 267332 265004
rect 267186 95976 267242 95985
rect 267186 95911 267242 95920
rect 267292 95062 267320 264998
rect 268396 240038 268424 700334
rect 283852 698970 283880 703520
rect 283840 698964 283892 698970
rect 283840 698906 283892 698912
rect 300136 697513 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 300122 697504 300178 697513
rect 300122 697439 300178 697448
rect 269764 630692 269816 630698
rect 269764 630634 269816 630640
rect 268476 299600 268528 299606
rect 268476 299542 268528 299548
rect 268384 240032 268436 240038
rect 268384 239974 268436 239980
rect 268488 178022 268516 299542
rect 269776 238542 269804 630634
rect 270500 514820 270552 514826
rect 270500 514762 270552 514768
rect 269856 296948 269908 296954
rect 269856 296890 269908 296896
rect 269764 238536 269816 238542
rect 269764 238478 269816 238484
rect 269764 228472 269816 228478
rect 269764 228414 269816 228420
rect 268476 178016 268528 178022
rect 268476 177958 268528 177964
rect 269776 175817 269804 228414
rect 269868 177449 269896 296890
rect 270512 248402 270540 514762
rect 331232 315314 331260 702986
rect 348804 702434 348832 703520
rect 347792 702406 348832 702434
rect 347792 693462 347820 702406
rect 364996 699718 365024 703520
rect 359464 699712 359516 699718
rect 359464 699654 359516 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 347780 693456 347832 693462
rect 347780 693398 347832 693404
rect 331220 315308 331272 315314
rect 331220 315250 331272 315256
rect 299480 303680 299532 303686
rect 299480 303622 299532 303628
rect 276664 302320 276716 302326
rect 276664 302262 276716 302268
rect 273904 301028 273956 301034
rect 273904 300970 273956 300976
rect 271236 292596 271288 292602
rect 271236 292538 271288 292544
rect 271144 267776 271196 267782
rect 271144 267718 271196 267724
rect 270500 248396 270552 248402
rect 270500 248338 270552 248344
rect 271156 178838 271184 267718
rect 271248 259418 271276 292538
rect 272524 288516 272576 288522
rect 272524 288458 272576 288464
rect 271236 259412 271288 259418
rect 271236 259354 271288 259360
rect 271236 253972 271288 253978
rect 271236 253914 271288 253920
rect 271144 178832 271196 178838
rect 271144 178774 271196 178780
rect 271248 177478 271276 253914
rect 272536 180198 272564 288458
rect 272524 180192 272576 180198
rect 272524 180134 272576 180140
rect 273916 178906 273944 300970
rect 273996 294364 274048 294370
rect 273996 294306 274048 294312
rect 273904 178900 273956 178906
rect 273904 178842 273956 178848
rect 271236 177472 271288 177478
rect 269854 177440 269910 177449
rect 271236 177414 271288 177420
rect 269854 177375 269910 177384
rect 274008 175953 274036 294306
rect 276676 176186 276704 302262
rect 280804 300960 280856 300966
rect 280804 300902 280856 300908
rect 278044 298308 278096 298314
rect 278044 298250 278096 298256
rect 276756 266484 276808 266490
rect 276756 266426 276808 266432
rect 276768 180334 276796 266426
rect 276848 258120 276900 258126
rect 276848 258062 276900 258068
rect 276756 180328 276808 180334
rect 276756 180270 276808 180276
rect 276860 177410 276888 258062
rect 276940 188420 276992 188426
rect 276940 188362 276992 188368
rect 276848 177404 276900 177410
rect 276848 177346 276900 177352
rect 276664 176180 276716 176186
rect 276664 176122 276716 176128
rect 276952 176050 276980 188362
rect 278056 176118 278084 298250
rect 278136 282940 278188 282946
rect 278136 282882 278188 282888
rect 278148 184346 278176 282882
rect 280160 196648 280212 196654
rect 280160 196590 280212 196596
rect 278136 184340 278188 184346
rect 278136 184282 278188 184288
rect 279422 177576 279478 177585
rect 279422 177511 279478 177520
rect 279332 176180 279384 176186
rect 279332 176122 279384 176128
rect 278044 176112 278096 176118
rect 278044 176054 278096 176060
rect 276940 176044 276992 176050
rect 276940 175986 276992 175992
rect 273994 175944 274050 175953
rect 273994 175879 274050 175888
rect 269762 175808 269818 175817
rect 269762 175743 269818 175752
rect 279344 173777 279372 176122
rect 279436 174457 279464 177511
rect 279422 174448 279478 174457
rect 279422 174383 279478 174392
rect 279330 173768 279386 173777
rect 279330 173703 279386 173712
rect 280172 136377 280200 196590
rect 280816 191185 280844 300902
rect 298100 299668 298152 299674
rect 298100 299610 298152 299616
rect 296720 295520 296772 295526
rect 282918 295488 282974 295497
rect 296720 295462 296772 295468
rect 282918 295423 282974 295432
rect 291200 295452 291252 295458
rect 281632 236700 281684 236706
rect 281632 236642 281684 236648
rect 281538 236600 281594 236609
rect 281538 236535 281594 236544
rect 280802 191176 280858 191185
rect 280802 191111 280858 191120
rect 280344 180260 280396 180266
rect 280344 180202 280396 180208
rect 280252 175976 280304 175982
rect 280252 175918 280304 175924
rect 280264 151745 280292 175918
rect 280356 172417 280384 180202
rect 280342 172408 280398 172417
rect 280342 172343 280398 172352
rect 281552 161474 281580 236535
rect 281644 167793 281672 236642
rect 281724 204944 281776 204950
rect 281724 204886 281776 204892
rect 281736 168609 281764 204886
rect 282736 171080 282788 171086
rect 282736 171022 282788 171028
rect 282748 170105 282776 171022
rect 282828 171012 282880 171018
rect 282828 170954 282880 170960
rect 282840 170921 282868 170954
rect 282826 170912 282882 170921
rect 282826 170847 282882 170856
rect 282734 170096 282790 170105
rect 282734 170031 282790 170040
rect 282828 169720 282880 169726
rect 282828 169662 282880 169668
rect 282840 169425 282868 169662
rect 282826 169416 282882 169425
rect 282826 169351 282882 169360
rect 281722 168600 281778 168609
rect 281722 168535 281778 168544
rect 282460 168360 282512 168366
rect 282460 168302 282512 168308
rect 281630 167784 281686 167793
rect 281630 167719 281686 167728
rect 282472 167113 282500 168302
rect 282458 167104 282514 167113
rect 282458 167039 282514 167048
rect 282092 167000 282144 167006
rect 282092 166942 282144 166948
rect 282104 166297 282132 166942
rect 282090 166288 282146 166297
rect 282090 166223 282146 166232
rect 282000 165572 282052 165578
rect 282000 165514 282052 165520
rect 282012 164801 282040 165514
rect 282828 165504 282880 165510
rect 282826 165472 282828 165481
rect 282880 165472 282882 165481
rect 282826 165407 282882 165416
rect 281998 164792 282054 164801
rect 281998 164727 282054 164736
rect 282828 164212 282880 164218
rect 282828 164154 282880 164160
rect 282090 163976 282146 163985
rect 282090 163911 282146 163920
rect 282104 163266 282132 163911
rect 282092 163260 282144 163266
rect 282092 163202 282144 163208
rect 282840 163169 282868 164154
rect 282826 163160 282882 163169
rect 282826 163095 282882 163104
rect 282092 162852 282144 162858
rect 282092 162794 282144 162800
rect 282104 162489 282132 162794
rect 282828 162784 282880 162790
rect 282828 162726 282880 162732
rect 282090 162480 282146 162489
rect 282090 162415 282146 162424
rect 282840 161673 282868 162726
rect 282826 161664 282882 161673
rect 282826 161599 282882 161608
rect 281552 161446 281672 161474
rect 281540 160676 281592 160682
rect 281540 160618 281592 160624
rect 281552 160177 281580 160618
rect 281538 160168 281594 160177
rect 281538 160103 281594 160112
rect 281540 160064 281592 160070
rect 281540 160006 281592 160012
rect 281552 159361 281580 160006
rect 281538 159352 281594 159361
rect 281538 159287 281594 159296
rect 281644 154737 281672 161446
rect 282828 161424 282880 161430
rect 282828 161366 282880 161372
rect 282840 160857 282868 161366
rect 282826 160848 282882 160857
rect 282826 160783 282882 160792
rect 282736 158704 282788 158710
rect 282736 158646 282788 158652
rect 282748 157865 282776 158646
rect 282828 158636 282880 158642
rect 282828 158578 282880 158584
rect 282840 158545 282868 158578
rect 282826 158536 282882 158545
rect 282826 158471 282882 158480
rect 282734 157856 282790 157865
rect 282734 157791 282790 157800
rect 281724 156596 281776 156602
rect 281724 156538 281776 156544
rect 281736 156369 281764 156538
rect 281722 156360 281778 156369
rect 281722 156295 281778 156304
rect 281630 154728 281686 154737
rect 281630 154663 281686 154672
rect 281724 154556 281776 154562
rect 281724 154498 281776 154504
rect 281736 154057 281764 154498
rect 281722 154048 281778 154057
rect 281722 153983 281778 153992
rect 282828 153468 282880 153474
rect 282828 153410 282880 153416
rect 282840 153241 282868 153410
rect 282826 153232 282882 153241
rect 282736 153196 282788 153202
rect 282826 153167 282882 153176
rect 282736 153138 282788 153144
rect 282748 152425 282776 153138
rect 282734 152416 282790 152425
rect 282734 152351 282790 152360
rect 282828 151768 282880 151774
rect 280250 151736 280306 151745
rect 282828 151710 282880 151716
rect 280250 151671 280306 151680
rect 282840 150929 282868 151710
rect 282826 150920 282882 150929
rect 282826 150855 282882 150864
rect 282828 150408 282880 150414
rect 282828 150350 282880 150356
rect 282840 150113 282868 150350
rect 282826 150104 282882 150113
rect 282826 150039 282882 150048
rect 281540 149660 281592 149666
rect 281540 149602 281592 149608
rect 281552 149433 281580 149602
rect 281538 149424 281594 149433
rect 281538 149359 281594 149368
rect 282828 149048 282880 149054
rect 282828 148990 282880 148996
rect 282276 148640 282328 148646
rect 282840 148617 282868 148990
rect 282276 148582 282328 148588
rect 282826 148608 282882 148617
rect 282288 147801 282316 148582
rect 282826 148543 282882 148552
rect 282274 147792 282330 147801
rect 282274 147727 282330 147736
rect 281724 147620 281776 147626
rect 281724 147562 281776 147568
rect 281736 147121 281764 147562
rect 281722 147112 281778 147121
rect 281722 147047 281778 147056
rect 282826 146296 282882 146305
rect 282000 146260 282052 146266
rect 282826 146231 282882 146240
rect 282000 146202 282052 146208
rect 282012 145489 282040 146202
rect 282840 146198 282868 146231
rect 282828 146192 282880 146198
rect 282828 146134 282880 146140
rect 281998 145480 282054 145489
rect 281998 145415 282054 145424
rect 282552 144832 282604 144838
rect 282550 144800 282552 144809
rect 282604 144800 282606 144809
rect 282550 144735 282606 144744
rect 282826 143984 282882 143993
rect 282826 143919 282882 143928
rect 282840 143750 282868 143919
rect 282828 143744 282880 143750
rect 282828 143686 282880 143692
rect 281632 143540 281684 143546
rect 281632 143482 281684 143488
rect 281644 142497 281672 143482
rect 281630 142488 281686 142497
rect 281630 142423 281686 142432
rect 282828 142112 282880 142118
rect 282828 142054 282880 142060
rect 282840 141681 282868 142054
rect 282826 141672 282882 141681
rect 282826 141607 282882 141616
rect 281908 140752 281960 140758
rect 281908 140694 281960 140700
rect 281920 140185 281948 140694
rect 281906 140176 281962 140185
rect 281906 140111 281962 140120
rect 282828 139392 282880 139398
rect 282826 139360 282828 139369
rect 282880 139360 282882 139369
rect 282736 139324 282788 139330
rect 282826 139295 282882 139304
rect 282736 139266 282788 139272
rect 282748 138553 282776 139266
rect 282734 138544 282790 138553
rect 282734 138479 282790 138488
rect 282184 137964 282236 137970
rect 282184 137906 282236 137912
rect 282196 137057 282224 137906
rect 282828 137896 282880 137902
rect 282826 137864 282828 137873
rect 282880 137864 282882 137873
rect 282826 137799 282882 137808
rect 282182 137048 282238 137057
rect 282182 136983 282238 136992
rect 280158 136368 280214 136377
rect 280158 136303 280214 136312
rect 282826 134056 282882 134065
rect 282932 134042 282960 295423
rect 291200 295394 291252 295400
rect 285678 292360 285734 292369
rect 285678 292295 285734 292304
rect 283104 277432 283156 277438
rect 283104 277374 283156 277380
rect 283012 273964 283064 273970
rect 283012 273906 283064 273912
rect 282882 134014 282960 134042
rect 282826 133991 282882 134000
rect 282828 133884 282880 133890
rect 282828 133826 282880 133832
rect 282840 133249 282868 133826
rect 282826 133240 282882 133249
rect 282826 133175 282882 133184
rect 283024 132494 283052 273906
rect 283116 155553 283144 277374
rect 284300 250504 284352 250510
rect 284300 250446 284352 250452
rect 283194 177304 283250 177313
rect 283194 177239 283250 177248
rect 283208 160682 283236 177239
rect 283196 160676 283248 160682
rect 283196 160618 283248 160624
rect 283102 155544 283158 155553
rect 283102 155479 283158 155488
rect 284312 149666 284340 250446
rect 284484 231124 284536 231130
rect 284484 231066 284536 231072
rect 284392 188488 284444 188494
rect 284392 188430 284444 188436
rect 284300 149660 284352 149666
rect 284300 149602 284352 149608
rect 282932 132466 283052 132494
rect 282828 132456 282880 132462
rect 282826 132424 282828 132433
rect 282880 132424 282882 132433
rect 282826 132359 282882 132368
rect 282828 131096 282880 131102
rect 282828 131038 282880 131044
rect 282840 130937 282868 131038
rect 282826 130928 282882 130937
rect 282826 130863 282882 130872
rect 282276 130620 282328 130626
rect 282276 130562 282328 130568
rect 282288 130121 282316 130562
rect 282274 130112 282330 130121
rect 282274 130047 282330 130056
rect 282826 128616 282882 128625
rect 282826 128551 282882 128560
rect 282840 128518 282868 128551
rect 282828 128512 282880 128518
rect 282828 128454 282880 128460
rect 281724 128308 281776 128314
rect 281724 128250 281776 128256
rect 281736 127809 281764 128250
rect 281722 127800 281778 127809
rect 281722 127735 281778 127744
rect 282826 126304 282882 126313
rect 282932 126290 282960 132466
rect 282882 126262 282960 126290
rect 282826 126239 282882 126248
rect 282092 125588 282144 125594
rect 282092 125530 282144 125536
rect 282104 124817 282132 125530
rect 282826 125488 282882 125497
rect 282826 125423 282882 125432
rect 282090 124808 282146 124817
rect 282090 124743 282146 124752
rect 282840 124710 282868 125423
rect 282828 124704 282880 124710
rect 282828 124646 282880 124652
rect 282736 124160 282788 124166
rect 282736 124102 282788 124108
rect 282748 123185 282776 124102
rect 282828 124092 282880 124098
rect 282828 124034 282880 124040
rect 282840 124001 282868 124034
rect 282826 123992 282882 124001
rect 282826 123927 282882 123936
rect 282734 123176 282790 123185
rect 282734 123111 282790 123120
rect 282092 122800 282144 122806
rect 282092 122742 282144 122748
rect 282104 122505 282132 122742
rect 282090 122496 282146 122505
rect 282090 122431 282146 122440
rect 282460 121440 282512 121446
rect 282460 121382 282512 121388
rect 281724 121372 281776 121378
rect 281724 121314 281776 121320
rect 281736 120873 281764 121314
rect 281722 120864 281778 120873
rect 281722 120799 281778 120808
rect 282472 120193 282500 121382
rect 282458 120184 282514 120193
rect 282458 120119 282514 120128
rect 282092 120080 282144 120086
rect 282092 120022 282144 120028
rect 282104 119377 282132 120022
rect 282090 119368 282146 119377
rect 282090 119303 282146 119312
rect 282828 118652 282880 118658
rect 282828 118594 282880 118600
rect 282736 118584 282788 118590
rect 282840 118561 282868 118594
rect 282736 118526 282788 118532
rect 282826 118552 282882 118561
rect 282748 117881 282776 118526
rect 282826 118487 282882 118496
rect 282734 117872 282790 117881
rect 282734 117807 282790 117816
rect 282828 117292 282880 117298
rect 282828 117234 282880 117240
rect 282736 117224 282788 117230
rect 282736 117166 282788 117172
rect 282748 116385 282776 117166
rect 282840 117065 282868 117234
rect 282826 117056 282882 117065
rect 282826 116991 282882 117000
rect 282734 116376 282790 116385
rect 282734 116311 282790 116320
rect 281724 115932 281776 115938
rect 281724 115874 281776 115880
rect 281736 114753 281764 115874
rect 282092 115864 282144 115870
rect 282092 115806 282144 115812
rect 282104 115569 282132 115806
rect 282090 115560 282146 115569
rect 282090 115495 282146 115504
rect 281722 114744 281778 114753
rect 281722 114679 281778 114688
rect 282826 114064 282882 114073
rect 282826 113999 282882 114008
rect 282840 113966 282868 113999
rect 282828 113960 282880 113966
rect 282828 113902 282880 113908
rect 282092 113144 282144 113150
rect 282092 113086 282144 113092
rect 282104 112441 282132 113086
rect 282090 112432 282146 112441
rect 282090 112367 282146 112376
rect 282828 111784 282880 111790
rect 282826 111752 282828 111761
rect 282880 111752 282882 111761
rect 282826 111687 282882 111696
rect 280158 110936 280214 110945
rect 280158 110871 280214 110880
rect 279422 98152 279478 98161
rect 279422 98087 279478 98096
rect 279330 96656 279386 96665
rect 279330 96591 279386 96600
rect 268016 95940 268068 95946
rect 268016 95882 268068 95888
rect 267280 95056 267332 95062
rect 267280 94998 267332 95004
rect 267096 94988 267148 94994
rect 267096 94930 267148 94936
rect 268028 93838 268056 95882
rect 268016 93832 268068 93838
rect 268016 93774 268068 93780
rect 270972 93770 271000 96016
rect 276952 93838 276980 96016
rect 279344 95985 279372 96591
rect 279330 95976 279386 95985
rect 279330 95911 279386 95920
rect 279436 95169 279464 98087
rect 279514 97336 279570 97345
rect 279514 97271 279570 97280
rect 279422 95160 279478 95169
rect 279422 95095 279478 95104
rect 279528 95062 279556 97271
rect 280066 95840 280122 95849
rect 280066 95775 280122 95784
rect 279516 95056 279568 95062
rect 279516 94998 279568 95004
rect 276940 93832 276992 93838
rect 276940 93774 276992 93780
rect 270960 93764 271012 93770
rect 270960 93706 271012 93712
rect 280080 93673 280108 95775
rect 280172 95198 280200 110871
rect 282828 108996 282880 109002
rect 282828 108938 282880 108944
rect 282840 108633 282868 108938
rect 282826 108624 282882 108633
rect 282826 108559 282882 108568
rect 284404 108050 284432 188430
rect 284496 160070 284524 231066
rect 284576 202156 284628 202162
rect 284576 202098 284628 202104
rect 284484 160064 284536 160070
rect 284484 160006 284536 160012
rect 284588 156602 284616 202098
rect 284576 156596 284628 156602
rect 284576 156538 284628 156544
rect 285692 125594 285720 292295
rect 287060 272536 287112 272542
rect 287060 272478 287112 272484
rect 285772 206304 285824 206310
rect 285772 206246 285824 206252
rect 285784 144838 285812 206246
rect 285864 185632 285916 185638
rect 285864 185574 285916 185580
rect 285772 144832 285824 144838
rect 285772 144774 285824 144780
rect 285876 130626 285904 185574
rect 287072 143750 287100 272478
rect 290096 266416 290148 266422
rect 290096 266358 290148 266364
rect 287152 232688 287204 232694
rect 287152 232630 287204 232636
rect 287060 143744 287112 143750
rect 287060 143686 287112 143692
rect 285864 130620 285916 130626
rect 285864 130562 285916 130568
rect 287164 128518 287192 232630
rect 287244 211812 287296 211818
rect 287244 211754 287296 211760
rect 287256 153474 287284 211754
rect 287336 200796 287388 200802
rect 287336 200738 287388 200744
rect 287244 153468 287296 153474
rect 287244 153410 287296 153416
rect 287348 148646 287376 200738
rect 288624 189916 288676 189922
rect 288624 189858 288676 189864
rect 288440 184272 288492 184278
rect 288440 184214 288492 184220
rect 287336 148640 287388 148646
rect 287336 148582 287388 148588
rect 287152 128512 287204 128518
rect 287152 128454 287204 128460
rect 285680 125588 285732 125594
rect 285680 125530 285732 125536
rect 288452 113966 288480 184214
rect 288532 177472 288584 177478
rect 288532 177414 288584 177420
rect 288544 124710 288572 177414
rect 288636 163266 288664 189858
rect 289912 184204 289964 184210
rect 289912 184146 289964 184152
rect 288716 180328 288768 180334
rect 288716 180270 288768 180276
rect 288624 163260 288676 163266
rect 288624 163202 288676 163208
rect 288728 158642 288756 180270
rect 289820 176044 289872 176050
rect 289820 175986 289872 175992
rect 289832 169726 289860 175986
rect 289820 169720 289872 169726
rect 289820 169662 289872 169668
rect 288716 158636 288768 158642
rect 288716 158578 288768 158584
rect 288532 124704 288584 124710
rect 288532 124646 288584 124652
rect 289924 118590 289952 184146
rect 290004 176112 290056 176118
rect 290004 176054 290056 176060
rect 290016 171018 290044 176054
rect 290004 171012 290056 171018
rect 290004 170954 290056 170960
rect 290108 149054 290136 266358
rect 291212 161430 291240 295394
rect 295340 280220 295392 280226
rect 295340 280162 295392 280168
rect 293960 260908 294012 260914
rect 293960 260850 294012 260856
rect 292856 244316 292908 244322
rect 292856 244258 292908 244264
rect 292764 195288 292816 195294
rect 292764 195230 292816 195236
rect 292672 187060 292724 187066
rect 292672 187002 292724 187008
rect 291384 185700 291436 185706
rect 291384 185642 291436 185648
rect 291292 180124 291344 180130
rect 291292 180066 291344 180072
rect 291200 161424 291252 161430
rect 291200 161366 291252 161372
rect 290096 149048 290148 149054
rect 290096 148990 290148 148996
rect 291304 121378 291332 180066
rect 291396 150414 291424 185642
rect 291476 178764 291528 178770
rect 291476 178706 291528 178712
rect 291488 165510 291516 178706
rect 292580 177336 292632 177342
rect 292580 177278 292632 177284
rect 292592 168366 292620 177278
rect 292580 168360 292632 168366
rect 292580 168302 292632 168308
rect 291476 165504 291528 165510
rect 291476 165446 291528 165452
rect 291384 150408 291436 150414
rect 291384 150350 291436 150356
rect 291292 121372 291344 121378
rect 291292 121314 291344 121320
rect 292684 118658 292712 187002
rect 292776 139330 292804 195230
rect 292868 162790 292896 244258
rect 292856 162784 292908 162790
rect 292856 162726 292908 162732
rect 292764 139324 292816 139330
rect 292764 139266 292816 139272
rect 293972 137902 294000 260850
rect 294144 185768 294196 185774
rect 294144 185710 294196 185716
rect 294052 178832 294104 178838
rect 294052 178774 294104 178780
rect 293960 137896 294012 137902
rect 293960 137838 294012 137844
rect 292672 118652 292724 118658
rect 292672 118594 292724 118600
rect 289912 118584 289964 118590
rect 289912 118526 289964 118532
rect 288440 113960 288492 113966
rect 288440 113902 288492 113908
rect 294064 113150 294092 178774
rect 294156 165578 294184 185710
rect 294234 178664 294290 178673
rect 294234 178599 294290 178608
rect 294248 167006 294276 178599
rect 294236 167000 294288 167006
rect 294236 166942 294288 166948
rect 294144 165572 294196 165578
rect 294144 165514 294196 165520
rect 295352 124098 295380 280162
rect 295524 189848 295576 189854
rect 295524 189790 295576 189796
rect 295432 181484 295484 181490
rect 295432 181426 295484 181432
rect 295340 124092 295392 124098
rect 295340 124034 295392 124040
rect 295444 117230 295472 181426
rect 295536 164218 295564 189790
rect 295616 178900 295668 178906
rect 295616 178842 295668 178848
rect 295524 164212 295576 164218
rect 295524 164154 295576 164160
rect 295628 158710 295656 178842
rect 296628 178016 296680 178022
rect 296628 177958 296680 177964
rect 296640 171193 296668 177958
rect 296626 171184 296682 171193
rect 296626 171119 296682 171128
rect 295616 158704 295668 158710
rect 295616 158646 295668 158652
rect 296732 146198 296760 295462
rect 296812 288448 296864 288454
rect 296812 288390 296864 288396
rect 296720 146192 296772 146198
rect 296720 146134 296772 146140
rect 296824 140758 296852 288390
rect 296904 188352 296956 188358
rect 296904 188294 296956 188300
rect 296812 140752 296864 140758
rect 296812 140694 296864 140700
rect 295432 117224 295484 117230
rect 295432 117166 295484 117172
rect 296916 115870 296944 188294
rect 296996 182844 297048 182850
rect 296996 182786 297048 182792
rect 297008 171086 297036 182786
rect 296996 171080 297048 171086
rect 296996 171022 297048 171028
rect 298112 162858 298140 299610
rect 298192 245676 298244 245682
rect 298192 245618 298244 245624
rect 298100 162852 298152 162858
rect 298100 162794 298152 162800
rect 298204 120086 298232 245618
rect 298284 182912 298336 182918
rect 298284 182854 298336 182860
rect 298192 120080 298244 120086
rect 298192 120022 298244 120028
rect 296904 115864 296956 115870
rect 296904 115806 296956 115812
rect 294052 113144 294104 113150
rect 294052 113086 294104 113092
rect 281540 108044 281592 108050
rect 281540 107986 281592 107992
rect 284392 108044 284444 108050
rect 284392 107986 284444 107992
rect 281552 107817 281580 107986
rect 281538 107808 281594 107817
rect 281538 107743 281594 107752
rect 298296 107642 298324 182854
rect 298374 180024 298430 180033
rect 298374 179959 298430 179968
rect 298388 137970 298416 179959
rect 298376 137964 298428 137970
rect 298376 137906 298428 137912
rect 282460 107636 282512 107642
rect 282460 107578 282512 107584
rect 298284 107636 298336 107642
rect 298284 107578 298336 107584
rect 280250 107128 280306 107137
rect 280250 107063 280306 107072
rect 280160 95192 280212 95198
rect 280160 95134 280212 95140
rect 280066 93664 280122 93673
rect 280066 93599 280122 93608
rect 280264 93537 280292 107063
rect 282472 106321 282500 107578
rect 282458 106312 282514 106321
rect 282458 106247 282514 106256
rect 282828 106276 282880 106282
rect 282828 106218 282880 106224
rect 282840 105505 282868 106218
rect 282826 105496 282882 105505
rect 282826 105431 282882 105440
rect 282458 104952 282514 104961
rect 282458 104887 282514 104896
rect 280342 104816 280398 104825
rect 280342 104751 280398 104760
rect 280356 94994 280384 104751
rect 282472 102513 282500 104887
rect 282828 103488 282880 103494
rect 282828 103430 282880 103436
rect 282840 103193 282868 103430
rect 282826 103184 282882 103193
rect 282826 103119 282882 103128
rect 282458 102504 282514 102513
rect 282458 102439 282514 102448
rect 281630 101688 281686 101697
rect 281630 101623 281686 101632
rect 281538 100192 281594 100201
rect 281538 100127 281594 100136
rect 281552 96422 281580 100127
rect 281540 96416 281592 96422
rect 281540 96358 281592 96364
rect 281644 95130 281672 101623
rect 281814 100872 281870 100881
rect 281814 100807 281870 100816
rect 281632 95124 281684 95130
rect 281632 95066 281684 95072
rect 280344 94988 280396 94994
rect 280344 94930 280396 94936
rect 280250 93528 280306 93537
rect 280250 93463 280306 93472
rect 281828 92478 281856 100807
rect 282826 99376 282882 99385
rect 299492 99346 299520 303622
rect 316040 302252 316092 302258
rect 316040 302194 316092 302200
rect 302240 299532 302292 299538
rect 302240 299474 302292 299480
rect 299572 298240 299624 298246
rect 299572 298182 299624 298188
rect 299584 111790 299612 298182
rect 300860 262268 300912 262274
rect 300860 262210 300912 262216
rect 299664 191140 299716 191146
rect 299664 191082 299716 191088
rect 299572 111784 299624 111790
rect 299572 111726 299624 111732
rect 299676 103494 299704 191082
rect 299756 189780 299808 189786
rect 299756 189722 299808 189728
rect 299768 146266 299796 189722
rect 299756 146260 299808 146266
rect 299756 146202 299808 146208
rect 300872 124166 300900 262210
rect 300952 238060 301004 238066
rect 300952 238002 301004 238008
rect 300964 154562 300992 238002
rect 301044 180192 301096 180198
rect 301044 180134 301096 180140
rect 300952 154556 301004 154562
rect 300952 154498 301004 154504
rect 301056 143546 301084 180134
rect 301136 178696 301188 178702
rect 301136 178638 301188 178644
rect 301148 151774 301176 178638
rect 301136 151768 301188 151774
rect 301136 151710 301188 151716
rect 301044 143540 301096 143546
rect 301044 143482 301096 143488
rect 300860 124160 300912 124166
rect 300860 124102 300912 124108
rect 302252 121446 302280 299474
rect 303620 298172 303672 298178
rect 303620 298114 303672 298120
rect 302884 232552 302936 232558
rect 302884 232494 302936 232500
rect 302332 177404 302384 177410
rect 302332 177346 302384 177352
rect 302344 131102 302372 177346
rect 302332 131096 302384 131102
rect 302332 131038 302384 131044
rect 302240 121440 302292 121446
rect 302240 121382 302292 121388
rect 299664 103488 299716 103494
rect 299664 103430 299716 103436
rect 282826 99311 282828 99320
rect 282880 99311 282882 99320
rect 299480 99340 299532 99346
rect 282828 99282 282880 99288
rect 299480 99282 299532 99288
rect 281816 92472 281868 92478
rect 281816 92414 281868 92420
rect 265992 90364 266044 90370
rect 265992 90306 266044 90312
rect 265900 89004 265952 89010
rect 265900 88946 265952 88952
rect 302896 33114 302924 232494
rect 303632 115938 303660 298114
rect 309140 295384 309192 295390
rect 309140 295326 309192 295332
rect 305644 287088 305696 287094
rect 305644 287030 305696 287036
rect 303712 264988 303764 264994
rect 303712 264930 303764 264936
rect 303724 142118 303752 264930
rect 305000 252612 305052 252618
rect 305000 252554 305052 252560
rect 303804 186992 303856 186998
rect 303804 186934 303856 186940
rect 303712 142112 303764 142118
rect 303712 142054 303764 142060
rect 303816 128314 303844 186934
rect 305012 153202 305040 252554
rect 305092 193860 305144 193866
rect 305092 193802 305144 193808
rect 305000 153196 305052 153202
rect 305000 153138 305052 153144
rect 303804 128308 303856 128314
rect 303804 128250 303856 128256
rect 303620 115932 303672 115938
rect 303620 115874 303672 115880
rect 305104 106282 305132 193802
rect 305656 126954 305684 287030
rect 306380 248464 306432 248470
rect 306380 248406 306432 248412
rect 305644 126948 305696 126954
rect 305644 126890 305696 126896
rect 306392 109002 306420 248406
rect 306472 233912 306524 233918
rect 306472 233854 306524 233860
rect 306484 117298 306512 233854
rect 307760 184340 307812 184346
rect 307760 184282 307812 184288
rect 307772 132462 307800 184282
rect 307760 132456 307812 132462
rect 307760 132398 307812 132404
rect 309152 122806 309180 295326
rect 313278 292224 313334 292233
rect 313278 292159 313334 292168
rect 311900 240168 311952 240174
rect 311900 240110 311952 240116
rect 311912 133890 311940 240110
rect 313292 139398 313320 292159
rect 316052 147626 316080 302194
rect 359476 238610 359504 699654
rect 397472 697610 397500 703520
rect 397460 697604 397512 697610
rect 397460 697546 397512 697552
rect 367744 696992 367796 696998
rect 367744 696934 367796 696940
rect 367756 301510 367784 696934
rect 411904 683188 411956 683194
rect 411904 683130 411956 683136
rect 410524 470620 410576 470626
rect 410524 470562 410576 470568
rect 407764 378208 407816 378214
rect 407764 378150 407816 378156
rect 367744 301504 367796 301510
rect 367744 301446 367796 301452
rect 407776 291174 407804 378150
rect 407764 291168 407816 291174
rect 407764 291110 407816 291116
rect 381544 285728 381596 285734
rect 381544 285670 381596 285676
rect 359464 238604 359516 238610
rect 359464 238546 359516 238552
rect 322204 235272 322256 235278
rect 322204 235214 322256 235220
rect 316040 147620 316092 147626
rect 316040 147562 316092 147568
rect 313280 139392 313332 139398
rect 313280 139334 313332 139340
rect 311900 133884 311952 133890
rect 311900 133826 311952 133832
rect 309140 122800 309192 122806
rect 309140 122742 309192 122748
rect 306472 117292 306524 117298
rect 306472 117234 306524 117240
rect 306380 108996 306432 109002
rect 306380 108938 306432 108944
rect 305092 106276 305144 106282
rect 305092 106218 305144 106224
rect 322216 46918 322244 235214
rect 381556 153202 381584 285670
rect 410536 285666 410564 470562
rect 410524 285660 410576 285666
rect 410524 285602 410576 285608
rect 385684 274712 385736 274718
rect 385684 274654 385736 274660
rect 382924 259480 382976 259486
rect 382924 259422 382976 259428
rect 382936 167006 382964 259422
rect 382924 167000 382976 167006
rect 382924 166942 382976 166948
rect 381544 153196 381596 153202
rect 381544 153138 381596 153144
rect 385696 100706 385724 274654
rect 411916 252550 411944 683130
rect 412652 309806 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700330 429884 703520
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 462332 696250 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 696244 462372 696250
rect 462320 696186 462372 696192
rect 477512 694822 477540 702406
rect 494808 700398 494836 703520
rect 494796 700392 494848 700398
rect 494796 700334 494848 700340
rect 527192 700330 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 504364 700324 504416 700330
rect 504364 700266 504416 700272
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 477500 694816 477552 694822
rect 477500 694758 477552 694764
rect 428464 484424 428516 484430
rect 428464 484366 428516 484372
rect 425704 430636 425756 430642
rect 425704 430578 425756 430584
rect 412640 309800 412692 309806
rect 412640 309742 412692 309748
rect 425716 256630 425744 430578
rect 428476 264926 428504 484366
rect 504376 300150 504404 700266
rect 504364 300144 504416 300150
rect 504364 300086 504416 300092
rect 428464 264920 428516 264926
rect 428464 264862 428516 264868
rect 425704 256624 425756 256630
rect 425704 256566 425756 256572
rect 411904 252544 411956 252550
rect 411904 252486 411956 252492
rect 542372 234598 542400 702406
rect 559668 700330 559696 703520
rect 547144 700324 547196 700330
rect 547144 700266 547196 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 547156 242894 547184 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 582378 617536 582434 617545
rect 582378 617471 582434 617480
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580264 282192 580316 282198
rect 580264 282134 580316 282140
rect 566464 276072 566516 276078
rect 566464 276014 566516 276020
rect 547144 242888 547196 242894
rect 547144 242830 547196 242836
rect 542360 234592 542412 234598
rect 542360 234534 542412 234540
rect 566476 233238 566504 276014
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 574744 271924 574796 271930
rect 574744 271866 574796 271872
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 574756 238678 574784 271866
rect 579620 259412 579672 259418
rect 579620 259354 579672 259360
rect 579632 258913 579660 259354
rect 579618 258904 579674 258913
rect 579618 258839 579674 258848
rect 579894 245576 579950 245585
rect 579894 245511 579950 245520
rect 579908 244322 579936 245511
rect 579896 244316 579948 244322
rect 579896 244258 579948 244264
rect 574744 238672 574796 238678
rect 574744 238614 574796 238620
rect 566464 233232 566516 233238
rect 566464 233174 566516 233180
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 579896 206984 579948 206990
rect 579896 206926 579948 206932
rect 579908 205737 579936 206926
rect 579894 205728 579950 205737
rect 579894 205663 579950 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579804 153196 579856 153202
rect 579804 153138 579856 153144
rect 579816 152697 579844 153138
rect 579802 152688 579858 152697
rect 579802 152623 579858 152632
rect 580276 139369 580304 282134
rect 580356 271176 580408 271182
rect 580356 271118 580408 271124
rect 580368 179217 580396 271118
rect 582392 256698 582420 617471
rect 582470 591016 582526 591025
rect 582470 590951 582526 590960
rect 582380 256692 582432 256698
rect 582380 256634 582432 256640
rect 582484 240106 582512 590951
rect 582562 537840 582618 537849
rect 582562 537775 582618 537784
rect 582472 240100 582524 240106
rect 582472 240042 582524 240048
rect 582576 237386 582604 537775
rect 582930 365120 582986 365129
rect 582930 365055 582986 365064
rect 582840 300892 582892 300898
rect 582840 300834 582892 300840
rect 582746 295352 582802 295361
rect 582746 295287 582802 295296
rect 582654 293992 582710 294001
rect 582654 293927 582710 293936
rect 582564 237380 582616 237386
rect 582564 237322 582616 237328
rect 582378 182880 582434 182889
rect 582378 182815 582434 182824
rect 580354 179208 580410 179217
rect 580354 179143 580410 179152
rect 580262 139360 580318 139369
rect 580262 139295 580318 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 385684 100700 385736 100706
rect 385684 100642 385736 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 582392 86193 582420 182815
rect 582378 86184 582434 86193
rect 582378 86119 582434 86128
rect 322204 46912 322256 46918
rect 322204 46854 322256 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 302884 33108 302936 33114
rect 580170 33079 580172 33088
rect 302884 33050 302936 33056
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 265716 32428 265768 32434
rect 265716 32370 265768 32376
rect 264428 26988 264480 26994
rect 264428 26930 264480 26936
rect 582668 19825 582696 293927
rect 582760 73001 582788 295287
rect 582852 112849 582880 300834
rect 582944 235958 582972 365055
rect 583114 298752 583170 298761
rect 583114 298687 583170 298696
rect 583024 296744 583076 296750
rect 583024 296686 583076 296692
rect 582932 235952 582984 235958
rect 582932 235894 582984 235900
rect 583036 219065 583064 296686
rect 583128 238746 583156 298687
rect 583116 238740 583168 238746
rect 583116 238682 583168 238688
rect 583022 219056 583078 219065
rect 583022 218991 583078 219000
rect 582838 112840 582894 112849
rect 582838 112775 582894 112784
rect 582746 72992 582802 73001
rect 582746 72927 582802 72936
rect 582654 19816 582710 19825
rect 582654 19751 582710 19760
rect 264244 18692 264296 18698
rect 264244 18634 264296 18640
rect 260196 7608 260248 7614
rect 260196 7550 260248 7556
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 249064 6248 249116 6254
rect 249064 6190 249116 6196
rect 238024 4820 238076 4826
rect 238024 4762 238076 4768
rect 233976 3528 234028 3534
rect 233976 3470 234028 3476
rect 235816 3528 235868 3534
rect 235816 3470 235868 3476
rect 215944 3460 215996 3466
rect 215944 3402 215996 3408
rect 235828 480 235856 3470
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 2962 527856 3018 527912
rect 3054 501744 3110 501800
rect 3054 475632 3110 475688
rect 3146 449520 3202 449576
rect 2778 423564 2834 423600
rect 2778 423544 2780 423564
rect 2780 423544 2832 423564
rect 2832 423544 2834 423564
rect 2870 410488 2926 410544
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3238 306176 3294 306232
rect 3514 671200 3570 671256
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 462576 3570 462632
rect 3514 371320 3570 371376
rect 3422 293120 3478 293176
rect 3422 290808 3478 290864
rect 3146 254088 3202 254144
rect 3054 241032 3110 241088
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3606 267144 3662 267200
rect 3514 188808 3570 188864
rect 3422 162832 3478 162888
rect 3422 149776 3478 149832
rect 3422 136720 3478 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3422 84632 3478 84688
rect 3514 71576 3570 71632
rect 3054 58520 3110 58576
rect 2778 55800 2834 55856
rect 1398 44784 1454 44840
rect 39302 292848 39358 292904
rect 2870 45500 2872 45520
rect 2872 45500 2924 45520
rect 2924 45500 2926 45520
rect 2870 45464 2926 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 2870 10240 2926 10296
rect 3422 6432 3478 6488
rect 7654 11600 7710 11656
rect 6458 4800 6514 4856
rect 27618 71032 27674 71088
rect 19430 36488 19486 36544
rect 27710 40568 27766 40624
rect 31758 43424 31814 43480
rect 34794 7520 34850 7576
rect 37278 33768 37334 33824
rect 40038 238584 40094 238640
rect 40038 57160 40094 57216
rect 104898 242120 104954 242176
rect 179326 273808 179382 273864
rect 99102 179424 99158 179480
rect 97538 176976 97594 177032
rect 99102 176976 99158 177032
rect 105910 177656 105966 177712
rect 108118 177656 108174 177712
rect 114466 177656 114522 177712
rect 114374 177112 114430 177168
rect 119526 177656 119582 177712
rect 124954 177656 125010 177712
rect 127070 177656 127126 177712
rect 130750 177656 130806 177712
rect 132406 177656 132462 177712
rect 123758 177112 123814 177168
rect 129462 177112 129518 177168
rect 100666 176704 100722 176760
rect 103334 176704 103390 176760
rect 104622 176704 104678 176760
rect 107014 176704 107070 176760
rect 109590 176704 109646 176760
rect 110694 176704 110750 176760
rect 112258 176704 112314 176760
rect 118422 176704 118478 176760
rect 125874 176740 125876 176760
rect 125876 176740 125928 176760
rect 125928 176740 125930 176760
rect 125874 176704 125930 176740
rect 128174 176704 128230 176760
rect 133142 176704 133198 176760
rect 136086 176724 136142 176760
rect 136086 176704 136088 176724
rect 136088 176704 136140 176724
rect 136140 176704 136142 176724
rect 148230 176704 148286 176760
rect 158994 176724 159050 176760
rect 158994 176704 158996 176724
rect 158996 176704 159048 176724
rect 159048 176704 159050 176724
rect 116950 175344 117006 175400
rect 120814 175344 120870 175400
rect 121918 175344 121974 175400
rect 134430 175344 134486 175400
rect 115754 174936 115810 174992
rect 165342 173168 165398 173224
rect 167734 176976 167790 177032
rect 168010 171536 168066 171592
rect 66074 129240 66130 129296
rect 65154 126248 65210 126304
rect 65982 123528 66038 123584
rect 64786 102176 64842 102232
rect 66166 128016 66222 128072
rect 66074 94832 66130 94888
rect 67638 125160 67694 125216
rect 67546 122576 67602 122632
rect 67454 120808 67510 120864
rect 66166 93744 66222 93800
rect 65982 90888 66038 90944
rect 67730 100680 67786 100736
rect 67638 91024 67694 91080
rect 105726 94696 105782 94752
rect 112350 94696 112406 94752
rect 128082 94696 128138 94752
rect 151726 94696 151782 94752
rect 106462 94016 106518 94072
rect 88982 93472 89038 93528
rect 103426 93200 103482 93256
rect 86590 92384 86646 92440
rect 98550 92404 98606 92440
rect 98550 92384 98552 92404
rect 98552 92384 98604 92404
rect 98604 92384 98606 92404
rect 75826 91160 75882 91216
rect 84658 91160 84714 91216
rect 67730 88168 67786 88224
rect 90362 91704 90418 91760
rect 86866 91160 86922 91216
rect 101862 91432 101918 91488
rect 95054 91296 95110 91352
rect 99194 91296 99250 91352
rect 100574 91296 100630 91352
rect 92294 91160 92350 91216
rect 93766 91160 93822 91216
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 97078 91160 97134 91216
rect 97906 91160 97962 91216
rect 99286 91160 99342 91216
rect 99194 82728 99250 82784
rect 100666 91160 100722 91216
rect 101954 91296 102010 91352
rect 102046 91160 102102 91216
rect 103058 91160 103114 91216
rect 101954 81368 102010 81424
rect 121734 93608 121790 93664
rect 111246 93472 111302 93528
rect 110142 93200 110198 93256
rect 104346 92384 104402 92440
rect 104622 92384 104678 92440
rect 106646 92384 106702 92440
rect 106002 91568 106058 91624
rect 109498 91432 109554 91488
rect 108854 91296 108910 91352
rect 108946 91160 109002 91216
rect 110694 92384 110750 92440
rect 118054 92384 118110 92440
rect 134430 93472 134486 93528
rect 126702 92384 126758 92440
rect 133142 92384 133198 92440
rect 151542 92384 151598 92440
rect 115478 91976 115534 92032
rect 126518 91976 126574 92032
rect 151358 91976 151414 92032
rect 114374 91296 114430 91352
rect 110326 91160 110382 91216
rect 113086 91160 113142 91216
rect 114466 91160 114522 91216
rect 119894 91704 119950 91760
rect 117134 91296 117190 91352
rect 115570 91160 115626 91216
rect 115846 91160 115902 91216
rect 115478 89664 115534 89720
rect 117226 91160 117282 91216
rect 113086 81232 113142 81288
rect 118606 91160 118662 91216
rect 70398 72392 70454 72448
rect 42798 46144 42854 46200
rect 44178 22616 44234 22672
rect 45558 17176 45614 17232
rect 62118 51720 62174 51776
rect 77298 47504 77354 47560
rect 124126 91432 124182 91488
rect 120814 91296 120870 91352
rect 121366 91160 121422 91216
rect 123758 91160 123814 91216
rect 124034 91160 124090 91216
rect 125414 91296 125470 91352
rect 125506 91160 125562 91216
rect 132406 91568 132462 91624
rect 126702 91160 126758 91216
rect 129646 91160 129702 91216
rect 130750 91160 130806 91216
rect 126702 86808 126758 86864
rect 136546 91160 136602 91216
rect 130750 85448 130806 85504
rect 152646 91160 152702 91216
rect 167458 110064 167514 110120
rect 167918 111696 167974 111752
rect 167918 108704 167974 108760
rect 179326 181464 179382 181520
rect 171966 93608 172022 93664
rect 182086 178744 182142 178800
rect 186134 178608 186190 178664
rect 190550 240080 190606 240136
rect 190366 177248 190422 177304
rect 103334 10376 103390 10432
rect 124218 62736 124274 62792
rect 192942 239536 192998 239592
rect 193034 182824 193090 182880
rect 191746 175888 191802 175944
rect 196990 272856 197046 272912
rect 197358 291236 197414 291272
rect 197358 291216 197360 291236
rect 197360 291216 197412 291236
rect 197412 291216 197414 291236
rect 197358 290536 197414 290592
rect 197358 289176 197414 289232
rect 197726 288496 197782 288552
rect 197450 287816 197506 287872
rect 197358 287156 197414 287192
rect 197358 287136 197360 287156
rect 197360 287136 197412 287156
rect 197412 287136 197414 287156
rect 197358 286456 197414 286512
rect 198002 285776 198058 285832
rect 197358 285096 197414 285152
rect 197266 284416 197322 284472
rect 197358 280336 197414 280392
rect 197358 279656 197414 279712
rect 197450 278296 197506 278352
rect 197358 277616 197414 277672
rect 197358 276936 197414 276992
rect 197726 276256 197782 276312
rect 197450 275576 197506 275632
rect 197358 274896 197414 274952
rect 197358 274216 197414 274272
rect 197266 272176 197322 272232
rect 197174 248376 197230 248432
rect 197082 239672 197138 239728
rect 195886 185544 195942 185600
rect 197450 271496 197506 271552
rect 197358 270816 197414 270872
rect 197450 270136 197506 270192
rect 197358 269456 197414 269512
rect 197358 268096 197414 268152
rect 197450 267416 197506 267472
rect 197358 266736 197414 266792
rect 197450 266056 197506 266112
rect 197358 265376 197414 265432
rect 197450 264696 197506 264752
rect 197358 264016 197414 264072
rect 197358 263336 197414 263392
rect 197358 262656 197414 262712
rect 197450 261976 197506 262032
rect 197542 261296 197598 261352
rect 197358 260616 197414 260672
rect 197358 259936 197414 259992
rect 197358 259256 197414 259312
rect 197450 258576 197506 258632
rect 197450 257896 197506 257952
rect 197358 257216 197414 257272
rect 197450 255856 197506 255912
rect 197358 255212 197360 255232
rect 197360 255212 197412 255232
rect 197412 255212 197414 255232
rect 197358 255176 197414 255212
rect 197358 254496 197414 254552
rect 197358 253816 197414 253872
rect 197450 252456 197506 252512
rect 197358 251776 197414 251832
rect 198554 283056 198610 283112
rect 198646 281696 198702 281752
rect 198646 281016 198702 281072
rect 198094 273536 198150 273592
rect 198002 252320 198058 252376
rect 198554 251096 198610 251152
rect 197450 250416 197506 250472
rect 197358 249756 197414 249792
rect 197358 249736 197360 249756
rect 197360 249736 197412 249756
rect 197412 249736 197414 249756
rect 197358 249056 197414 249112
rect 197542 247696 197598 247752
rect 197450 247016 197506 247072
rect 197358 245656 197414 245712
rect 197450 244316 197506 244352
rect 197450 244296 197452 244316
rect 197452 244296 197504 244316
rect 197504 244296 197506 244316
rect 197358 243616 197414 243672
rect 197358 242256 197414 242312
rect 200854 295432 200910 295488
rect 201406 292476 201408 292496
rect 201408 292476 201460 292496
rect 201460 292476 201462 292496
rect 201406 292440 201462 292476
rect 211158 296928 211214 296984
rect 209226 293936 209282 293992
rect 216954 298152 217010 298208
rect 220174 299512 220230 299568
rect 229834 294208 229890 294264
rect 236274 293936 236330 293992
rect 235630 292712 235686 292768
rect 238206 296792 238262 296848
rect 243358 295296 243414 295352
rect 242346 292168 242402 292224
rect 244646 294072 244702 294128
rect 244002 292576 244058 292632
rect 248510 292848 248566 292904
rect 249154 292304 249210 292360
rect 200118 291488 200174 291544
rect 249982 287544 250038 287600
rect 200026 278976 200082 279032
rect 249982 269728 250038 269784
rect 200026 268776 200082 268832
rect 199934 256536 199990 256592
rect 199842 253136 199898 253192
rect 199750 244976 199806 245032
rect 199750 239400 199806 239456
rect 200762 240080 200818 240136
rect 198646 193840 198702 193896
rect 204718 190984 204774 191040
rect 205362 186904 205418 186960
rect 197174 177384 197230 177440
rect 207294 197920 207350 197976
rect 207938 184184 207994 184240
rect 206374 181328 206430 181384
rect 209226 180104 209282 180160
rect 213090 228248 213146 228304
rect 209870 179968 209926 180024
rect 213918 175752 213974 175808
rect 213918 175072 213974 175128
rect 214010 174664 214066 174720
rect 213918 173712 213974 173768
rect 214010 173304 214066 173360
rect 214194 172352 214250 172408
rect 214102 171944 214158 172000
rect 213918 170720 213974 170776
rect 214010 170584 214066 170640
rect 213918 169360 213974 169416
rect 214010 169224 214066 169280
rect 213918 168000 213974 168056
rect 214010 167864 214066 167920
rect 213274 166912 213330 166968
rect 213918 166640 213974 166696
rect 214010 166096 214066 166152
rect 213918 164736 213974 164792
rect 214470 164092 214472 164112
rect 214472 164092 214524 164112
rect 214524 164092 214526 164112
rect 214470 164056 214526 164092
rect 213918 163376 213974 163432
rect 213918 162560 213974 162616
rect 213182 162016 213238 162072
rect 213918 161372 213920 161392
rect 213920 161372 213972 161392
rect 213972 161372 213974 161392
rect 213918 161336 213974 161372
rect 213918 160012 213920 160032
rect 213920 160012 213972 160032
rect 213972 160012 213974 160032
rect 213918 159976 213974 160012
rect 214010 159432 214066 159488
rect 213918 158652 213920 158672
rect 213920 158652 213972 158672
rect 213972 158652 213974 158672
rect 213918 158616 213974 158652
rect 214102 158072 214158 158128
rect 213918 156848 213974 156904
rect 213918 155488 213974 155544
rect 214010 153856 214066 153912
rect 213918 153332 213974 153368
rect 213918 153312 213920 153332
rect 213920 153312 213972 153332
rect 213972 153312 213974 153332
rect 214010 152632 214066 152688
rect 213918 151952 213974 152008
rect 214010 150728 214066 150784
rect 213918 150592 213974 150648
rect 214654 165452 214656 165472
rect 214656 165452 214708 165472
rect 214708 165452 214710 165472
rect 214654 165416 214710 165452
rect 214562 150184 214618 150240
rect 213918 149504 213974 149560
rect 215022 151816 215078 151872
rect 214746 148824 214802 148880
rect 213918 148008 213974 148064
rect 213918 146648 213974 146704
rect 214562 146376 214618 146432
rect 213918 145288 213974 145344
rect 214010 143928 214066 143984
rect 213918 143556 213920 143576
rect 213920 143556 213972 143576
rect 213972 143556 213974 143576
rect 213918 143520 213974 143556
rect 213918 142704 213974 142760
rect 214010 141344 214066 141400
rect 213918 140936 213974 140992
rect 213918 139460 213974 139496
rect 213918 139440 213920 139460
rect 213920 139440 213972 139460
rect 213972 139440 213974 139460
rect 204994 94832 205050 94888
rect 214010 138760 214066 138816
rect 213918 138100 213974 138136
rect 213918 138080 213920 138100
rect 213920 138080 213972 138100
rect 213972 138080 213974 138100
rect 213918 137400 213974 137456
rect 213182 136040 213238 136096
rect 213918 134000 213974 134056
rect 214010 132776 214066 132832
rect 213918 132540 213920 132560
rect 213920 132540 213972 132560
rect 213972 132540 213974 132560
rect 213918 132504 213974 132540
rect 214010 131416 214066 131472
rect 213918 131180 213920 131200
rect 213920 131180 213972 131200
rect 213972 131180 213974 131200
rect 213918 131144 213974 131180
rect 214010 130056 214066 130112
rect 213918 129804 213974 129840
rect 213918 129784 213920 129804
rect 213920 129784 213972 129804
rect 213972 129784 213974 129804
rect 213918 128424 213974 128480
rect 213918 127064 213974 127120
rect 214010 126112 214066 126168
rect 213918 125704 213974 125760
rect 214010 124752 214066 124808
rect 213918 124344 213974 124400
rect 214010 123528 214066 123584
rect 213918 123120 213974 123176
rect 213918 122168 213974 122224
rect 214470 121624 214526 121680
rect 214010 120808 214066 120864
rect 213918 120400 213974 120456
rect 214010 119584 214066 119640
rect 213274 119040 213330 119096
rect 213918 118904 213974 118960
rect 214010 117544 214066 117600
rect 213918 117308 213920 117328
rect 213920 117308 213972 117328
rect 213972 117308 213974 117328
rect 213918 117272 213974 117308
rect 213918 116184 213974 116240
rect 213366 115912 213422 115968
rect 214010 114960 214066 115016
rect 213918 114572 213974 114608
rect 213918 114552 213920 114572
rect 213920 114552 213972 114572
rect 213972 114552 213974 114572
rect 214010 113600 214066 113656
rect 213918 113228 213920 113248
rect 213920 113228 213972 113248
rect 213972 113228 213974 113248
rect 213918 113192 213974 113228
rect 214010 112240 214066 112296
rect 213918 111852 213974 111888
rect 213918 111832 213920 111852
rect 213920 111832 213972 111852
rect 213972 111832 213974 111852
rect 214010 110880 214066 110936
rect 213918 110508 213920 110528
rect 213920 110508 213972 110528
rect 213972 110508 213974 110528
rect 213918 110472 213974 110508
rect 214010 109656 214066 109712
rect 213918 109132 213974 109168
rect 213918 109112 213920 109132
rect 213920 109112 213972 109132
rect 213972 109112 213974 109132
rect 214010 108296 214066 108352
rect 213918 107888 213974 107944
rect 214010 106936 214066 106992
rect 213918 106528 213974 106584
rect 214010 105712 214066 105768
rect 213918 105304 213974 105360
rect 213458 105168 213514 105224
rect 213918 103672 213974 103728
rect 214746 135496 214802 135552
rect 214654 134136 214710 134192
rect 214010 101224 214066 101280
rect 213918 101088 213974 101144
rect 213918 99728 213974 99784
rect 214102 99456 214158 99512
rect 214010 98368 214066 98424
rect 213918 97960 213974 98016
rect 213918 97008 213974 97064
rect 214102 95784 214158 95840
rect 214562 95784 214618 95840
rect 213458 93744 213514 93800
rect 214746 108432 214802 108488
rect 214746 102448 214802 102504
rect 214838 96600 214894 96656
rect 219530 238448 219586 238504
rect 225970 238584 226026 238640
rect 227626 175752 227682 175808
rect 229190 168952 229246 169008
rect 229098 154264 229154 154320
rect 231766 175208 231822 175264
rect 231122 174664 231178 174720
rect 231674 173732 231730 173768
rect 231674 173712 231676 173732
rect 231676 173712 231728 173732
rect 231728 173712 231730 173732
rect 231214 173304 231270 173360
rect 231766 172760 231822 172816
rect 231766 172352 231822 172408
rect 231674 171808 231730 171864
rect 231674 171400 231730 171456
rect 230662 164328 230718 164384
rect 230662 158616 230718 158672
rect 230754 157664 230810 157720
rect 231766 170856 231822 170912
rect 231766 170484 231768 170504
rect 231768 170484 231820 170504
rect 231820 170484 231822 170504
rect 231766 170448 231822 170484
rect 231306 169904 231362 169960
rect 231674 169532 231676 169552
rect 231676 169532 231728 169552
rect 231728 169532 231730 169552
rect 231674 169496 231730 169532
rect 231766 168544 231822 168600
rect 231766 168000 231822 168056
rect 231674 167592 231730 167648
rect 231582 167048 231638 167104
rect 231766 166640 231822 166696
rect 231122 166096 231178 166152
rect 231490 165688 231546 165744
rect 231766 165144 231822 165200
rect 231306 164736 231362 164792
rect 231674 162832 231730 162888
rect 231766 162424 231822 162480
rect 231766 161880 231822 161936
rect 231674 161472 231730 161528
rect 231766 160928 231822 160984
rect 231398 160520 231454 160576
rect 231766 159568 231822 159624
rect 231490 159024 231546 159080
rect 231766 158072 231822 158128
rect 231766 157120 231822 157176
rect 231674 156712 231730 156768
rect 230938 156168 230994 156224
rect 231122 155796 231124 155816
rect 231124 155796 231176 155816
rect 231176 155796 231178 155816
rect 231122 155760 231178 155796
rect 230570 155216 230626 155272
rect 231582 155216 231638 155272
rect 231766 154808 231822 154864
rect 231766 152904 231822 152960
rect 231674 152496 231730 152552
rect 231582 151952 231638 152008
rect 231674 151544 231730 151600
rect 231766 151000 231822 151056
rect 231766 150592 231822 150648
rect 231950 153312 232006 153368
rect 230938 149640 230994 149696
rect 230478 147736 230534 147792
rect 230938 146784 230994 146840
rect 231030 145288 231086 145344
rect 214838 88168 214894 88224
rect 231122 142432 231178 142488
rect 231766 150048 231822 150104
rect 231674 149096 231730 149152
rect 231766 148144 231822 148200
rect 231766 147192 231822 147248
rect 231766 146260 231822 146296
rect 231766 146240 231768 146260
rect 231768 146240 231820 146260
rect 231820 146240 231822 146260
rect 231674 145832 231730 145888
rect 231766 145560 231822 145616
rect 231766 144336 231822 144392
rect 231582 143928 231638 143984
rect 231766 143420 231768 143440
rect 231768 143420 231820 143440
rect 231820 143420 231822 143440
rect 231766 143384 231822 143420
rect 231674 142976 231730 143032
rect 231030 134000 231086 134056
rect 230938 133048 230994 133104
rect 231122 126384 231178 126440
rect 231030 125976 231086 126032
rect 230662 118360 230718 118416
rect 230662 117000 230718 117056
rect 230570 116492 230572 116512
rect 230572 116492 230624 116512
rect 230624 116492 230626 116512
rect 230570 116456 230626 116492
rect 231766 141072 231822 141128
rect 231766 140684 231822 140720
rect 231766 140664 231768 140684
rect 231768 140664 231820 140684
rect 231820 140664 231822 140684
rect 231674 140120 231730 140176
rect 231398 137264 231454 137320
rect 231398 135904 231454 135960
rect 231490 134408 231546 134464
rect 231766 136856 231822 136912
rect 231766 135360 231822 135416
rect 231582 133456 231638 133512
rect 231674 132504 231730 132560
rect 231306 131552 231362 131608
rect 231766 132096 231822 132152
rect 231674 131144 231730 131200
rect 231398 130192 231454 130248
rect 231306 129240 231362 129296
rect 231766 130600 231822 130656
rect 231674 129784 231730 129840
rect 231490 128832 231546 128888
rect 231306 124480 231362 124536
rect 230846 121624 230902 121680
rect 230938 120672 230994 120728
rect 231766 128288 231822 128344
rect 231674 127880 231730 127936
rect 231674 127336 231730 127392
rect 231766 126928 231822 126984
rect 231766 125024 231822 125080
rect 231582 124072 231638 124128
rect 231582 123564 231584 123584
rect 231584 123564 231636 123584
rect 231636 123564 231638 123584
rect 231582 123528 231638 123564
rect 231766 123120 231822 123176
rect 231490 122576 231546 122632
rect 231306 122168 231362 122224
rect 231122 120264 231178 120320
rect 230938 119720 230994 119776
rect 230938 117408 230994 117464
rect 231490 118904 231546 118960
rect 230754 116048 230810 116104
rect 230662 114144 230718 114200
rect 230570 113192 230626 113248
rect 231490 113600 231546 113656
rect 230938 112648 230994 112704
rect 230570 106528 230626 106584
rect 229926 101768 229982 101824
rect 230846 105168 230902 105224
rect 230570 100816 230626 100872
rect 231122 109792 231178 109848
rect 231122 108432 231178 108488
rect 231030 103672 231086 103728
rect 231766 121216 231822 121272
rect 231766 119312 231822 119368
rect 231766 117952 231822 118008
rect 231766 115504 231822 115560
rect 231766 115132 231768 115152
rect 231768 115132 231820 115152
rect 231820 115132 231822 115152
rect 231766 115096 231822 115132
rect 231674 114552 231730 114608
rect 231674 112240 231730 112296
rect 231766 111732 231768 111752
rect 231768 111732 231820 111752
rect 231820 111732 231822 111752
rect 231766 111696 231822 111732
rect 231674 111288 231730 111344
rect 231582 110744 231638 110800
rect 231490 109384 231546 109440
rect 231766 110372 231768 110392
rect 231768 110372 231820 110392
rect 231820 110372 231822 110392
rect 231766 110336 231822 110372
rect 231766 108876 231768 108896
rect 231768 108876 231820 108896
rect 231820 108876 231822 108896
rect 231766 108840 231822 108876
rect 231674 107888 231730 107944
rect 234986 181464 235042 181520
rect 233790 151000 233846 151056
rect 231766 107480 231822 107536
rect 231582 107072 231638 107128
rect 231306 102312 231362 102368
rect 231122 101360 231178 101416
rect 231674 106156 231676 106176
rect 231676 106156 231728 106176
rect 231728 106156 231730 106176
rect 231674 106120 231730 106156
rect 231766 105576 231822 105632
rect 231582 104660 231584 104680
rect 231584 104660 231636 104680
rect 231636 104660 231638 104680
rect 231582 104624 231638 104660
rect 231766 104216 231822 104272
rect 231582 103300 231584 103320
rect 231584 103300 231636 103320
rect 231636 103300 231638 103320
rect 231582 103264 231638 103300
rect 231766 102720 231822 102776
rect 231766 100408 231822 100464
rect 231674 99864 231730 99920
rect 231398 99456 231454 99512
rect 230662 98912 230718 98968
rect 231490 98504 231546 98560
rect 230478 97552 230534 97608
rect 230478 97008 230534 97064
rect 231122 96600 231178 96656
rect 230478 95648 230534 95704
rect 238758 239672 238814 239728
rect 238022 135224 238078 135280
rect 241426 153176 241482 153232
rect 248518 239944 248574 240000
rect 249154 238584 249210 238640
rect 250074 253408 250130 253464
rect 250442 281968 250498 282024
rect 250350 258848 250406 258904
rect 250258 240352 250314 240408
rect 251270 286456 251326 286512
rect 251270 273536 251326 273592
rect 251178 261296 251234 261352
rect 251178 257896 251234 257952
rect 251086 240488 251142 240544
rect 252558 291896 252614 291952
rect 252926 289176 252982 289232
rect 252558 280356 252614 280392
rect 252558 280336 252560 280356
rect 252560 280336 252612 280356
rect 252612 280336 252614 280356
rect 252006 278976 252062 279032
rect 251362 271496 251418 271552
rect 252650 274252 252652 274272
rect 252652 274252 252704 274272
rect 252704 274252 252706 274272
rect 252650 274216 252706 274252
rect 253294 283736 253350 283792
rect 253754 291216 253810 291272
rect 253754 289856 253810 289912
rect 253754 288516 253810 288552
rect 253754 288496 253756 288516
rect 253756 288496 253808 288516
rect 253808 288496 253810 288516
rect 253754 287816 253810 287872
rect 253754 285776 253810 285832
rect 253846 284416 253902 284472
rect 253754 283056 253810 283112
rect 253754 281016 253810 281072
rect 253754 278296 253810 278352
rect 253294 276936 253350 276992
rect 253478 276256 253534 276312
rect 253294 275576 253350 275632
rect 253202 272856 253258 272912
rect 253846 277616 253902 277672
rect 252650 272196 252706 272232
rect 252650 272176 252652 272196
rect 252652 272176 252704 272196
rect 252704 272176 252706 272196
rect 252650 268776 252706 268832
rect 253202 268096 253258 268152
rect 253294 267416 253350 267472
rect 253754 266736 253810 266792
rect 253846 266056 253902 266112
rect 253754 265376 253810 265432
rect 253754 264696 253810 264752
rect 252742 264016 252798 264072
rect 252558 263336 252614 263392
rect 252558 258576 252614 258632
rect 253754 262656 253810 262712
rect 253386 261976 253442 262032
rect 252834 260616 252890 260672
rect 253202 259936 253258 259992
rect 252742 250416 252798 250472
rect 252650 248376 252706 248432
rect 252558 241596 252614 241632
rect 252558 241576 252560 241596
rect 252560 241576 252612 241596
rect 252612 241576 252614 241596
rect 253018 257216 253074 257272
rect 253754 256572 253756 256592
rect 253756 256572 253808 256592
rect 253808 256572 253810 256592
rect 253754 256536 253810 256572
rect 253110 255856 253166 255912
rect 253754 255176 253810 255232
rect 253018 254496 253074 254552
rect 253846 253136 253902 253192
rect 253754 252492 253756 252512
rect 253756 252492 253808 252512
rect 253808 252492 253810 252512
rect 253754 252456 253810 252492
rect 253478 251776 253534 251832
rect 253386 251096 253442 251152
rect 253754 249756 253810 249792
rect 253754 249736 253756 249756
rect 253756 249736 253808 249756
rect 253808 249736 253810 249756
rect 253754 249056 253810 249112
rect 253846 247696 253902 247752
rect 253754 247052 253756 247072
rect 253756 247052 253808 247072
rect 253808 247052 253810 247072
rect 253754 247016 253810 247052
rect 253754 245676 253810 245712
rect 253754 245656 253756 245676
rect 253756 245656 253808 245676
rect 253808 245656 253810 245676
rect 253846 244976 253902 245032
rect 253754 244316 253810 244352
rect 253754 244296 253756 244316
rect 253756 244296 253808 244316
rect 253808 244296 253810 244316
rect 253754 243616 253810 243672
rect 253386 242936 253442 242992
rect 253754 242256 253810 242312
rect 253754 240216 253810 240272
rect 254122 290536 254178 290592
rect 257342 292712 257398 292768
rect 256882 240352 256938 240408
rect 258170 235184 258226 235240
rect 261390 166776 261446 166832
rect 261666 157256 261722 157312
rect 262402 268368 262458 268424
rect 261574 146104 261630 146160
rect 261482 144064 261538 144120
rect 260470 140120 260526 140176
rect 260470 139712 260526 139768
rect 261666 119856 261722 119912
rect 262862 239944 262918 240000
rect 265806 175344 265862 175400
rect 265346 174936 265402 174992
rect 265806 174528 265862 174584
rect 265622 174120 265678 174176
rect 265898 173984 265954 174040
rect 265714 173168 265770 173224
rect 265346 171944 265402 172000
rect 265346 170584 265402 170640
rect 264242 170176 264298 170232
rect 265898 172760 265954 172816
rect 265806 172524 265808 172544
rect 265808 172524 265860 172544
rect 265860 172524 265862 172544
rect 265806 172488 265862 172524
rect 265806 171536 265862 171592
rect 265898 171164 265900 171184
rect 265900 171164 265952 171184
rect 265952 171164 265954 171184
rect 265898 171128 265954 171164
rect 265622 169768 265678 169824
rect 265438 169360 265494 169416
rect 265346 168952 265402 169008
rect 264426 168136 264482 168192
rect 265162 167592 265218 167648
rect 265806 168544 265862 168600
rect 265806 167184 265862 167240
rect 265990 166368 266046 166424
rect 265714 165960 265770 166016
rect 265806 165708 265862 165744
rect 265806 165688 265808 165708
rect 265808 165688 265860 165708
rect 265860 165688 265862 165708
rect 265438 165008 265494 165064
rect 265714 164600 265770 164656
rect 265530 163376 265586 163432
rect 265346 162988 265402 163024
rect 265346 162968 265348 162988
rect 265348 162968 265400 162988
rect 265400 162968 265402 162988
rect 265346 162016 265402 162072
rect 265346 160792 265402 160848
rect 265622 160384 265678 160440
rect 265346 159432 265402 159488
rect 265622 159024 265678 159080
rect 265622 158208 265678 158264
rect 265254 157800 265310 157856
rect 265530 157412 265586 157448
rect 265530 157392 265532 157412
rect 265532 157392 265584 157412
rect 265584 157392 265586 157412
rect 265806 164192 265862 164248
rect 265898 163784 265954 163840
rect 265806 162832 265862 162888
rect 265806 161608 265862 161664
rect 265806 160132 265862 160168
rect 265806 160112 265808 160132
rect 265808 160112 265860 160132
rect 265860 160112 265862 160132
rect 265806 158772 265862 158808
rect 265806 158752 265808 158772
rect 265808 158752 265860 158772
rect 265860 158752 265862 158772
rect 265530 156440 265586 156496
rect 264426 152088 264482 152144
rect 264334 141888 264390 141944
rect 264334 123800 264390 123856
rect 264242 107480 264298 107536
rect 265346 150048 265402 150104
rect 265438 148688 265494 148744
rect 265162 148280 265218 148336
rect 265530 147056 265586 147112
rect 264518 145696 264574 145752
rect 265530 144880 265586 144936
rect 265438 144472 265494 144528
rect 265898 156848 265954 156904
rect 265806 156032 265862 156088
rect 265806 155624 265862 155680
rect 265714 155216 265770 155272
rect 265990 154672 266046 154728
rect 265898 153856 265954 153912
rect 265806 153448 265862 153504
rect 265898 153176 265954 153232
rect 265714 152632 265770 152688
rect 265806 151836 265862 151872
rect 265806 151816 265808 151836
rect 265808 151816 265860 151836
rect 265860 151816 265862 151836
rect 266082 154536 266138 154592
rect 265990 151272 266046 151328
rect 265898 150864 265954 150920
rect 265806 150476 265862 150512
rect 265806 150456 265808 150476
rect 265808 150456 265860 150476
rect 265860 150456 265862 150476
rect 265898 149640 265954 149696
rect 265806 149232 265862 149288
rect 265806 147872 265862 147928
rect 265806 146648 265862 146704
rect 266082 146512 266138 146568
rect 265806 145288 265862 145344
rect 265806 143928 265862 143984
rect 265898 143520 265954 143576
rect 265714 143112 265770 143168
rect 265346 142704 265402 142760
rect 264610 142296 264666 142352
rect 264518 115912 264574 115968
rect 264518 110064 264574 110120
rect 264426 104488 264482 104544
rect 265438 139460 265494 139496
rect 265438 139440 265440 139460
rect 265440 139440 265492 139460
rect 265492 139440 265494 139460
rect 265438 138760 265494 138816
rect 265162 138352 265218 138408
rect 265622 138116 265624 138136
rect 265624 138116 265676 138136
rect 265676 138116 265678 138136
rect 265622 138080 265678 138116
rect 265622 137536 265678 137592
rect 265530 136740 265586 136776
rect 265530 136720 265532 136740
rect 265532 136720 265584 136740
rect 265584 136720 265586 136740
rect 265622 136312 265678 136368
rect 265346 135904 265402 135960
rect 265530 134544 265586 134600
rect 265622 132776 265678 132832
rect 265162 131552 265218 131608
rect 265622 131180 265624 131200
rect 265624 131180 265676 131200
rect 265676 131180 265678 131200
rect 265622 131144 265678 131180
rect 265530 130600 265586 130656
rect 265622 128968 265678 129024
rect 265346 127608 265402 127664
rect 265254 125976 265310 126032
rect 265530 124616 265586 124672
rect 265530 123392 265586 123448
rect 265070 123004 265126 123040
rect 265070 122984 265072 123004
rect 265072 122984 265124 123004
rect 265124 122984 265126 123004
rect 265254 119040 265310 119096
rect 265530 118224 265586 118280
rect 265162 117816 265218 117872
rect 265254 114824 265310 114880
rect 265254 113464 265310 113520
rect 265438 113212 265494 113248
rect 265438 113192 265440 113212
rect 265440 113192 265492 113212
rect 265492 113192 265494 113212
rect 265530 112648 265586 112704
rect 265530 111288 265586 111344
rect 265162 110880 265218 110936
rect 265530 109656 265586 109712
rect 265438 108296 265494 108352
rect 265346 107908 265402 107944
rect 265346 107888 265348 107908
rect 265348 107888 265400 107908
rect 265400 107888 265402 107908
rect 265530 107072 265586 107128
rect 265530 101904 265586 101960
rect 265530 99456 265586 99512
rect 265438 97996 265440 98016
rect 265440 97996 265492 98016
rect 265492 97996 265494 98016
rect 265438 97960 265494 97996
rect 265162 97144 265218 97200
rect 265806 140936 265862 140992
rect 265990 141344 266046 141400
rect 265714 119448 265770 119504
rect 265714 117408 265770 117464
rect 265714 113872 265770 113928
rect 265714 112240 265770 112296
rect 265714 110492 265770 110528
rect 265714 110472 265716 110492
rect 265716 110472 265768 110492
rect 265768 110472 265770 110492
rect 265714 109248 265770 109304
rect 265714 108704 265770 108760
rect 265898 135360 265954 135416
rect 265898 134136 265954 134192
rect 265898 133900 265900 133920
rect 265900 133900 265952 133920
rect 265952 133900 265954 133920
rect 265898 133864 265954 133900
rect 265898 132524 265954 132560
rect 265898 132504 265900 132524
rect 265900 132504 265952 132524
rect 265952 132504 265954 132524
rect 265898 131960 265954 132016
rect 265898 129376 265954 129432
rect 265898 127200 265954 127256
rect 265898 126384 265954 126440
rect 266082 135768 266138 135824
rect 266174 125568 266230 125624
rect 265898 125024 265954 125080
rect 265990 124208 266046 124264
rect 265990 122032 266046 122088
rect 265898 121624 265954 121680
rect 265990 120808 266046 120864
rect 265898 120148 265954 120184
rect 265898 120128 265900 120148
rect 265900 120128 265952 120148
rect 265952 120128 265954 120148
rect 266266 122848 266322 122904
rect 265806 106664 265862 106720
rect 265714 106528 265770 106584
rect 265714 105712 265770 105768
rect 265806 105304 265862 105360
rect 265806 103556 265862 103592
rect 265806 103536 265808 103556
rect 265808 103536 265860 103556
rect 265860 103536 265862 103556
rect 265714 103128 265770 103184
rect 265806 102312 265862 102368
rect 265714 101496 265770 101552
rect 265806 100952 265862 101008
rect 265714 100136 265770 100192
rect 265806 99728 265862 99784
rect 265806 98368 265862 98424
rect 265806 97552 265862 97608
rect 265806 96328 265862 96384
rect 266174 116864 266230 116920
rect 266082 116456 266138 116512
rect 266082 112104 266138 112160
rect 266082 104896 266138 104952
rect 266082 103944 266138 104000
rect 267186 95920 267242 95976
rect 300122 697448 300178 697504
rect 269854 177384 269910 177440
rect 279422 177520 279478 177576
rect 273994 175888 274050 175944
rect 269762 175752 269818 175808
rect 279422 174392 279478 174448
rect 279330 173712 279386 173768
rect 282918 295432 282974 295488
rect 281538 236544 281594 236600
rect 280802 191120 280858 191176
rect 280342 172352 280398 172408
rect 282826 170856 282882 170912
rect 282734 170040 282790 170096
rect 282826 169360 282882 169416
rect 281722 168544 281778 168600
rect 281630 167728 281686 167784
rect 282458 167048 282514 167104
rect 282090 166232 282146 166288
rect 282826 165452 282828 165472
rect 282828 165452 282880 165472
rect 282880 165452 282882 165472
rect 282826 165416 282882 165452
rect 281998 164736 282054 164792
rect 282090 163920 282146 163976
rect 282826 163104 282882 163160
rect 282090 162424 282146 162480
rect 282826 161608 282882 161664
rect 281538 160112 281594 160168
rect 281538 159296 281594 159352
rect 282826 160792 282882 160848
rect 282826 158480 282882 158536
rect 282734 157800 282790 157856
rect 281722 156304 281778 156360
rect 281630 154672 281686 154728
rect 281722 153992 281778 154048
rect 282826 153176 282882 153232
rect 282734 152360 282790 152416
rect 280250 151680 280306 151736
rect 282826 150864 282882 150920
rect 282826 150048 282882 150104
rect 281538 149368 281594 149424
rect 282826 148552 282882 148608
rect 282274 147736 282330 147792
rect 281722 147056 281778 147112
rect 282826 146240 282882 146296
rect 281998 145424 282054 145480
rect 282550 144780 282552 144800
rect 282552 144780 282604 144800
rect 282604 144780 282606 144800
rect 282550 144744 282606 144780
rect 282826 143928 282882 143984
rect 281630 142432 281686 142488
rect 282826 141616 282882 141672
rect 281906 140120 281962 140176
rect 282826 139340 282828 139360
rect 282828 139340 282880 139360
rect 282880 139340 282882 139360
rect 282826 139304 282882 139340
rect 282734 138488 282790 138544
rect 282826 137844 282828 137864
rect 282828 137844 282880 137864
rect 282880 137844 282882 137864
rect 282826 137808 282882 137844
rect 282182 136992 282238 137048
rect 280158 136312 280214 136368
rect 282826 134000 282882 134056
rect 285678 292304 285734 292360
rect 282826 133184 282882 133240
rect 283194 177248 283250 177304
rect 283102 155488 283158 155544
rect 282826 132404 282828 132424
rect 282828 132404 282880 132424
rect 282880 132404 282882 132424
rect 282826 132368 282882 132404
rect 282826 130872 282882 130928
rect 282274 130056 282330 130112
rect 282826 128560 282882 128616
rect 281722 127744 281778 127800
rect 282826 126248 282882 126304
rect 282826 125432 282882 125488
rect 282090 124752 282146 124808
rect 282826 123936 282882 123992
rect 282734 123120 282790 123176
rect 282090 122440 282146 122496
rect 281722 120808 281778 120864
rect 282458 120128 282514 120184
rect 282090 119312 282146 119368
rect 282826 118496 282882 118552
rect 282734 117816 282790 117872
rect 282826 117000 282882 117056
rect 282734 116320 282790 116376
rect 282090 115504 282146 115560
rect 281722 114688 281778 114744
rect 282826 114008 282882 114064
rect 282090 112376 282146 112432
rect 282826 111732 282828 111752
rect 282828 111732 282880 111752
rect 282880 111732 282882 111752
rect 282826 111696 282882 111732
rect 280158 110880 280214 110936
rect 279422 98096 279478 98152
rect 279330 96600 279386 96656
rect 279330 95920 279386 95976
rect 279514 97280 279570 97336
rect 279422 95104 279478 95160
rect 280066 95784 280122 95840
rect 282826 108568 282882 108624
rect 294234 178608 294290 178664
rect 296626 171128 296682 171184
rect 281538 107752 281594 107808
rect 298374 179968 298430 180024
rect 280250 107072 280306 107128
rect 280066 93608 280122 93664
rect 282458 106256 282514 106312
rect 282826 105440 282882 105496
rect 282458 104896 282514 104952
rect 280342 104760 280398 104816
rect 282826 103128 282882 103184
rect 282458 102448 282514 102504
rect 281630 101632 281686 101688
rect 281538 100136 281594 100192
rect 281814 100816 281870 100872
rect 280250 93472 280306 93528
rect 282826 99340 282882 99376
rect 282826 99320 282828 99340
rect 282828 99320 282880 99340
rect 282880 99320 282882 99340
rect 313278 292168 313334 292224
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 582378 617480 582434 617536
rect 579802 564304 579858 564360
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 272176 580226 272232
rect 579618 258848 579674 258904
rect 579894 245520 579950 245576
rect 580170 232328 580226 232384
rect 579894 205672 579950 205728
rect 580170 192480 580226 192536
rect 580170 165824 580226 165880
rect 579802 152632 579858 152688
rect 582470 590960 582526 591016
rect 582562 537784 582618 537840
rect 582930 365064 582986 365120
rect 582746 295296 582802 295352
rect 582654 293936 582710 293992
rect 582378 182824 582434 182880
rect 580354 179152 580410 179208
rect 580262 139304 580318 139360
rect 580170 125976 580226 126032
rect 580170 99456 580226 99512
rect 582378 86128 582434 86184
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 583114 298696 583170 298752
rect 583022 219000 583078 219056
rect 582838 112784 582894 112840
rect 582746 72936 582802 72992
rect 582654 19760 582710 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 191598 697444 191604 697508
rect 191668 697506 191674 697508
rect 300117 697506 300183 697509
rect 191668 697504 300183 697506
rect 191668 697448 300122 697504
rect 300178 697448 300183 697504
rect 191668 697446 300183 697448
rect 191668 697444 191674 697446
rect 300117 697443 300183 697446
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 582373 617538 582439 617541
rect 583520 617538 584960 617628
rect 582373 617536 584960 617538
rect 582373 617480 582378 617536
rect 582434 617480 584960 617536
rect 582373 617478 584960 617480
rect 582373 617475 582439 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 582465 591018 582531 591021
rect 583520 591018 584960 591108
rect 582465 591016 584960 591018
rect 582465 590960 582470 591016
rect 582526 590960 584960 591016
rect 582465 590958 584960 590960
rect 582465 590955 582531 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 583520 577690 584960 577780
rect 583342 577630 584960 577690
rect 583342 577554 583402 577630
rect 583520 577554 584960 577630
rect 583342 577540 584960 577554
rect 583342 577494 583586 577540
rect 255814 576812 255820 576876
rect 255884 576874 255890 576876
rect 583526 576874 583586 577494
rect 255884 576814 583586 576874
rect 255884 576812 255890 576814
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 582557 537842 582623 537845
rect 583520 537842 584960 537932
rect 582557 537840 584960 537842
rect 582557 537784 582562 537840
rect 582618 537784 584960 537840
rect 582557 537782 584960 537784
rect 582557 537779 582623 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 583520 458146 584960 458236
rect 583342 458086 584960 458146
rect 583342 458010 583402 458086
rect 583520 458010 584960 458086
rect 583342 457996 584960 458010
rect 583342 457950 583586 457996
rect 187550 456860 187556 456924
rect 187620 456922 187626 456924
rect 583526 456922 583586 457950
rect 187620 456862 583586 456922
rect 187620 456860 187626 456862
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 190494 397490 190500 397492
rect -960 397430 190500 397490
rect -960 397340 480 397430
rect 190494 397428 190500 397430
rect 190564 397428 190570 397492
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 582925 365122 582991 365125
rect 583520 365122 584960 365212
rect 582925 365120 584960 365122
rect 582925 365064 582930 365120
rect 582986 365064 584960 365120
rect 582925 365062 584960 365064
rect 582925 365059 582991 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 220169 299570 220235 299573
rect 291142 299570 291148 299572
rect 220169 299568 291148 299570
rect 220169 299512 220174 299568
rect 220230 299512 291148 299568
rect 220169 299510 291148 299512
rect 220169 299507 220235 299510
rect 291142 299508 291148 299510
rect 291212 299508 291218 299572
rect 583109 298754 583175 298757
rect 583520 298754 584960 298844
rect 583109 298752 584960 298754
rect 583109 298696 583114 298752
rect 583170 298696 584960 298752
rect 583109 298694 584960 298696
rect 583109 298691 583175 298694
rect 583520 298604 584960 298694
rect 216949 298210 217015 298213
rect 295558 298210 295564 298212
rect 216949 298208 295564 298210
rect 216949 298152 216954 298208
rect 217010 298152 295564 298208
rect 216949 298150 295564 298152
rect 216949 298147 217015 298150
rect 295558 298148 295564 298150
rect 295628 298148 295634 298212
rect 211153 296986 211219 296989
rect 258390 296986 258396 296988
rect 211153 296984 258396 296986
rect 211153 296928 211158 296984
rect 211214 296928 258396 296984
rect 211153 296926 258396 296928
rect 211153 296923 211219 296926
rect 258390 296924 258396 296926
rect 258460 296924 258466 296988
rect 238201 296850 238267 296853
rect 295374 296850 295380 296852
rect 238201 296848 295380 296850
rect 238201 296792 238206 296848
rect 238262 296792 295380 296848
rect 238201 296790 295380 296792
rect 238201 296787 238267 296790
rect 295374 296788 295380 296790
rect 295444 296788 295450 296852
rect 200849 295490 200915 295493
rect 282913 295490 282979 295493
rect 200849 295488 282979 295490
rect 200849 295432 200854 295488
rect 200910 295432 282918 295488
rect 282974 295432 282979 295488
rect 200849 295430 282979 295432
rect 200849 295427 200915 295430
rect 282913 295427 282979 295430
rect 243353 295354 243419 295357
rect 582741 295354 582807 295357
rect 243353 295352 582807 295354
rect 243353 295296 243358 295352
rect 243414 295296 582746 295352
rect 582802 295296 582807 295352
rect 243353 295294 582807 295296
rect 243353 295291 243419 295294
rect 582741 295291 582807 295294
rect 229829 294266 229895 294269
rect 249006 294266 249012 294268
rect 229829 294264 249012 294266
rect 229829 294208 229834 294264
rect 229890 294208 249012 294264
rect 229829 294206 249012 294208
rect 229829 294203 229895 294206
rect 249006 294204 249012 294206
rect 249076 294204 249082 294268
rect 244641 294130 244707 294133
rect 288382 294130 288388 294132
rect 244641 294128 288388 294130
rect 244641 294072 244646 294128
rect 244702 294072 288388 294128
rect 244641 294070 288388 294072
rect 244641 294067 244707 294070
rect 288382 294068 288388 294070
rect 288452 294068 288458 294132
rect 200246 293932 200252 293996
rect 200316 293994 200322 293996
rect 209221 293994 209287 293997
rect 200316 293992 209287 293994
rect 200316 293936 209226 293992
rect 209282 293936 209287 293992
rect 200316 293934 209287 293936
rect 200316 293932 200322 293934
rect 209221 293931 209287 293934
rect 236269 293994 236335 293997
rect 582649 293994 582715 293997
rect 236269 293992 582715 293994
rect 236269 293936 236274 293992
rect 236330 293936 582654 293992
rect 582710 293936 582715 293992
rect 236269 293934 582715 293936
rect 236269 293931 236335 293934
rect 582649 293931 582715 293934
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 39297 292906 39363 292909
rect 248505 292906 248571 292909
rect 39297 292904 248571 292906
rect 39297 292848 39302 292904
rect 39358 292848 248510 292904
rect 248566 292848 248571 292904
rect 39297 292846 248571 292848
rect 39297 292843 39363 292846
rect 248505 292843 248571 292846
rect 235625 292770 235691 292773
rect 257337 292770 257403 292773
rect 235625 292768 257403 292770
rect 235625 292712 235630 292768
rect 235686 292712 257342 292768
rect 257398 292712 257403 292768
rect 235625 292710 257403 292712
rect 235625 292707 235691 292710
rect 257337 292707 257403 292710
rect 243997 292634 244063 292637
rect 288566 292634 288572 292636
rect 243997 292632 288572 292634
rect 243997 292576 244002 292632
rect 244058 292576 288572 292632
rect 243997 292574 288572 292576
rect 243997 292571 244063 292574
rect 288566 292572 288572 292574
rect 288636 292572 288642 292636
rect 201401 292498 201467 292501
rect 200806 292496 201467 292498
rect 200806 292440 201406 292496
rect 201462 292440 201467 292496
rect 200806 292438 201467 292440
rect 200806 291924 200866 292438
rect 201401 292435 201467 292438
rect 249149 292362 249215 292365
rect 285673 292362 285739 292365
rect 249149 292360 285739 292362
rect 249149 292304 249154 292360
rect 249210 292304 285678 292360
rect 285734 292304 285739 292360
rect 249149 292302 285739 292304
rect 249149 292299 249215 292302
rect 285673 292299 285739 292302
rect 242341 292226 242407 292229
rect 313273 292226 313339 292229
rect 242341 292224 313339 292226
rect 242341 292168 242346 292224
rect 242402 292168 313278 292224
rect 313334 292168 313339 292224
rect 242341 292166 313339 292168
rect 242341 292163 242407 292166
rect 313273 292163 313339 292166
rect 252553 291954 252619 291957
rect 250148 291952 252619 291954
rect 250148 291896 252558 291952
rect 252614 291896 252619 291952
rect 250148 291894 252619 291896
rect 252553 291891 252619 291894
rect 200113 291548 200179 291549
rect 200062 291484 200068 291548
rect 200132 291546 200179 291548
rect 200132 291544 200224 291546
rect 200174 291488 200224 291544
rect 200132 291486 200224 291488
rect 200132 291484 200179 291486
rect 200113 291483 200179 291484
rect 197353 291274 197419 291277
rect 253749 291274 253815 291277
rect 197353 291272 200284 291274
rect 197353 291216 197358 291272
rect 197414 291216 200284 291272
rect 197353 291214 200284 291216
rect 250148 291272 253815 291274
rect 250148 291216 253754 291272
rect 253810 291216 253815 291272
rect 250148 291214 253815 291216
rect 197353 291211 197419 291214
rect 253749 291211 253815 291214
rect 3417 290866 3483 290869
rect 3417 290864 200130 290866
rect 3417 290808 3422 290864
rect 3478 290808 200130 290864
rect 3417 290806 200130 290808
rect 3417 290803 3483 290806
rect 200070 290732 200130 290806
rect 200062 290668 200068 290732
rect 200132 290668 200138 290732
rect 197353 290594 197419 290597
rect 254117 290594 254183 290597
rect 197353 290592 200284 290594
rect 197353 290536 197358 290592
rect 197414 290536 200284 290592
rect 197353 290534 200284 290536
rect 250148 290592 254183 290594
rect 250148 290536 254122 290592
rect 254178 290536 254183 290592
rect 250148 290534 254183 290536
rect 197353 290531 197419 290534
rect 254117 290531 254183 290534
rect 195830 289852 195836 289916
rect 195900 289914 195906 289916
rect 253749 289914 253815 289917
rect 195900 289854 200284 289914
rect 250148 289912 253815 289914
rect 250148 289856 253754 289912
rect 253810 289856 253815 289912
rect 250148 289854 253815 289856
rect 195900 289852 195906 289854
rect 253749 289851 253815 289854
rect 197353 289234 197419 289237
rect 252921 289234 252987 289237
rect 197353 289232 200284 289234
rect 197353 289176 197358 289232
rect 197414 289176 200284 289232
rect 197353 289174 200284 289176
rect 250148 289232 252987 289234
rect 250148 289176 252926 289232
rect 252982 289176 252987 289232
rect 250148 289174 252987 289176
rect 197353 289171 197419 289174
rect 252921 289171 252987 289174
rect 197721 288554 197787 288557
rect 253749 288554 253815 288557
rect 197721 288552 200284 288554
rect 197721 288496 197726 288552
rect 197782 288496 200284 288552
rect 197721 288494 200284 288496
rect 250148 288552 253815 288554
rect 250148 288496 253754 288552
rect 253810 288496 253815 288552
rect 250148 288494 253815 288496
rect 197721 288491 197787 288494
rect 253749 288491 253815 288494
rect 197445 287874 197511 287877
rect 253749 287874 253815 287877
rect 197445 287872 200284 287874
rect 197445 287816 197450 287872
rect 197506 287816 200284 287872
rect 197445 287814 200284 287816
rect 250148 287872 253815 287874
rect 250148 287816 253754 287872
rect 253810 287816 253815 287872
rect 250148 287814 253815 287816
rect 197445 287811 197511 287814
rect 253749 287811 253815 287814
rect 249977 287602 250043 287605
rect 249934 287600 250043 287602
rect 249934 287544 249982 287600
rect 250038 287544 250043 287600
rect 249934 287539 250043 287544
rect 197353 287194 197419 287197
rect 197353 287192 200284 287194
rect 197353 287136 197358 287192
rect 197414 287136 200284 287192
rect 249934 287164 249994 287539
rect 197353 287134 200284 287136
rect 197353 287131 197419 287134
rect 197353 286514 197419 286517
rect 251265 286514 251331 286517
rect 197353 286512 200284 286514
rect 197353 286456 197358 286512
rect 197414 286456 200284 286512
rect 197353 286454 200284 286456
rect 250148 286512 251331 286514
rect 250148 286456 251270 286512
rect 251326 286456 251331 286512
rect 250148 286454 251331 286456
rect 197353 286451 197419 286454
rect 251265 286451 251331 286454
rect 197997 285834 198063 285837
rect 253749 285834 253815 285837
rect 197997 285832 200284 285834
rect 197997 285776 198002 285832
rect 198058 285776 200284 285832
rect 197997 285774 200284 285776
rect 250148 285832 253815 285834
rect 250148 285776 253754 285832
rect 253810 285776 253815 285832
rect 250148 285774 253815 285776
rect 197997 285771 198063 285774
rect 253749 285771 253815 285774
rect 583520 285276 584960 285516
rect 197353 285154 197419 285157
rect 253054 285154 253060 285156
rect 197353 285152 200284 285154
rect 197353 285096 197358 285152
rect 197414 285096 200284 285152
rect 197353 285094 200284 285096
rect 250148 285094 253060 285154
rect 197353 285091 197419 285094
rect 253054 285092 253060 285094
rect 253124 285092 253130 285156
rect 197261 284474 197327 284477
rect 253841 284474 253907 284477
rect 197261 284472 200284 284474
rect 197261 284416 197266 284472
rect 197322 284416 200284 284472
rect 197261 284414 200284 284416
rect 250148 284472 253907 284474
rect 250148 284416 253846 284472
rect 253902 284416 253907 284472
rect 250148 284414 253907 284416
rect 197261 284411 197327 284414
rect 253841 284411 253907 284414
rect 195646 283732 195652 283796
rect 195716 283794 195722 283796
rect 253289 283794 253355 283797
rect 195716 283734 200284 283794
rect 250148 283792 253355 283794
rect 250148 283736 253294 283792
rect 253350 283736 253355 283792
rect 250148 283734 253355 283736
rect 195716 283732 195722 283734
rect 253289 283731 253355 283734
rect 198549 283114 198615 283117
rect 253749 283114 253815 283117
rect 198549 283112 200284 283114
rect 198549 283056 198554 283112
rect 198610 283056 200284 283112
rect 198549 283054 200284 283056
rect 250148 283112 253815 283114
rect 250148 283056 253754 283112
rect 253810 283056 253815 283112
rect 250148 283054 253815 283056
rect 198549 283051 198615 283054
rect 253749 283051 253815 283054
rect 250118 282026 250178 282404
rect 250437 282026 250503 282029
rect 250118 282024 250503 282026
rect 250118 281968 250442 282024
rect 250498 281968 250503 282024
rect 250118 281966 250503 281968
rect 250437 281963 250503 281966
rect 198641 281754 198707 281757
rect 250294 281754 250300 281756
rect 198641 281752 200284 281754
rect 198641 281696 198646 281752
rect 198702 281696 200284 281752
rect 198641 281694 200284 281696
rect 250148 281694 250300 281754
rect 198641 281691 198707 281694
rect 250294 281692 250300 281694
rect 250364 281692 250370 281756
rect 198641 281074 198707 281077
rect 253749 281074 253815 281077
rect 198641 281072 200284 281074
rect 198641 281016 198646 281072
rect 198702 281016 200284 281072
rect 198641 281014 200284 281016
rect 250148 281072 253815 281074
rect 250148 281016 253754 281072
rect 253810 281016 253815 281072
rect 250148 281014 253815 281016
rect 198641 281011 198707 281014
rect 253749 281011 253815 281014
rect 197353 280394 197419 280397
rect 252553 280394 252619 280397
rect 197353 280392 200284 280394
rect 197353 280336 197358 280392
rect 197414 280336 200284 280392
rect 197353 280334 200284 280336
rect 250148 280392 252619 280394
rect 250148 280336 252558 280392
rect 252614 280336 252619 280392
rect 250148 280334 252619 280336
rect 197353 280331 197419 280334
rect 252553 280331 252619 280334
rect -960 279972 480 280212
rect 197353 279714 197419 279717
rect 197353 279712 200284 279714
rect 197353 279656 197358 279712
rect 197414 279656 200284 279712
rect 197353 279654 200284 279656
rect 197353 279651 197419 279654
rect 250118 279306 250178 279684
rect 250118 279246 258090 279306
rect 200021 279034 200087 279037
rect 252001 279034 252067 279037
rect 200021 279032 200284 279034
rect 200021 278976 200026 279032
rect 200082 278976 200284 279032
rect 200021 278974 200284 278976
rect 250148 279032 252067 279034
rect 250148 278976 252006 279032
rect 252062 278976 252067 279032
rect 250148 278974 252067 278976
rect 258030 279034 258090 279246
rect 278814 279034 278820 279036
rect 258030 278974 278820 279034
rect 200021 278971 200087 278974
rect 252001 278971 252067 278974
rect 278814 278972 278820 278974
rect 278884 278972 278890 279036
rect 197445 278354 197511 278357
rect 253749 278354 253815 278357
rect 197445 278352 200284 278354
rect 197445 278296 197450 278352
rect 197506 278296 200284 278352
rect 197445 278294 200284 278296
rect 250148 278352 253815 278354
rect 250148 278296 253754 278352
rect 253810 278296 253815 278352
rect 250148 278294 253815 278296
rect 197445 278291 197511 278294
rect 253749 278291 253815 278294
rect 197353 277674 197419 277677
rect 253841 277674 253907 277677
rect 197353 277672 200284 277674
rect 197353 277616 197358 277672
rect 197414 277616 200284 277672
rect 197353 277614 200284 277616
rect 250148 277672 253907 277674
rect 250148 277616 253846 277672
rect 253902 277616 253907 277672
rect 250148 277614 253907 277616
rect 197353 277611 197419 277614
rect 253841 277611 253907 277614
rect 197353 276994 197419 276997
rect 253289 276994 253355 276997
rect 197353 276992 200284 276994
rect 197353 276936 197358 276992
rect 197414 276936 200284 276992
rect 197353 276934 200284 276936
rect 250148 276992 253355 276994
rect 250148 276936 253294 276992
rect 253350 276936 253355 276992
rect 250148 276934 253355 276936
rect 197353 276931 197419 276934
rect 253289 276931 253355 276934
rect 197721 276314 197787 276317
rect 253473 276314 253539 276317
rect 197721 276312 200284 276314
rect 197721 276256 197726 276312
rect 197782 276256 200284 276312
rect 197721 276254 200284 276256
rect 250148 276312 253539 276314
rect 250148 276256 253478 276312
rect 253534 276256 253539 276312
rect 250148 276254 253539 276256
rect 197721 276251 197787 276254
rect 253473 276251 253539 276254
rect 197445 275634 197511 275637
rect 253289 275634 253355 275637
rect 197445 275632 200284 275634
rect 197445 275576 197450 275632
rect 197506 275576 200284 275632
rect 197445 275574 200284 275576
rect 250148 275632 253355 275634
rect 250148 275576 253294 275632
rect 253350 275576 253355 275632
rect 250148 275574 253355 275576
rect 197445 275571 197511 275574
rect 253289 275571 253355 275574
rect 197353 274954 197419 274957
rect 251214 274954 251220 274956
rect 197353 274952 200284 274954
rect 197353 274896 197358 274952
rect 197414 274896 200284 274952
rect 197353 274894 200284 274896
rect 250148 274894 251220 274954
rect 197353 274891 197419 274894
rect 251214 274892 251220 274894
rect 251284 274892 251290 274956
rect 197353 274274 197419 274277
rect 252645 274274 252711 274277
rect 197353 274272 200284 274274
rect 197353 274216 197358 274272
rect 197414 274216 200284 274272
rect 197353 274214 200284 274216
rect 250148 274272 252711 274274
rect 250148 274216 252650 274272
rect 252706 274216 252711 274272
rect 250148 274214 252711 274216
rect 197353 274211 197419 274214
rect 252645 274211 252711 274214
rect 179321 273866 179387 273869
rect 199878 273866 199884 273868
rect 179321 273864 199884 273866
rect 179321 273808 179326 273864
rect 179382 273808 199884 273864
rect 179321 273806 199884 273808
rect 179321 273803 179387 273806
rect 199878 273804 199884 273806
rect 199948 273804 199954 273868
rect 198089 273594 198155 273597
rect 251265 273594 251331 273597
rect 198089 273592 200284 273594
rect 198089 273536 198094 273592
rect 198150 273536 200284 273592
rect 198089 273534 200284 273536
rect 250148 273592 251331 273594
rect 250148 273536 251270 273592
rect 251326 273536 251331 273592
rect 250148 273534 251331 273536
rect 198089 273531 198155 273534
rect 251265 273531 251331 273534
rect 196985 272914 197051 272917
rect 253197 272914 253263 272917
rect 196985 272912 200284 272914
rect 196985 272856 196990 272912
rect 197046 272856 200284 272912
rect 196985 272854 200284 272856
rect 250148 272912 253263 272914
rect 250148 272856 253202 272912
rect 253258 272856 253263 272912
rect 250148 272854 253263 272856
rect 196985 272851 197051 272854
rect 253197 272851 253263 272854
rect 197261 272234 197327 272237
rect 252645 272234 252711 272237
rect 197261 272232 200284 272234
rect 197261 272176 197266 272232
rect 197322 272176 200284 272232
rect 197261 272174 200284 272176
rect 250148 272232 252711 272234
rect 250148 272176 252650 272232
rect 252706 272176 252711 272232
rect 250148 272174 252711 272176
rect 197261 272171 197327 272174
rect 252645 272171 252711 272174
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 197445 271554 197511 271557
rect 251357 271554 251423 271557
rect 197445 271552 200284 271554
rect 197445 271496 197450 271552
rect 197506 271496 200284 271552
rect 197445 271494 200284 271496
rect 250148 271552 251423 271554
rect 250148 271496 251362 271552
rect 251418 271496 251423 271552
rect 250148 271494 251423 271496
rect 197445 271491 197511 271494
rect 251357 271491 251423 271494
rect 197353 270874 197419 270877
rect 197353 270872 200284 270874
rect 197353 270816 197358 270872
rect 197414 270816 200284 270872
rect 197353 270814 200284 270816
rect 197353 270811 197419 270814
rect 197445 270194 197511 270197
rect 197445 270192 200284 270194
rect 197445 270136 197450 270192
rect 197506 270136 200284 270192
rect 197445 270134 200284 270136
rect 197445 270131 197511 270134
rect 249934 269789 249994 270164
rect 249934 269784 250043 269789
rect 249934 269728 249982 269784
rect 250038 269728 250043 269784
rect 249934 269726 250043 269728
rect 249977 269723 250043 269726
rect 197353 269514 197419 269517
rect 197353 269512 200284 269514
rect 197353 269456 197358 269512
rect 197414 269456 200284 269512
rect 197353 269454 200284 269456
rect 197353 269451 197419 269454
rect 249750 269244 249810 269484
rect 249742 269180 249748 269244
rect 249812 269180 249818 269244
rect 200021 268834 200087 268837
rect 252645 268834 252711 268837
rect 200021 268832 200284 268834
rect 200021 268776 200026 268832
rect 200082 268776 200284 268832
rect 200021 268774 200284 268776
rect 250148 268832 252711 268834
rect 250148 268776 252650 268832
rect 252706 268776 252711 268832
rect 250148 268774 252711 268776
rect 200021 268771 200087 268774
rect 252645 268771 252711 268774
rect 249558 268364 249564 268428
rect 249628 268426 249634 268428
rect 262397 268426 262463 268429
rect 249628 268424 262463 268426
rect 249628 268368 262402 268424
rect 262458 268368 262463 268424
rect 249628 268366 262463 268368
rect 249628 268364 249634 268366
rect 262397 268363 262463 268366
rect 197353 268154 197419 268157
rect 253197 268154 253263 268157
rect 197353 268152 200284 268154
rect 197353 268096 197358 268152
rect 197414 268096 200284 268152
rect 197353 268094 200284 268096
rect 250148 268152 253263 268154
rect 250148 268096 253202 268152
rect 253258 268096 253263 268152
rect 250148 268094 253263 268096
rect 197353 268091 197419 268094
rect 253197 268091 253263 268094
rect 197445 267474 197511 267477
rect 253289 267474 253355 267477
rect 197445 267472 200284 267474
rect 197445 267416 197450 267472
rect 197506 267416 200284 267472
rect 197445 267414 200284 267416
rect 250148 267472 253355 267474
rect 250148 267416 253294 267472
rect 253350 267416 253355 267472
rect 250148 267414 253355 267416
rect 197445 267411 197511 267414
rect 253289 267411 253355 267414
rect -960 267202 480 267292
rect 3601 267202 3667 267205
rect -960 267200 3667 267202
rect -960 267144 3606 267200
rect 3662 267144 3667 267200
rect -960 267142 3667 267144
rect -960 267052 480 267142
rect 3601 267139 3667 267142
rect 197353 266794 197419 266797
rect 253749 266794 253815 266797
rect 197353 266792 200284 266794
rect 197353 266736 197358 266792
rect 197414 266736 200284 266792
rect 197353 266734 200284 266736
rect 250148 266792 253815 266794
rect 250148 266736 253754 266792
rect 253810 266736 253815 266792
rect 250148 266734 253815 266736
rect 197353 266731 197419 266734
rect 253749 266731 253815 266734
rect 197445 266114 197511 266117
rect 253841 266114 253907 266117
rect 197445 266112 200284 266114
rect 197445 266056 197450 266112
rect 197506 266056 200284 266112
rect 197445 266054 200284 266056
rect 250148 266112 253907 266114
rect 250148 266056 253846 266112
rect 253902 266056 253907 266112
rect 250148 266054 253907 266056
rect 197445 266051 197511 266054
rect 253841 266051 253907 266054
rect 197353 265434 197419 265437
rect 253749 265434 253815 265437
rect 197353 265432 200284 265434
rect 197353 265376 197358 265432
rect 197414 265376 200284 265432
rect 197353 265374 200284 265376
rect 250148 265432 253815 265434
rect 250148 265376 253754 265432
rect 253810 265376 253815 265432
rect 250148 265374 253815 265376
rect 197353 265371 197419 265374
rect 253749 265371 253815 265374
rect 197445 264754 197511 264757
rect 253749 264754 253815 264757
rect 197445 264752 200284 264754
rect 197445 264696 197450 264752
rect 197506 264696 200284 264752
rect 197445 264694 200284 264696
rect 250148 264752 253815 264754
rect 250148 264696 253754 264752
rect 253810 264696 253815 264752
rect 250148 264694 253815 264696
rect 197445 264691 197511 264694
rect 253749 264691 253815 264694
rect 197353 264074 197419 264077
rect 252737 264074 252803 264077
rect 197353 264072 200284 264074
rect 197353 264016 197358 264072
rect 197414 264016 200284 264072
rect 197353 264014 200284 264016
rect 250148 264072 252803 264074
rect 250148 264016 252742 264072
rect 252798 264016 252803 264072
rect 250148 264014 252803 264016
rect 197353 264011 197419 264014
rect 252737 264011 252803 264014
rect 197353 263394 197419 263397
rect 252553 263394 252619 263397
rect 197353 263392 200284 263394
rect 197353 263336 197358 263392
rect 197414 263336 200284 263392
rect 197353 263334 200284 263336
rect 250148 263392 252619 263394
rect 250148 263336 252558 263392
rect 252614 263336 252619 263392
rect 250148 263334 252619 263336
rect 197353 263331 197419 263334
rect 252553 263331 252619 263334
rect 197353 262714 197419 262717
rect 253749 262714 253815 262717
rect 197353 262712 200284 262714
rect 197353 262656 197358 262712
rect 197414 262656 200284 262712
rect 197353 262654 200284 262656
rect 250148 262712 253815 262714
rect 250148 262656 253754 262712
rect 253810 262656 253815 262712
rect 250148 262654 253815 262656
rect 197353 262651 197419 262654
rect 253749 262651 253815 262654
rect 197445 262034 197511 262037
rect 253381 262034 253447 262037
rect 197445 262032 200284 262034
rect 197445 261976 197450 262032
rect 197506 261976 200284 262032
rect 197445 261974 200284 261976
rect 250148 262032 253447 262034
rect 250148 261976 253386 262032
rect 253442 261976 253447 262032
rect 250148 261974 253447 261976
rect 197445 261971 197511 261974
rect 253381 261971 253447 261974
rect 197537 261354 197603 261357
rect 251173 261354 251239 261357
rect 197537 261352 200284 261354
rect 197537 261296 197542 261352
rect 197598 261296 200284 261352
rect 197537 261294 200284 261296
rect 250148 261352 251239 261354
rect 250148 261296 251178 261352
rect 251234 261296 251239 261352
rect 250148 261294 251239 261296
rect 197537 261291 197603 261294
rect 251173 261291 251239 261294
rect 197353 260674 197419 260677
rect 252829 260674 252895 260677
rect 197353 260672 200284 260674
rect 197353 260616 197358 260672
rect 197414 260616 200284 260672
rect 197353 260614 200284 260616
rect 250148 260672 252895 260674
rect 250148 260616 252834 260672
rect 252890 260616 252895 260672
rect 250148 260614 252895 260616
rect 197353 260611 197419 260614
rect 252829 260611 252895 260614
rect 197353 259994 197419 259997
rect 253197 259994 253263 259997
rect 197353 259992 200284 259994
rect 197353 259936 197358 259992
rect 197414 259936 200284 259992
rect 197353 259934 200284 259936
rect 250148 259992 253263 259994
rect 250148 259936 253202 259992
rect 253258 259936 253263 259992
rect 250148 259934 253263 259936
rect 197353 259931 197419 259934
rect 253197 259931 253263 259934
rect 197353 259314 197419 259317
rect 197353 259312 200284 259314
rect 197353 259256 197358 259312
rect 197414 259256 200284 259312
rect 197353 259254 200284 259256
rect 197353 259251 197419 259254
rect 250118 258906 250178 259284
rect 250345 258906 250411 258909
rect 250118 258904 250411 258906
rect 250118 258848 250350 258904
rect 250406 258848 250411 258904
rect 250118 258846 250411 258848
rect 250345 258843 250411 258846
rect 579613 258906 579679 258909
rect 583520 258906 584960 258996
rect 579613 258904 584960 258906
rect 579613 258848 579618 258904
rect 579674 258848 584960 258904
rect 579613 258846 584960 258848
rect 579613 258843 579679 258846
rect 583520 258756 584960 258846
rect 197445 258634 197511 258637
rect 252553 258634 252619 258637
rect 197445 258632 200284 258634
rect 197445 258576 197450 258632
rect 197506 258576 200284 258632
rect 197445 258574 200284 258576
rect 250148 258632 252619 258634
rect 250148 258576 252558 258632
rect 252614 258576 252619 258632
rect 250148 258574 252619 258576
rect 197445 258571 197511 258574
rect 252553 258571 252619 258574
rect 197445 257954 197511 257957
rect 251173 257954 251239 257957
rect 197445 257952 200284 257954
rect 197445 257896 197450 257952
rect 197506 257896 200284 257952
rect 197445 257894 200284 257896
rect 250148 257952 251239 257954
rect 250148 257896 251178 257952
rect 251234 257896 251239 257952
rect 250148 257894 251239 257896
rect 197445 257891 197511 257894
rect 251173 257891 251239 257894
rect 197353 257274 197419 257277
rect 253013 257274 253079 257277
rect 197353 257272 200284 257274
rect 197353 257216 197358 257272
rect 197414 257216 200284 257272
rect 197353 257214 200284 257216
rect 250148 257272 253079 257274
rect 250148 257216 253018 257272
rect 253074 257216 253079 257272
rect 250148 257214 253079 257216
rect 197353 257211 197419 257214
rect 253013 257211 253079 257214
rect 199929 256594 199995 256597
rect 253749 256594 253815 256597
rect 199929 256592 200284 256594
rect 199929 256536 199934 256592
rect 199990 256536 200284 256592
rect 199929 256534 200284 256536
rect 250148 256592 253815 256594
rect 250148 256536 253754 256592
rect 253810 256536 253815 256592
rect 250148 256534 253815 256536
rect 199929 256531 199995 256534
rect 253749 256531 253815 256534
rect 197445 255914 197511 255917
rect 253105 255914 253171 255917
rect 197445 255912 200284 255914
rect 197445 255856 197450 255912
rect 197506 255856 200284 255912
rect 197445 255854 200284 255856
rect 250148 255912 253171 255914
rect 250148 255856 253110 255912
rect 253166 255856 253171 255912
rect 250148 255854 253171 255856
rect 197445 255851 197511 255854
rect 253105 255851 253171 255854
rect 197353 255234 197419 255237
rect 253749 255234 253815 255237
rect 197353 255232 200284 255234
rect 197353 255176 197358 255232
rect 197414 255176 200284 255232
rect 197353 255174 200284 255176
rect 250148 255232 253815 255234
rect 250148 255176 253754 255232
rect 253810 255176 253815 255232
rect 250148 255174 253815 255176
rect 197353 255171 197419 255174
rect 253749 255171 253815 255174
rect 197353 254554 197419 254557
rect 253013 254554 253079 254557
rect 197353 254552 200284 254554
rect 197353 254496 197358 254552
rect 197414 254496 200284 254552
rect 197353 254494 200284 254496
rect 250148 254552 253079 254554
rect 250148 254496 253018 254552
rect 253074 254496 253079 254552
rect 250148 254494 253079 254496
rect 197353 254491 197419 254494
rect 253013 254491 253079 254494
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 197353 253874 197419 253877
rect 197353 253872 200284 253874
rect 197353 253816 197358 253872
rect 197414 253816 200284 253872
rect 197353 253814 200284 253816
rect 197353 253811 197419 253814
rect 250118 253469 250178 253844
rect 250069 253464 250178 253469
rect 250069 253408 250074 253464
rect 250130 253408 250178 253464
rect 250069 253406 250178 253408
rect 250069 253403 250135 253406
rect 199837 253194 199903 253197
rect 253841 253194 253907 253197
rect 199837 253192 200284 253194
rect 199837 253136 199842 253192
rect 199898 253136 200284 253192
rect 199837 253134 200284 253136
rect 250148 253192 253907 253194
rect 250148 253136 253846 253192
rect 253902 253136 253907 253192
rect 250148 253134 253907 253136
rect 199837 253131 199903 253134
rect 253841 253131 253907 253134
rect 197445 252514 197511 252517
rect 253749 252514 253815 252517
rect 197445 252512 200284 252514
rect 197445 252456 197450 252512
rect 197506 252456 200284 252512
rect 197445 252454 200284 252456
rect 250148 252512 253815 252514
rect 250148 252456 253754 252512
rect 253810 252456 253815 252512
rect 250148 252454 253815 252456
rect 197445 252451 197511 252454
rect 253749 252451 253815 252454
rect 197118 252316 197124 252380
rect 197188 252378 197194 252380
rect 197997 252378 198063 252381
rect 197188 252376 198063 252378
rect 197188 252320 198002 252376
rect 198058 252320 198063 252376
rect 197188 252318 198063 252320
rect 197188 252316 197194 252318
rect 197997 252315 198063 252318
rect 197353 251834 197419 251837
rect 253473 251834 253539 251837
rect 197353 251832 200284 251834
rect 197353 251776 197358 251832
rect 197414 251776 200284 251832
rect 197353 251774 200284 251776
rect 250148 251832 253539 251834
rect 250148 251776 253478 251832
rect 253534 251776 253539 251832
rect 250148 251774 253539 251776
rect 197353 251771 197419 251774
rect 253473 251771 253539 251774
rect 198549 251154 198615 251157
rect 253381 251154 253447 251157
rect 198549 251152 200284 251154
rect 198549 251096 198554 251152
rect 198610 251096 200284 251152
rect 198549 251094 200284 251096
rect 250148 251152 253447 251154
rect 250148 251096 253386 251152
rect 253442 251096 253447 251152
rect 250148 251094 253447 251096
rect 198549 251091 198615 251094
rect 253381 251091 253447 251094
rect 197445 250474 197511 250477
rect 252737 250474 252803 250477
rect 197445 250472 200284 250474
rect 197445 250416 197450 250472
rect 197506 250416 200284 250472
rect 197445 250414 200284 250416
rect 250148 250472 252803 250474
rect 250148 250416 252742 250472
rect 252798 250416 252803 250472
rect 250148 250414 252803 250416
rect 197445 250411 197511 250414
rect 252737 250411 252803 250414
rect 197353 249794 197419 249797
rect 253749 249794 253815 249797
rect 197353 249792 200284 249794
rect 197353 249736 197358 249792
rect 197414 249736 200284 249792
rect 197353 249734 200284 249736
rect 250148 249792 253815 249794
rect 250148 249736 253754 249792
rect 253810 249736 253815 249792
rect 250148 249734 253815 249736
rect 197353 249731 197419 249734
rect 253749 249731 253815 249734
rect 197353 249114 197419 249117
rect 253749 249114 253815 249117
rect 197353 249112 200284 249114
rect 197353 249056 197358 249112
rect 197414 249056 200284 249112
rect 197353 249054 200284 249056
rect 250148 249112 253815 249114
rect 250148 249056 253754 249112
rect 253810 249056 253815 249112
rect 250148 249054 253815 249056
rect 197353 249051 197419 249054
rect 253749 249051 253815 249054
rect 197169 248434 197235 248437
rect 252645 248434 252711 248437
rect 197169 248432 200284 248434
rect 197169 248376 197174 248432
rect 197230 248376 200284 248432
rect 197169 248374 200284 248376
rect 250148 248432 252711 248434
rect 250148 248376 252650 248432
rect 252706 248376 252711 248432
rect 250148 248374 252711 248376
rect 197169 248371 197235 248374
rect 252645 248371 252711 248374
rect 197537 247754 197603 247757
rect 253841 247754 253907 247757
rect 197537 247752 200284 247754
rect 197537 247696 197542 247752
rect 197598 247696 200284 247752
rect 197537 247694 200284 247696
rect 250148 247752 253907 247754
rect 250148 247696 253846 247752
rect 253902 247696 253907 247752
rect 250148 247694 253907 247696
rect 197537 247691 197603 247694
rect 253841 247691 253907 247694
rect 197445 247074 197511 247077
rect 253749 247074 253815 247077
rect 197445 247072 200284 247074
rect 197445 247016 197450 247072
rect 197506 247016 200284 247072
rect 197445 247014 200284 247016
rect 250148 247072 253815 247074
rect 250148 247016 253754 247072
rect 253810 247016 253815 247072
rect 250148 247014 253815 247016
rect 197445 247011 197511 247014
rect 253749 247011 253815 247014
rect 252502 246394 252508 246396
rect 200622 245988 200682 246364
rect 250148 246334 252508 246394
rect 252502 246332 252508 246334
rect 252572 246332 252578 246396
rect 200614 245924 200620 245988
rect 200684 245924 200690 245988
rect 197353 245714 197419 245717
rect 253749 245714 253815 245717
rect 197353 245712 200284 245714
rect 197353 245656 197358 245712
rect 197414 245656 200284 245712
rect 197353 245654 200284 245656
rect 250148 245712 253815 245714
rect 250148 245656 253754 245712
rect 253810 245656 253815 245712
rect 250148 245654 253815 245656
rect 197353 245651 197419 245654
rect 253749 245651 253815 245654
rect 579889 245578 579955 245581
rect 583520 245578 584960 245668
rect 579889 245576 584960 245578
rect 579889 245520 579894 245576
rect 579950 245520 584960 245576
rect 579889 245518 584960 245520
rect 579889 245515 579955 245518
rect 583520 245428 584960 245518
rect 199745 245034 199811 245037
rect 253841 245034 253907 245037
rect 199745 245032 200284 245034
rect 199745 244976 199750 245032
rect 199806 244976 200284 245032
rect 199745 244974 200284 244976
rect 250148 245032 253907 245034
rect 250148 244976 253846 245032
rect 253902 244976 253907 245032
rect 250148 244974 253907 244976
rect 199745 244971 199811 244974
rect 253841 244971 253907 244974
rect 197445 244354 197511 244357
rect 253749 244354 253815 244357
rect 197445 244352 200284 244354
rect 197445 244296 197450 244352
rect 197506 244296 200284 244352
rect 197445 244294 200284 244296
rect 250148 244352 253815 244354
rect 250148 244296 253754 244352
rect 253810 244296 253815 244352
rect 250148 244294 253815 244296
rect 197445 244291 197511 244294
rect 253749 244291 253815 244294
rect 197353 243674 197419 243677
rect 253749 243674 253815 243677
rect 197353 243672 200284 243674
rect 197353 243616 197358 243672
rect 197414 243616 200284 243672
rect 197353 243614 200284 243616
rect 250148 243672 253815 243674
rect 250148 243616 253754 243672
rect 253810 243616 253815 243672
rect 250148 243614 253815 243616
rect 197353 243611 197419 243614
rect 253749 243611 253815 243614
rect 191598 242932 191604 242996
rect 191668 242994 191674 242996
rect 253381 242994 253447 242997
rect 191668 242934 200284 242994
rect 250148 242992 253447 242994
rect 250148 242936 253386 242992
rect 253442 242936 253447 242992
rect 250148 242934 253447 242936
rect 191668 242932 191674 242934
rect 253381 242931 253447 242934
rect 197353 242314 197419 242317
rect 253749 242314 253815 242317
rect 197353 242312 200284 242314
rect 197353 242256 197358 242312
rect 197414 242256 200284 242312
rect 197353 242254 200284 242256
rect 250148 242312 253815 242314
rect 250148 242256 253754 242312
rect 253810 242256 253815 242312
rect 250148 242254 253815 242256
rect 197353 242251 197419 242254
rect 253749 242251 253815 242254
rect 104893 242178 104959 242181
rect 192334 242178 192340 242180
rect 104893 242176 192340 242178
rect 104893 242120 104898 242176
rect 104954 242120 192340 242176
rect 104893 242118 192340 242120
rect 104893 242115 104959 242118
rect 192334 242116 192340 242118
rect 192404 242116 192410 242180
rect 187550 241572 187556 241636
rect 187620 241634 187626 241636
rect 252553 241634 252619 241637
rect 187620 241574 200284 241634
rect 250148 241632 252619 241634
rect 250148 241576 252558 241632
rect 252614 241576 252619 241632
rect 250148 241574 252619 241576
rect 187620 241572 187626 241574
rect 252553 241571 252619 241574
rect -960 241090 480 241180
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 200806 240141 200866 240924
rect 250118 240546 250178 240924
rect 251081 240546 251147 240549
rect 250118 240544 251147 240546
rect 250118 240488 251086 240544
rect 251142 240488 251147 240544
rect 250118 240486 251147 240488
rect 251081 240483 251147 240486
rect 250253 240410 250319 240413
rect 256877 240410 256943 240413
rect 250253 240408 256943 240410
rect 250253 240352 250258 240408
rect 250314 240352 256882 240408
rect 256938 240352 256943 240408
rect 250253 240350 256943 240352
rect 250253 240347 250319 240350
rect 256877 240347 256943 240350
rect 253749 240274 253815 240277
rect 250148 240272 253815 240274
rect 250148 240216 253754 240272
rect 253810 240216 253815 240272
rect 250148 240214 253815 240216
rect 253749 240211 253815 240214
rect 190545 240140 190611 240141
rect 190494 240138 190500 240140
rect 190454 240078 190500 240138
rect 190564 240136 190611 240140
rect 190606 240080 190611 240136
rect 190494 240076 190500 240078
rect 190564 240076 190611 240080
rect 190545 240075 190611 240076
rect 200757 240136 200866 240141
rect 200757 240080 200762 240136
rect 200818 240080 200866 240136
rect 200757 240078 200866 240080
rect 200757 240075 200823 240078
rect 248513 240002 248579 240005
rect 262857 240002 262923 240005
rect 248513 240000 262923 240002
rect 248513 239944 248518 240000
rect 248574 239944 262862 240000
rect 262918 239944 262923 240000
rect 248513 239942 262923 239944
rect 248513 239939 248579 239942
rect 262857 239939 262923 239942
rect 197077 239730 197143 239733
rect 236494 239730 236500 239732
rect 197077 239728 236500 239730
rect 197077 239672 197082 239728
rect 197138 239672 236500 239728
rect 197077 239670 236500 239672
rect 197077 239667 197143 239670
rect 236494 239668 236500 239670
rect 236564 239668 236570 239732
rect 238518 239668 238524 239732
rect 238588 239730 238594 239732
rect 238753 239730 238819 239733
rect 238588 239728 238819 239730
rect 238588 239672 238758 239728
rect 238814 239672 238819 239728
rect 238588 239670 238819 239672
rect 238588 239668 238594 239670
rect 238753 239667 238819 239670
rect 192937 239594 193003 239597
rect 237414 239594 237420 239596
rect 192937 239592 237420 239594
rect 192937 239536 192942 239592
rect 192998 239536 237420 239592
rect 192937 239534 237420 239536
rect 192937 239531 193003 239534
rect 237414 239532 237420 239534
rect 237484 239532 237490 239596
rect 199745 239458 199811 239461
rect 241646 239458 241652 239460
rect 199745 239456 241652 239458
rect 199745 239400 199750 239456
rect 199806 239400 241652 239456
rect 199745 239398 241652 239400
rect 199745 239395 199811 239398
rect 241646 239396 241652 239398
rect 241716 239396 241722 239460
rect 40033 238642 40099 238645
rect 225965 238642 226031 238645
rect 40033 238640 226031 238642
rect 40033 238584 40038 238640
rect 40094 238584 225970 238640
rect 226026 238584 226031 238640
rect 40033 238582 226031 238584
rect 40033 238579 40099 238582
rect 225965 238579 226031 238582
rect 249149 238642 249215 238645
rect 255814 238642 255820 238644
rect 249149 238640 255820 238642
rect 249149 238584 249154 238640
rect 249210 238584 255820 238640
rect 249149 238582 255820 238584
rect 249149 238579 249215 238582
rect 255814 238580 255820 238582
rect 255884 238580 255890 238644
rect 192334 238444 192340 238508
rect 192404 238506 192410 238508
rect 219525 238506 219591 238509
rect 192404 238504 219591 238506
rect 192404 238448 219530 238504
rect 219586 238448 219591 238504
rect 192404 238446 219591 238448
rect 192404 238444 192410 238446
rect 219525 238443 219591 238446
rect 200614 236540 200620 236604
rect 200684 236602 200690 236604
rect 281533 236602 281599 236605
rect 200684 236600 281599 236602
rect 200684 236544 281538 236600
rect 281594 236544 281599 236600
rect 200684 236542 281599 236544
rect 200684 236540 200690 236542
rect 281533 236539 281599 236542
rect 244774 235180 244780 235244
rect 244844 235242 244850 235244
rect 258165 235242 258231 235245
rect 244844 235240 258231 235242
rect 244844 235184 258170 235240
rect 258226 235184 258231 235240
rect 244844 235182 258231 235184
rect 244844 235180 244850 235182
rect 258165 235179 258231 235182
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 213085 228306 213151 228309
rect 298686 228306 298692 228308
rect 213085 228304 298692 228306
rect 213085 228248 213090 228304
rect 213146 228248 298692 228304
rect 213085 228246 298692 228248
rect 213085 228243 213151 228246
rect 298686 228244 298692 228246
rect 298756 228244 298762 228308
rect -960 227884 480 228124
rect 583017 219058 583083 219061
rect 583520 219058 584960 219148
rect 583017 219056 584960 219058
rect 583017 219000 583022 219056
rect 583078 219000 584960 219056
rect 583017 218998 584960 219000
rect 583017 218995 583083 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579889 205730 579955 205733
rect 583520 205730 584960 205820
rect 579889 205728 584960 205730
rect 579889 205672 579894 205728
rect 579950 205672 584960 205728
rect 579889 205670 584960 205672
rect 579889 205667 579955 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 207289 197978 207355 197981
rect 287094 197978 287100 197980
rect 207289 197976 287100 197978
rect 207289 197920 207294 197976
rect 207350 197920 287100 197976
rect 207289 197918 287100 197920
rect 207289 197915 207355 197918
rect 287094 197916 287100 197918
rect 287164 197916 287170 197980
rect 198641 193898 198707 193901
rect 285622 193898 285628 193900
rect 198641 193896 285628 193898
rect 198641 193840 198646 193896
rect 198702 193840 285628 193896
rect 198641 193838 285628 193840
rect 198641 193835 198707 193838
rect 285622 193836 285628 193838
rect 285692 193836 285698 193900
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 280797 191178 280863 191181
rect 290590 191178 290596 191180
rect 280797 191176 290596 191178
rect 280797 191120 280802 191176
rect 280858 191120 290596 191176
rect 280797 191118 290596 191120
rect 280797 191115 280863 191118
rect 290590 191116 290596 191118
rect 290660 191116 290666 191180
rect 204713 191042 204779 191045
rect 294270 191042 294276 191044
rect 204713 191040 294276 191042
rect 204713 190984 204718 191040
rect 204774 190984 294276 191040
rect 204713 190982 294276 190984
rect 204713 190979 204779 190982
rect 294270 190980 294276 190982
rect 294340 190980 294346 191044
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 205357 186962 205423 186965
rect 233366 186962 233372 186964
rect 205357 186960 233372 186962
rect 205357 186904 205362 186960
rect 205418 186904 233372 186960
rect 205357 186902 233372 186904
rect 205357 186899 205423 186902
rect 233366 186900 233372 186902
rect 233436 186900 233442 186964
rect 195881 185602 195947 185605
rect 276606 185602 276612 185604
rect 195881 185600 276612 185602
rect 195881 185544 195886 185600
rect 195942 185544 276612 185600
rect 195881 185542 276612 185544
rect 195881 185539 195947 185542
rect 276606 185540 276612 185542
rect 276676 185540 276682 185604
rect 207933 184242 207999 184245
rect 287278 184242 287284 184244
rect 207933 184240 287284 184242
rect 207933 184184 207938 184240
rect 207994 184184 287284 184240
rect 207933 184182 287284 184184
rect 207933 184179 207999 184182
rect 287278 184180 287284 184182
rect 287348 184180 287354 184244
rect 193029 182882 193095 182885
rect 582373 182882 582439 182885
rect 193029 182880 582439 182882
rect 193029 182824 193034 182880
rect 193090 182824 582378 182880
rect 582434 182824 582439 182880
rect 193029 182822 582439 182824
rect 193029 182819 193095 182822
rect 582373 182819 582439 182822
rect 179321 181522 179387 181525
rect 228766 181522 228772 181524
rect 179321 181520 228772 181522
rect 179321 181464 179326 181520
rect 179382 181464 228772 181520
rect 179321 181462 228772 181464
rect 179321 181459 179387 181462
rect 228766 181460 228772 181462
rect 228836 181460 228842 181524
rect 234981 181522 235047 181525
rect 284334 181522 284340 181524
rect 234981 181520 284340 181522
rect 234981 181464 234986 181520
rect 235042 181464 284340 181520
rect 234981 181462 284340 181464
rect 234981 181459 235047 181462
rect 284334 181460 284340 181462
rect 284404 181460 284410 181524
rect 206369 181386 206435 181389
rect 292614 181386 292620 181388
rect 206369 181384 292620 181386
rect 206369 181328 206374 181384
rect 206430 181328 292620 181384
rect 206369 181326 292620 181328
rect 206369 181323 206435 181326
rect 292614 181324 292620 181326
rect 292684 181324 292690 181388
rect 209221 180162 209287 180165
rect 241646 180162 241652 180164
rect 209221 180160 241652 180162
rect 209221 180104 209226 180160
rect 209282 180104 241652 180160
rect 209221 180102 241652 180104
rect 209221 180099 209287 180102
rect 241646 180100 241652 180102
rect 241716 180100 241722 180164
rect 209865 180026 209931 180029
rect 298369 180026 298435 180029
rect 209865 180024 298435 180026
rect 209865 179968 209870 180024
rect 209926 179968 298374 180024
rect 298430 179968 298435 180024
rect 209865 179966 298435 179968
rect 209865 179963 209931 179966
rect 298369 179963 298435 179966
rect 99097 179482 99163 179485
rect 166206 179482 166212 179484
rect 99097 179480 166212 179482
rect 99097 179424 99102 179480
rect 99158 179424 166212 179480
rect 99097 179422 166212 179424
rect 99097 179419 99163 179422
rect 166206 179420 166212 179422
rect 166276 179420 166282 179484
rect 580349 179210 580415 179213
rect 583520 179210 584960 179300
rect 580349 179208 584960 179210
rect 580349 179152 580354 179208
rect 580410 179152 584960 179208
rect 580349 179150 584960 179152
rect 580349 179147 580415 179150
rect 583520 179060 584960 179150
rect 182081 178802 182147 178805
rect 234654 178802 234660 178804
rect 182081 178800 234660 178802
rect 182081 178744 182086 178800
rect 182142 178744 234660 178800
rect 182081 178742 234660 178744
rect 182081 178739 182147 178742
rect 234654 178740 234660 178742
rect 234724 178740 234730 178804
rect 186129 178666 186195 178669
rect 294229 178666 294295 178669
rect 186129 178664 294295 178666
rect 186129 178608 186134 178664
rect 186190 178608 294234 178664
rect 294290 178608 294295 178664
rect 186129 178606 294295 178608
rect 186129 178603 186195 178606
rect 294229 178603 294295 178606
rect 105670 177652 105676 177716
rect 105740 177714 105746 177716
rect 105905 177714 105971 177717
rect 108113 177716 108179 177717
rect 108062 177714 108068 177716
rect 105740 177712 105971 177714
rect 105740 177656 105910 177712
rect 105966 177656 105971 177712
rect 105740 177654 105971 177656
rect 108022 177654 108068 177714
rect 108132 177712 108179 177716
rect 108174 177656 108179 177712
rect 105740 177652 105746 177654
rect 105905 177651 105971 177654
rect 108062 177652 108068 177654
rect 108132 177652 108179 177656
rect 114318 177652 114324 177716
rect 114388 177714 114394 177716
rect 114461 177714 114527 177717
rect 119521 177716 119587 177717
rect 119470 177714 119476 177716
rect 114388 177712 114527 177714
rect 114388 177656 114466 177712
rect 114522 177656 114527 177712
rect 114388 177654 114527 177656
rect 119430 177654 119476 177714
rect 119540 177712 119587 177716
rect 119582 177656 119587 177712
rect 114388 177652 114394 177654
rect 108113 177651 108179 177652
rect 114461 177651 114527 177654
rect 119470 177652 119476 177654
rect 119540 177652 119587 177656
rect 124438 177652 124444 177716
rect 124508 177714 124514 177716
rect 124949 177714 125015 177717
rect 127065 177716 127131 177717
rect 130745 177716 130811 177717
rect 132401 177716 132467 177717
rect 127014 177714 127020 177716
rect 124508 177712 125015 177714
rect 124508 177656 124954 177712
rect 125010 177656 125015 177712
rect 124508 177654 125015 177656
rect 126974 177654 127020 177714
rect 127084 177712 127131 177716
rect 130694 177714 130700 177716
rect 127126 177656 127131 177712
rect 124508 177652 124514 177654
rect 119521 177651 119587 177652
rect 124949 177651 125015 177654
rect 127014 177652 127020 177654
rect 127084 177652 127131 177656
rect 130654 177654 130700 177714
rect 130764 177712 130811 177716
rect 132350 177714 132356 177716
rect 130806 177656 130811 177712
rect 130694 177652 130700 177654
rect 130764 177652 130811 177656
rect 132310 177654 132356 177714
rect 132420 177712 132467 177716
rect 132462 177656 132467 177712
rect 132350 177652 132356 177654
rect 132420 177652 132467 177656
rect 127065 177651 127131 177652
rect 130745 177651 130811 177652
rect 132401 177651 132467 177652
rect 276606 177516 276612 177580
rect 276676 177578 276682 177580
rect 279417 177578 279483 177581
rect 276676 177576 279483 177578
rect 276676 177520 279422 177576
rect 279478 177520 279483 177576
rect 276676 177518 279483 177520
rect 276676 177516 276682 177518
rect 279417 177515 279483 177518
rect 197169 177442 197235 177445
rect 233182 177442 233188 177444
rect 197169 177440 233188 177442
rect 197169 177384 197174 177440
rect 197230 177384 233188 177440
rect 197169 177382 233188 177384
rect 197169 177379 197235 177382
rect 233182 177380 233188 177382
rect 233252 177380 233258 177444
rect 269849 177442 269915 177445
rect 291326 177442 291332 177444
rect 269849 177440 291332 177442
rect 269849 177384 269854 177440
rect 269910 177384 291332 177440
rect 269849 177382 291332 177384
rect 269849 177379 269915 177382
rect 291326 177380 291332 177382
rect 291396 177380 291402 177444
rect 190361 177306 190427 177309
rect 237598 177306 237604 177308
rect 190361 177304 237604 177306
rect 190361 177248 190366 177304
rect 190422 177248 237604 177304
rect 190361 177246 237604 177248
rect 190361 177243 190427 177246
rect 237598 177244 237604 177246
rect 237668 177244 237674 177308
rect 253054 177244 253060 177308
rect 253124 177306 253130 177308
rect 283189 177306 283255 177309
rect 253124 177304 283255 177306
rect 253124 177248 283194 177304
rect 283250 177248 283255 177304
rect 253124 177246 283255 177248
rect 253124 177244 253130 177246
rect 283189 177243 283255 177246
rect 113214 177108 113220 177172
rect 113284 177170 113290 177172
rect 114369 177170 114435 177173
rect 113284 177168 114435 177170
rect 113284 177112 114374 177168
rect 114430 177112 114435 177168
rect 113284 177110 114435 177112
rect 113284 177108 113290 177110
rect 114369 177107 114435 177110
rect 123150 177108 123156 177172
rect 123220 177170 123226 177172
rect 123753 177170 123819 177173
rect 129457 177172 129523 177173
rect 129406 177170 129412 177172
rect 123220 177168 123819 177170
rect 123220 177112 123758 177168
rect 123814 177112 123819 177168
rect 123220 177110 123819 177112
rect 129366 177110 129412 177170
rect 129476 177168 129523 177172
rect 129518 177112 129523 177168
rect 123220 177108 123226 177110
rect 123753 177107 123819 177110
rect 129406 177108 129412 177110
rect 129476 177108 129523 177112
rect 129457 177107 129523 177108
rect 97022 176972 97028 177036
rect 97092 177034 97098 177036
rect 97533 177034 97599 177037
rect 97092 177032 97599 177034
rect 97092 176976 97538 177032
rect 97594 176976 97599 177032
rect 97092 176974 97599 176976
rect 97092 176972 97098 176974
rect 97533 176971 97599 176974
rect 98310 176972 98316 177036
rect 98380 177034 98386 177036
rect 99097 177034 99163 177037
rect 98380 177032 99163 177034
rect 98380 176976 99102 177032
rect 99158 176976 99163 177032
rect 98380 176974 99163 176976
rect 98380 176972 98386 176974
rect 99097 176971 99163 176974
rect 101990 176972 101996 177036
rect 102060 177034 102066 177036
rect 167729 177034 167795 177037
rect 102060 177032 167795 177034
rect 102060 176976 167734 177032
rect 167790 176976 167795 177032
rect 102060 176974 167795 176976
rect 102060 176972 102066 176974
rect 167729 176971 167795 176974
rect 100702 176836 100708 176900
rect 100772 176898 100778 176900
rect 166390 176898 166396 176900
rect 100772 176838 166396 176898
rect 100772 176836 100778 176838
rect 166390 176836 166396 176838
rect 166460 176836 166466 176900
rect 100661 176762 100727 176765
rect 103329 176762 103395 176765
rect 104617 176764 104683 176765
rect 107009 176764 107075 176765
rect 109585 176764 109651 176765
rect 110689 176764 110755 176765
rect 104566 176762 104572 176764
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 103286 176760 103395 176762
rect 103286 176704 103334 176760
rect 103390 176704 103395 176760
rect 103286 176699 103395 176704
rect 104526 176702 104572 176762
rect 104636 176760 104683 176764
rect 106958 176762 106964 176764
rect 104678 176704 104683 176760
rect 104566 176700 104572 176702
rect 104636 176700 104683 176704
rect 106918 176702 106964 176762
rect 107028 176760 107075 176764
rect 109534 176762 109540 176764
rect 107070 176704 107075 176760
rect 106958 176700 106964 176702
rect 107028 176700 107075 176704
rect 109494 176702 109540 176762
rect 109604 176760 109651 176764
rect 110638 176762 110644 176764
rect 109646 176704 109651 176760
rect 109534 176700 109540 176702
rect 109604 176700 109651 176704
rect 110598 176702 110644 176762
rect 110708 176760 110755 176764
rect 110750 176704 110755 176760
rect 110638 176700 110644 176702
rect 110708 176700 110755 176704
rect 112110 176700 112116 176764
rect 112180 176762 112186 176764
rect 112253 176762 112319 176765
rect 118417 176764 118483 176765
rect 118366 176762 118372 176764
rect 112180 176760 112319 176762
rect 112180 176704 112258 176760
rect 112314 176704 112319 176760
rect 112180 176702 112319 176704
rect 118326 176702 118372 176762
rect 118436 176760 118483 176764
rect 118478 176704 118483 176760
rect 112180 176700 112186 176702
rect 104617 176699 104683 176700
rect 107009 176699 107075 176700
rect 109585 176699 109651 176700
rect 110689 176699 110755 176700
rect 112253 176699 112319 176702
rect 118366 176700 118372 176702
rect 118436 176700 118483 176704
rect 125726 176700 125732 176764
rect 125796 176762 125802 176764
rect 125869 176762 125935 176765
rect 128169 176762 128235 176765
rect 133137 176764 133203 176765
rect 136081 176764 136147 176765
rect 148225 176764 148291 176765
rect 133086 176762 133092 176764
rect 125796 176760 125935 176762
rect 125796 176704 125874 176760
rect 125930 176704 125935 176760
rect 125796 176702 125935 176704
rect 125796 176700 125802 176702
rect 118417 176699 118483 176700
rect 125869 176699 125935 176702
rect 128126 176760 128235 176762
rect 128126 176704 128174 176760
rect 128230 176704 128235 176760
rect 128126 176699 128235 176704
rect 133046 176702 133092 176762
rect 133156 176760 133203 176764
rect 136030 176762 136036 176764
rect 133198 176704 133203 176760
rect 133086 176700 133092 176702
rect 133156 176700 133203 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 148174 176762 148180 176764
rect 136142 176704 136147 176760
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 158989 176762 159055 176765
rect 158916 176760 159055 176762
rect 158916 176704 158994 176760
rect 159050 176704 159055 176760
rect 158916 176702 159055 176704
rect 158916 176700 158922 176702
rect 133137 176699 133203 176700
rect 136081 176699 136147 176700
rect 148225 176699 148291 176700
rect 158989 176699 159055 176702
rect 103286 176492 103346 176699
rect 128126 176492 128186 176699
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect -960 175796 480 176036
rect 191741 175946 191807 175949
rect 240358 175946 240364 175948
rect 191741 175944 240364 175946
rect 191741 175888 191746 175944
rect 191802 175888 240364 175944
rect 191741 175886 240364 175888
rect 191741 175883 191807 175886
rect 240358 175884 240364 175886
rect 240428 175884 240434 175948
rect 273989 175946 274055 175949
rect 281574 175946 281580 175948
rect 273989 175944 281580 175946
rect 273989 175888 273994 175944
rect 274050 175888 281580 175944
rect 273989 175886 281580 175888
rect 273989 175883 274055 175886
rect 281574 175884 281580 175886
rect 281644 175884 281650 175948
rect 213913 175810 213979 175813
rect 227621 175810 227687 175813
rect 269757 175810 269823 175813
rect 213913 175808 217242 175810
rect 213913 175752 213918 175808
rect 213974 175752 217242 175808
rect 213913 175750 217242 175752
rect 213913 175747 213979 175750
rect 217182 175644 217242 175750
rect 227621 175808 228282 175810
rect 227621 175752 227626 175808
rect 227682 175752 228282 175808
rect 227621 175750 228282 175752
rect 227621 175747 227687 175750
rect 228222 175644 228282 175750
rect 269757 175808 279434 175810
rect 269757 175752 269762 175808
rect 269818 175752 279434 175808
rect 269757 175750 279434 175752
rect 269757 175747 269823 175750
rect 116945 175404 117011 175405
rect 120809 175404 120875 175405
rect 121913 175404 121979 175405
rect 134425 175404 134491 175405
rect 116894 175402 116900 175404
rect 116854 175342 116900 175402
rect 116964 175400 117011 175404
rect 120758 175402 120764 175404
rect 117006 175344 117011 175400
rect 116894 175340 116900 175342
rect 116964 175340 117011 175344
rect 120718 175342 120764 175402
rect 120828 175400 120875 175404
rect 121862 175402 121868 175404
rect 120870 175344 120875 175400
rect 120758 175340 120764 175342
rect 120828 175340 120875 175344
rect 121822 175342 121868 175402
rect 121932 175400 121979 175404
rect 134374 175402 134380 175404
rect 121974 175344 121979 175400
rect 121862 175340 121868 175342
rect 121932 175340 121979 175344
rect 134334 175342 134380 175402
rect 134444 175400 134491 175404
rect 134486 175344 134491 175400
rect 134374 175340 134380 175342
rect 134444 175340 134491 175344
rect 116945 175339 117011 175340
rect 120809 175339 120875 175340
rect 121913 175339 121979 175340
rect 134425 175339 134491 175340
rect 265801 175402 265867 175405
rect 268150 175402 268210 175644
rect 279374 175508 279434 175750
rect 265801 175400 268210 175402
rect 265801 175344 265806 175400
rect 265862 175344 268210 175400
rect 265801 175342 268210 175344
rect 265801 175339 265867 175342
rect 231761 175266 231827 175269
rect 228968 175264 231827 175266
rect 228968 175208 231766 175264
rect 231822 175208 231827 175264
rect 228968 175206 231827 175208
rect 231761 175203 231827 175206
rect 213913 175130 213979 175133
rect 213913 175128 217242 175130
rect 213913 175072 213918 175128
rect 213974 175072 217242 175128
rect 213913 175070 217242 175072
rect 213913 175067 213979 175070
rect 115749 174996 115815 174997
rect 115720 174994 115726 174996
rect 115658 174934 115726 174994
rect 115790 174992 115815 174996
rect 115810 174936 115815 174992
rect 217182 174964 217242 175070
rect 265341 174994 265407 174997
rect 268150 174994 268210 175236
rect 279366 175068 279372 175132
rect 279436 175068 279442 175132
rect 265341 174992 268210 174994
rect 115720 174932 115726 174934
rect 115790 174932 115815 174936
rect 115749 174931 115815 174932
rect 265341 174936 265346 174992
rect 265402 174936 268210 174992
rect 265341 174934 268210 174936
rect 265341 174931 265407 174934
rect 214005 174722 214071 174725
rect 231117 174722 231183 174725
rect 214005 174720 217242 174722
rect 214005 174664 214010 174720
rect 214066 174664 217242 174720
rect 214005 174662 217242 174664
rect 228968 174720 231183 174722
rect 228968 174664 231122 174720
rect 231178 174664 231183 174720
rect 228968 174662 231183 174664
rect 214005 174659 214071 174662
rect 217182 174284 217242 174662
rect 231117 174659 231183 174662
rect 265801 174586 265867 174589
rect 268150 174586 268210 174828
rect 279374 174692 279434 175068
rect 265801 174584 268210 174586
rect 265801 174528 265806 174584
rect 265862 174528 268210 174584
rect 265801 174526 268210 174528
rect 265801 174523 265867 174526
rect 279417 174450 279483 174453
rect 279374 174448 279483 174450
rect 229134 174314 229140 174316
rect 228968 174254 229140 174314
rect 229134 174252 229140 174254
rect 229204 174252 229210 174316
rect 265617 174178 265683 174181
rect 268150 174178 268210 174420
rect 265617 174176 268210 174178
rect 265617 174120 265622 174176
rect 265678 174120 268210 174176
rect 265617 174118 268210 174120
rect 279374 174392 279422 174448
rect 279478 174392 279483 174448
rect 279374 174387 279483 174392
rect 265617 174115 265683 174118
rect 265893 174042 265959 174045
rect 265893 174040 267842 174042
rect 265893 173984 265898 174040
rect 265954 173984 267842 174040
rect 279374 174012 279434 174387
rect 265893 173982 267842 173984
rect 265893 173979 265959 173982
rect 213913 173770 213979 173773
rect 231669 173770 231735 173773
rect 213913 173768 217242 173770
rect 213913 173712 213918 173768
rect 213974 173712 217242 173768
rect 213913 173710 217242 173712
rect 228968 173768 231735 173770
rect 228968 173712 231674 173768
rect 231730 173712 231735 173768
rect 228968 173710 231735 173712
rect 267782 173770 267842 173982
rect 268334 173770 268394 174012
rect 267782 173710 268394 173770
rect 279325 173770 279391 173773
rect 279325 173768 279434 173770
rect 279325 173712 279330 173768
rect 279386 173712 279434 173768
rect 213913 173707 213979 173710
rect 217182 173604 217242 173710
rect 231669 173707 231735 173710
rect 279325 173707 279434 173712
rect 214005 173362 214071 173365
rect 231209 173362 231275 173365
rect 214005 173360 217242 173362
rect 214005 173304 214010 173360
rect 214066 173304 217242 173360
rect 214005 173302 217242 173304
rect 228968 173360 231275 173362
rect 228968 173304 231214 173360
rect 231270 173304 231275 173360
rect 228968 173302 231275 173304
rect 214005 173299 214071 173302
rect 165337 173226 165403 173229
rect 214414 173226 214420 173228
rect 165337 173224 214420 173226
rect 165337 173168 165342 173224
rect 165398 173168 214420 173224
rect 165337 173166 214420 173168
rect 165337 173163 165403 173166
rect 214414 173164 214420 173166
rect 214484 173164 214490 173228
rect 217182 172924 217242 173302
rect 231209 173299 231275 173302
rect 265709 173226 265775 173229
rect 268150 173226 268210 173604
rect 265709 173224 268210 173226
rect 265709 173168 265714 173224
rect 265770 173168 268210 173224
rect 279374 173196 279434 173707
rect 265709 173166 268210 173168
rect 265709 173163 265775 173166
rect 231761 172818 231827 172821
rect 228968 172816 231827 172818
rect 228968 172760 231766 172816
rect 231822 172760 231827 172816
rect 228968 172758 231827 172760
rect 231761 172755 231827 172758
rect 265893 172818 265959 172821
rect 268150 172818 268210 173060
rect 265893 172816 268210 172818
rect 265893 172760 265898 172816
rect 265954 172760 268210 172816
rect 265893 172758 268210 172760
rect 265893 172755 265959 172758
rect 265801 172546 265867 172549
rect 265801 172544 267842 172546
rect 265801 172488 265806 172544
rect 265862 172488 267842 172544
rect 265801 172486 267842 172488
rect 265801 172483 265867 172486
rect 214189 172410 214255 172413
rect 231761 172410 231827 172413
rect 214189 172408 217242 172410
rect 214189 172352 214194 172408
rect 214250 172352 217242 172408
rect 214189 172350 217242 172352
rect 228968 172408 231827 172410
rect 228968 172352 231766 172408
rect 231822 172352 231827 172408
rect 228968 172350 231827 172352
rect 267782 172410 267842 172486
rect 268334 172410 268394 172652
rect 280337 172410 280403 172413
rect 267782 172350 268394 172410
rect 279956 172408 280403 172410
rect 279956 172352 280342 172408
rect 280398 172352 280403 172408
rect 279956 172350 280403 172352
rect 214189 172347 214255 172350
rect 217182 172244 217242 172350
rect 231761 172347 231827 172350
rect 280337 172347 280403 172350
rect 214097 172002 214163 172005
rect 265341 172002 265407 172005
rect 268150 172002 268210 172244
rect 214097 172000 217242 172002
rect 214097 171944 214102 172000
rect 214158 171944 217242 172000
rect 214097 171942 217242 171944
rect 214097 171939 214163 171942
rect 168005 171594 168071 171597
rect 164694 171592 168071 171594
rect 164694 171536 168010 171592
rect 168066 171536 168071 171592
rect 217182 171564 217242 171942
rect 265341 172000 268210 172002
rect 265341 171944 265346 172000
rect 265402 171944 268210 172000
rect 265341 171942 268210 171944
rect 265341 171939 265407 171942
rect 231669 171866 231735 171869
rect 228968 171864 231735 171866
rect 228968 171808 231674 171864
rect 231730 171808 231735 171864
rect 228968 171806 231735 171808
rect 231669 171803 231735 171806
rect 265801 171594 265867 171597
rect 268150 171594 268210 171836
rect 265801 171592 268210 171594
rect 164694 171534 168071 171536
rect 168005 171531 168071 171534
rect 265801 171536 265806 171592
rect 265862 171536 268210 171592
rect 265801 171534 268210 171536
rect 265801 171531 265867 171534
rect 231669 171458 231735 171461
rect 228968 171456 231735 171458
rect 228968 171400 231674 171456
rect 231730 171400 231735 171456
rect 228968 171398 231735 171400
rect 231669 171395 231735 171398
rect 265893 171186 265959 171189
rect 268334 171186 268394 171428
rect 265893 171184 268394 171186
rect 265893 171128 265898 171184
rect 265954 171128 268394 171184
rect 265893 171126 268394 171128
rect 279926 171186 279986 171700
rect 296621 171188 296687 171189
rect 295558 171186 295564 171188
rect 279926 171126 295564 171186
rect 265893 171123 265959 171126
rect 295558 171124 295564 171126
rect 295628 171124 295634 171188
rect 296621 171186 296668 171188
rect 296576 171184 296668 171186
rect 296732 171186 296738 171188
rect 296576 171128 296626 171184
rect 296576 171126 296668 171128
rect 296621 171124 296668 171126
rect 296732 171126 296814 171186
rect 296732 171124 296738 171126
rect 296621 171123 296687 171124
rect 213913 170778 213979 170781
rect 217366 170778 217426 171020
rect 231761 170914 231827 170917
rect 228968 170912 231827 170914
rect 228968 170856 231766 170912
rect 231822 170856 231827 170912
rect 228968 170854 231827 170856
rect 231761 170851 231827 170854
rect 213913 170776 217426 170778
rect 213913 170720 213918 170776
rect 213974 170720 217426 170776
rect 213913 170718 217426 170720
rect 213913 170715 213979 170718
rect 214005 170642 214071 170645
rect 265341 170642 265407 170645
rect 268150 170642 268210 171020
rect 282821 170914 282887 170917
rect 279956 170912 282887 170914
rect 279956 170856 282826 170912
rect 282882 170856 282887 170912
rect 279956 170854 282887 170856
rect 282821 170851 282887 170854
rect 214005 170640 217242 170642
rect 214005 170584 214010 170640
rect 214066 170584 217242 170640
rect 214005 170582 217242 170584
rect 214005 170579 214071 170582
rect 217182 170340 217242 170582
rect 265341 170640 268210 170642
rect 265341 170584 265346 170640
rect 265402 170584 268210 170640
rect 265341 170582 268210 170584
rect 265341 170579 265407 170582
rect 231761 170506 231827 170509
rect 228968 170504 231827 170506
rect 228968 170448 231766 170504
rect 231822 170448 231827 170504
rect 228968 170446 231827 170448
rect 231761 170443 231827 170446
rect 264237 170234 264303 170237
rect 268150 170234 268210 170476
rect 264237 170232 268210 170234
rect 264237 170176 264242 170232
rect 264298 170176 268210 170232
rect 264237 170174 268210 170176
rect 264237 170171 264303 170174
rect 282729 170098 282795 170101
rect 279956 170096 282795 170098
rect 231301 169962 231367 169965
rect 228968 169960 231367 169962
rect 228968 169904 231306 169960
rect 231362 169904 231367 169960
rect 228968 169902 231367 169904
rect 231301 169899 231367 169902
rect 265617 169826 265683 169829
rect 268150 169826 268210 170068
rect 279956 170040 282734 170096
rect 282790 170040 282795 170096
rect 279956 170038 282795 170040
rect 282729 170035 282795 170038
rect 265617 169824 268210 169826
rect 265617 169768 265622 169824
rect 265678 169768 268210 169824
rect 265617 169766 268210 169768
rect 265617 169763 265683 169766
rect 213913 169418 213979 169421
rect 217366 169418 217426 169660
rect 231669 169554 231735 169557
rect 228968 169552 231735 169554
rect 228968 169496 231674 169552
rect 231730 169496 231735 169552
rect 228968 169494 231735 169496
rect 231669 169491 231735 169494
rect 213913 169416 217426 169418
rect 213913 169360 213918 169416
rect 213974 169360 217426 169416
rect 213913 169358 217426 169360
rect 265433 169418 265499 169421
rect 268150 169418 268210 169660
rect 282821 169418 282887 169421
rect 265433 169416 268210 169418
rect 265433 169360 265438 169416
rect 265494 169360 268210 169416
rect 265433 169358 268210 169360
rect 279956 169416 282887 169418
rect 279956 169360 282826 169416
rect 282882 169360 282887 169416
rect 279956 169358 282887 169360
rect 213913 169355 213979 169358
rect 265433 169355 265499 169358
rect 282821 169355 282887 169358
rect 214005 169282 214071 169285
rect 214005 169280 217242 169282
rect 214005 169224 214010 169280
rect 214066 169224 217242 169280
rect 214005 169222 217242 169224
rect 214005 169219 214071 169222
rect 217182 168980 217242 169222
rect 229185 169010 229251 169013
rect 228968 169008 229251 169010
rect 228968 168952 229190 169008
rect 229246 168952 229251 169008
rect 228968 168950 229251 168952
rect 229185 168947 229251 168950
rect 265341 169010 265407 169013
rect 268150 169010 268210 169252
rect 265341 169008 268210 169010
rect 265341 168952 265346 169008
rect 265402 168952 268210 169008
rect 265341 168950 268210 168952
rect 265341 168947 265407 168950
rect 231761 168602 231827 168605
rect 228968 168600 231827 168602
rect 228968 168544 231766 168600
rect 231822 168544 231827 168600
rect 228968 168542 231827 168544
rect 231761 168539 231827 168542
rect 265801 168602 265867 168605
rect 268518 168604 268578 168844
rect 265801 168600 268210 168602
rect 265801 168544 265806 168600
rect 265862 168544 268210 168600
rect 265801 168542 268210 168544
rect 265801 168539 265867 168542
rect 268150 168436 268210 168542
rect 268510 168540 268516 168604
rect 268580 168540 268586 168604
rect 281717 168602 281783 168605
rect 279956 168600 281783 168602
rect 279956 168544 281722 168600
rect 281778 168544 281783 168600
rect 279956 168542 281783 168544
rect 281717 168539 281783 168542
rect 213913 168058 213979 168061
rect 217366 168058 217426 168300
rect 264421 168194 264487 168197
rect 268510 168194 268516 168196
rect 264421 168192 268516 168194
rect 264421 168136 264426 168192
rect 264482 168136 268516 168192
rect 264421 168134 268516 168136
rect 264421 168131 264487 168134
rect 268510 168132 268516 168134
rect 268580 168132 268586 168196
rect 231761 168058 231827 168061
rect 213913 168056 217426 168058
rect 213913 168000 213918 168056
rect 213974 168000 217426 168056
rect 213913 167998 217426 168000
rect 228968 168056 231827 168058
rect 228968 168000 231766 168056
rect 231822 168000 231827 168056
rect 228968 167998 231827 168000
rect 213913 167995 213979 167998
rect 231761 167995 231827 167998
rect 214005 167922 214071 167925
rect 214005 167920 217242 167922
rect 214005 167864 214010 167920
rect 214066 167864 217242 167920
rect 214005 167862 217242 167864
rect 214005 167859 214071 167862
rect 217182 167620 217242 167862
rect 231669 167650 231735 167653
rect 228968 167648 231735 167650
rect 228968 167592 231674 167648
rect 231730 167592 231735 167648
rect 228968 167590 231735 167592
rect 231669 167587 231735 167590
rect 265157 167650 265223 167653
rect 268150 167650 268210 167892
rect 281625 167786 281691 167789
rect 279956 167784 281691 167786
rect 279956 167728 281630 167784
rect 281686 167728 281691 167784
rect 279956 167726 281691 167728
rect 281625 167723 281691 167726
rect 265157 167648 268210 167650
rect 265157 167592 265162 167648
rect 265218 167592 268210 167648
rect 265157 167590 268210 167592
rect 265157 167587 265223 167590
rect 265801 167242 265867 167245
rect 268518 167244 268578 167484
rect 265801 167240 268210 167242
rect 265801 167184 265806 167240
rect 265862 167184 268210 167240
rect 265801 167182 268210 167184
rect 265801 167179 265867 167182
rect 231577 167106 231643 167109
rect 216998 167046 217242 167106
rect 228968 167104 231643 167106
rect 228968 167048 231582 167104
rect 231638 167048 231643 167104
rect 268150 167076 268210 167182
rect 268510 167180 268516 167244
rect 268580 167180 268586 167244
rect 282453 167106 282519 167109
rect 279956 167104 282519 167106
rect 228968 167046 231643 167048
rect 279956 167048 282458 167104
rect 282514 167048 282519 167104
rect 279956 167046 282519 167048
rect 213269 166970 213335 166973
rect 216998 166970 217058 167046
rect 213269 166968 217058 166970
rect 213269 166912 213274 166968
rect 213330 166912 217058 166968
rect 217182 166940 217242 167046
rect 231577 167043 231643 167046
rect 282453 167043 282519 167046
rect 213269 166910 217058 166912
rect 213269 166907 213335 166910
rect 261385 166834 261451 166837
rect 268510 166834 268516 166836
rect 261385 166832 268516 166834
rect 261385 166776 261390 166832
rect 261446 166776 268516 166832
rect 261385 166774 268516 166776
rect 261385 166771 261451 166774
rect 268510 166772 268516 166774
rect 268580 166772 268586 166836
rect 213913 166698 213979 166701
rect 231761 166698 231827 166701
rect 213913 166696 217242 166698
rect 213913 166640 213918 166696
rect 213974 166640 217242 166696
rect 213913 166638 217242 166640
rect 228968 166696 231827 166698
rect 228968 166640 231766 166696
rect 231822 166640 231827 166696
rect 228968 166638 231827 166640
rect 213913 166635 213979 166638
rect 217182 166396 217242 166638
rect 231761 166635 231827 166638
rect 265985 166426 266051 166429
rect 268150 166426 268210 166668
rect 265985 166424 268210 166426
rect 265985 166368 265990 166424
rect 266046 166368 268210 166424
rect 265985 166366 268210 166368
rect 265985 166363 266051 166366
rect 282085 166290 282151 166293
rect 279956 166288 282151 166290
rect 214005 166154 214071 166157
rect 231117 166154 231183 166157
rect 214005 166152 217242 166154
rect 214005 166096 214010 166152
rect 214066 166096 217242 166152
rect 214005 166094 217242 166096
rect 228968 166152 231183 166154
rect 228968 166096 231122 166152
rect 231178 166096 231183 166152
rect 228968 166094 231183 166096
rect 214005 166091 214071 166094
rect 217182 165716 217242 166094
rect 231117 166091 231183 166094
rect 265709 166018 265775 166021
rect 268150 166018 268210 166260
rect 279956 166232 282090 166288
rect 282146 166232 282151 166288
rect 279956 166230 282151 166232
rect 282085 166227 282151 166230
rect 265709 166016 268210 166018
rect 265709 165960 265714 166016
rect 265770 165960 268210 166016
rect 265709 165958 268210 165960
rect 265709 165955 265775 165958
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 231485 165746 231551 165749
rect 228968 165744 231551 165746
rect 228968 165688 231490 165744
rect 231546 165688 231551 165744
rect 228968 165686 231551 165688
rect 231485 165683 231551 165686
rect 265801 165746 265867 165749
rect 265801 165744 267842 165746
rect 265801 165688 265806 165744
rect 265862 165688 267842 165744
rect 265801 165686 267842 165688
rect 265801 165683 265867 165686
rect 267782 165610 267842 165686
rect 268334 165610 268394 165852
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 267782 165550 268394 165610
rect 214649 165474 214715 165477
rect 282821 165474 282887 165477
rect 214649 165472 217242 165474
rect 214649 165416 214654 165472
rect 214710 165416 217242 165472
rect 214649 165414 217242 165416
rect 279956 165472 282887 165474
rect 279956 165416 282826 165472
rect 282882 165416 282887 165472
rect 279956 165414 282887 165416
rect 214649 165411 214715 165414
rect 217182 165036 217242 165414
rect 282821 165411 282887 165414
rect 231761 165202 231827 165205
rect 228968 165200 231827 165202
rect 228968 165144 231766 165200
rect 231822 165144 231827 165200
rect 228968 165142 231827 165144
rect 231761 165139 231827 165142
rect 265433 165066 265499 165069
rect 268150 165066 268210 165308
rect 265433 165064 268210 165066
rect 265433 165008 265438 165064
rect 265494 165008 268210 165064
rect 265433 165006 268210 165008
rect 265433 165003 265499 165006
rect 213913 164794 213979 164797
rect 231301 164794 231367 164797
rect 213913 164792 217242 164794
rect 213913 164736 213918 164792
rect 213974 164736 217242 164792
rect 213913 164734 217242 164736
rect 228968 164792 231367 164794
rect 228968 164736 231306 164792
rect 231362 164736 231367 164792
rect 228968 164734 231367 164736
rect 213913 164731 213979 164734
rect 217182 164356 217242 164734
rect 231301 164731 231367 164734
rect 265709 164658 265775 164661
rect 268150 164658 268210 164900
rect 281993 164794 282059 164797
rect 279956 164792 282059 164794
rect 279956 164736 281998 164792
rect 282054 164736 282059 164792
rect 279956 164734 282059 164736
rect 281993 164731 282059 164734
rect 265709 164656 268210 164658
rect 265709 164600 265714 164656
rect 265770 164600 268210 164656
rect 265709 164598 268210 164600
rect 265709 164595 265775 164598
rect 230657 164386 230723 164389
rect 228968 164384 230723 164386
rect 228968 164328 230662 164384
rect 230718 164328 230723 164384
rect 228968 164326 230723 164328
rect 230657 164323 230723 164326
rect 265801 164250 265867 164253
rect 268334 164250 268394 164492
rect 265801 164248 268394 164250
rect 265801 164192 265806 164248
rect 265862 164192 268394 164248
rect 265801 164190 268394 164192
rect 265801 164187 265867 164190
rect 214465 164114 214531 164117
rect 214465 164112 217242 164114
rect 214465 164056 214470 164112
rect 214526 164056 217242 164112
rect 214465 164054 217242 164056
rect 214465 164051 214531 164054
rect 217182 163676 217242 164054
rect 236494 163842 236500 163844
rect 228968 163782 236500 163842
rect 236494 163780 236500 163782
rect 236564 163780 236570 163844
rect 265893 163842 265959 163845
rect 268150 163842 268210 164084
rect 282085 163978 282151 163981
rect 279956 163976 282151 163978
rect 279956 163920 282090 163976
rect 282146 163920 282151 163976
rect 279956 163918 282151 163920
rect 282085 163915 282151 163918
rect 265893 163840 268210 163842
rect 265893 163784 265898 163840
rect 265954 163784 268210 163840
rect 265893 163782 268210 163784
rect 265893 163779 265959 163782
rect 213913 163434 213979 163437
rect 234654 163434 234660 163436
rect 213913 163432 217242 163434
rect 213913 163376 213918 163432
rect 213974 163376 217242 163432
rect 213913 163374 217242 163376
rect 228968 163374 234660 163434
rect 213913 163371 213979 163374
rect 217182 162996 217242 163374
rect 234654 163372 234660 163374
rect 234724 163372 234730 163436
rect 265525 163434 265591 163437
rect 268150 163434 268210 163676
rect 265525 163432 268210 163434
rect 265525 163376 265530 163432
rect 265586 163376 268210 163432
rect 265525 163374 268210 163376
rect 265525 163371 265591 163374
rect 265341 163026 265407 163029
rect 268150 163026 268210 163268
rect 282821 163162 282887 163165
rect 279956 163160 282887 163162
rect 279956 163104 282826 163160
rect 282882 163104 282887 163160
rect 279956 163102 282887 163104
rect 282821 163099 282887 163102
rect 265341 163024 268210 163026
rect -960 162890 480 162980
rect 265341 162968 265346 163024
rect 265402 162968 268210 163024
rect 265341 162966 268210 162968
rect 265341 162963 265407 162966
rect 3417 162890 3483 162893
rect 231669 162890 231735 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect 228968 162888 231735 162890
rect 228968 162832 231674 162888
rect 231730 162832 231735 162888
rect 228968 162830 231735 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 231669 162827 231735 162830
rect 265801 162890 265867 162893
rect 265801 162888 267842 162890
rect 265801 162832 265806 162888
rect 265862 162832 267842 162888
rect 265801 162830 267842 162832
rect 265801 162827 265867 162830
rect 213913 162618 213979 162621
rect 267782 162618 267842 162830
rect 268334 162618 268394 162860
rect 213913 162616 217242 162618
rect 213913 162560 213918 162616
rect 213974 162560 217242 162616
rect 213913 162558 217242 162560
rect 267782 162558 268394 162618
rect 213913 162555 213979 162558
rect 217182 162316 217242 162558
rect 231761 162482 231827 162485
rect 282085 162482 282151 162485
rect 228968 162480 231827 162482
rect 228968 162424 231766 162480
rect 231822 162424 231827 162480
rect 228968 162422 231827 162424
rect 279956 162480 282151 162482
rect 279956 162424 282090 162480
rect 282146 162424 282151 162480
rect 279956 162422 282151 162424
rect 231761 162419 231827 162422
rect 282085 162419 282151 162422
rect 213177 162074 213243 162077
rect 265341 162074 265407 162077
rect 268150 162074 268210 162316
rect 213177 162072 217242 162074
rect 213177 162016 213182 162072
rect 213238 162016 217242 162072
rect 213177 162014 217242 162016
rect 213177 162011 213243 162014
rect 217182 161772 217242 162014
rect 265341 162072 268210 162074
rect 265341 162016 265346 162072
rect 265402 162016 268210 162072
rect 265341 162014 268210 162016
rect 265341 162011 265407 162014
rect 231761 161938 231827 161941
rect 228968 161936 231827 161938
rect 228968 161880 231766 161936
rect 231822 161880 231827 161936
rect 228968 161878 231827 161880
rect 231761 161875 231827 161878
rect 265801 161666 265867 161669
rect 268518 161668 268578 161908
rect 265801 161664 268210 161666
rect 265801 161608 265806 161664
rect 265862 161608 268210 161664
rect 265801 161606 268210 161608
rect 265801 161603 265867 161606
rect 231669 161530 231735 161533
rect 228968 161528 231735 161530
rect 228968 161472 231674 161528
rect 231730 161472 231735 161528
rect 268150 161500 268210 161606
rect 268510 161604 268516 161668
rect 268580 161604 268586 161668
rect 282821 161666 282887 161669
rect 279956 161664 282887 161666
rect 279956 161608 282826 161664
rect 282882 161608 282887 161664
rect 279956 161606 282887 161608
rect 282821 161603 282887 161606
rect 228968 161470 231735 161472
rect 231669 161467 231735 161470
rect 213913 161394 213979 161397
rect 213913 161392 217242 161394
rect 213913 161336 213918 161392
rect 213974 161336 217242 161392
rect 213913 161334 217242 161336
rect 213913 161331 213979 161334
rect 217182 161092 217242 161334
rect 231761 160986 231827 160989
rect 228968 160984 231827 160986
rect 228968 160928 231766 160984
rect 231822 160928 231827 160984
rect 228968 160926 231827 160928
rect 231761 160923 231827 160926
rect 214414 160788 214420 160852
rect 214484 160850 214490 160852
rect 265341 160850 265407 160853
rect 268150 160850 268210 161092
rect 282821 160850 282887 160853
rect 214484 160790 217242 160850
rect 214484 160788 214490 160790
rect 217182 160412 217242 160790
rect 265341 160848 268210 160850
rect 265341 160792 265346 160848
rect 265402 160792 268210 160848
rect 265341 160790 268210 160792
rect 279956 160848 282887 160850
rect 279956 160792 282826 160848
rect 282882 160792 282887 160848
rect 279956 160790 282887 160792
rect 265341 160787 265407 160790
rect 282821 160787 282887 160790
rect 231393 160578 231459 160581
rect 228968 160576 231459 160578
rect 228968 160520 231398 160576
rect 231454 160520 231459 160576
rect 228968 160518 231459 160520
rect 231393 160515 231459 160518
rect 265617 160442 265683 160445
rect 268150 160442 268210 160684
rect 265617 160440 268210 160442
rect 265617 160384 265622 160440
rect 265678 160384 268210 160440
rect 265617 160382 268210 160384
rect 265617 160379 265683 160382
rect 265801 160170 265867 160173
rect 265801 160168 267842 160170
rect 265801 160112 265806 160168
rect 265862 160112 267842 160168
rect 265801 160110 267842 160112
rect 265801 160107 265867 160110
rect 213913 160034 213979 160037
rect 250294 160034 250300 160036
rect 213913 160032 217242 160034
rect 213913 159976 213918 160032
rect 213974 159976 217242 160032
rect 213913 159974 217242 159976
rect 228968 159974 250300 160034
rect 213913 159971 213979 159974
rect 217182 159732 217242 159974
rect 250294 159972 250300 159974
rect 250364 159972 250370 160036
rect 267782 160034 267842 160110
rect 268334 160034 268394 160276
rect 281533 160170 281599 160173
rect 279956 160168 281599 160170
rect 279956 160112 281538 160168
rect 281594 160112 281599 160168
rect 279956 160110 281599 160112
rect 281533 160107 281599 160110
rect 267782 159974 268394 160034
rect 231761 159626 231827 159629
rect 228968 159624 231827 159626
rect 228968 159568 231766 159624
rect 231822 159568 231827 159624
rect 228968 159566 231827 159568
rect 231761 159563 231827 159566
rect 214005 159490 214071 159493
rect 265341 159490 265407 159493
rect 268150 159490 268210 159732
rect 214005 159488 217242 159490
rect 214005 159432 214010 159488
rect 214066 159432 217242 159488
rect 214005 159430 217242 159432
rect 214005 159427 214071 159430
rect 217182 159052 217242 159430
rect 265341 159488 268210 159490
rect 265341 159432 265346 159488
rect 265402 159432 268210 159488
rect 265341 159430 268210 159432
rect 265341 159427 265407 159430
rect 281533 159354 281599 159357
rect 279956 159352 281599 159354
rect 231485 159082 231551 159085
rect 228968 159080 231551 159082
rect 228968 159024 231490 159080
rect 231546 159024 231551 159080
rect 228968 159022 231551 159024
rect 231485 159019 231551 159022
rect 265617 159082 265683 159085
rect 268150 159082 268210 159324
rect 279956 159296 281538 159352
rect 281594 159296 281599 159352
rect 279956 159294 281599 159296
rect 281533 159291 281599 159294
rect 265617 159080 268210 159082
rect 265617 159024 265622 159080
rect 265678 159024 268210 159080
rect 265617 159022 268210 159024
rect 265617 159019 265683 159022
rect 265801 158810 265867 158813
rect 265801 158808 267842 158810
rect 265801 158752 265806 158808
rect 265862 158752 267842 158808
rect 265801 158750 267842 158752
rect 265801 158747 265867 158750
rect 213913 158674 213979 158677
rect 230657 158674 230723 158677
rect 213913 158672 217242 158674
rect 213913 158616 213918 158672
rect 213974 158616 217242 158672
rect 213913 158614 217242 158616
rect 228968 158672 230723 158674
rect 228968 158616 230662 158672
rect 230718 158616 230723 158672
rect 228968 158614 230723 158616
rect 267782 158674 267842 158750
rect 268334 158674 268394 158916
rect 267782 158614 268394 158674
rect 213913 158611 213979 158614
rect 217182 158372 217242 158614
rect 230657 158611 230723 158614
rect 282821 158538 282887 158541
rect 279956 158536 282887 158538
rect 265617 158266 265683 158269
rect 268150 158266 268210 158508
rect 279956 158480 282826 158536
rect 282882 158480 282887 158536
rect 279956 158478 282887 158480
rect 282821 158475 282887 158478
rect 265617 158264 268210 158266
rect 265617 158208 265622 158264
rect 265678 158208 268210 158264
rect 265617 158206 268210 158208
rect 265617 158203 265683 158206
rect 214097 158130 214163 158133
rect 231761 158130 231827 158133
rect 214097 158128 217242 158130
rect 214097 158072 214102 158128
rect 214158 158072 217242 158128
rect 214097 158070 217242 158072
rect 228968 158128 231827 158130
rect 228968 158072 231766 158128
rect 231822 158072 231827 158128
rect 228968 158070 231827 158072
rect 214097 158067 214163 158070
rect 217182 157692 217242 158070
rect 231761 158067 231827 158070
rect 265249 157858 265315 157861
rect 268150 157858 268210 158100
rect 282729 157858 282795 157861
rect 265249 157856 268210 157858
rect 265249 157800 265254 157856
rect 265310 157800 268210 157856
rect 265249 157798 268210 157800
rect 279956 157856 282795 157858
rect 279956 157800 282734 157856
rect 282790 157800 282795 157856
rect 279956 157798 282795 157800
rect 265249 157795 265315 157798
rect 282729 157795 282795 157798
rect 230749 157722 230815 157725
rect 228968 157720 230815 157722
rect 228968 157664 230754 157720
rect 230810 157664 230815 157720
rect 228968 157662 230815 157664
rect 230749 157659 230815 157662
rect 265525 157450 265591 157453
rect 268150 157450 268210 157692
rect 265525 157448 268210 157450
rect 265525 157392 265530 157448
rect 265586 157392 268210 157448
rect 265525 157390 268210 157392
rect 265525 157387 265591 157390
rect 261661 157314 261727 157317
rect 268510 157314 268516 157316
rect 200070 157254 217242 157314
rect 166390 156028 166396 156092
rect 166460 156090 166466 156092
rect 200070 156090 200130 157254
rect 217182 157148 217242 157254
rect 261661 157312 268516 157314
rect 261661 157256 261666 157312
rect 261722 157256 268516 157312
rect 261661 157254 268516 157256
rect 261661 157251 261727 157254
rect 268510 157252 268516 157254
rect 268580 157252 268586 157316
rect 231761 157178 231827 157181
rect 228968 157176 231827 157178
rect 228968 157120 231766 157176
rect 231822 157120 231827 157176
rect 228968 157118 231827 157120
rect 231761 157115 231827 157118
rect 213913 156906 213979 156909
rect 265893 156906 265959 156909
rect 268150 156906 268210 157148
rect 281574 157042 281580 157044
rect 279956 156982 281580 157042
rect 281574 156980 281580 156982
rect 281644 156980 281650 157044
rect 213913 156904 217242 156906
rect 213913 156848 213918 156904
rect 213974 156848 217242 156904
rect 213913 156846 217242 156848
rect 213913 156843 213979 156846
rect 217182 156468 217242 156846
rect 265893 156904 268210 156906
rect 265893 156848 265898 156904
rect 265954 156848 268210 156904
rect 265893 156846 268210 156848
rect 265893 156843 265959 156846
rect 231669 156770 231735 156773
rect 228968 156768 231735 156770
rect 228968 156712 231674 156768
rect 231730 156712 231735 156768
rect 228968 156710 231735 156712
rect 231669 156707 231735 156710
rect 265525 156498 265591 156501
rect 268150 156498 268210 156740
rect 265525 156496 268210 156498
rect 265525 156440 265530 156496
rect 265586 156440 268210 156496
rect 265525 156438 268210 156440
rect 265525 156435 265591 156438
rect 281717 156362 281783 156365
rect 279956 156360 281783 156362
rect 230933 156226 230999 156229
rect 228968 156224 230999 156226
rect 228968 156168 230938 156224
rect 230994 156168 230999 156224
rect 228968 156166 230999 156168
rect 230933 156163 230999 156166
rect 166460 156030 200130 156090
rect 265801 156090 265867 156093
rect 268150 156090 268210 156332
rect 279956 156304 281722 156360
rect 281778 156304 281783 156360
rect 279956 156302 281783 156304
rect 281717 156299 281783 156302
rect 265801 156088 268210 156090
rect 265801 156032 265806 156088
rect 265862 156032 268210 156088
rect 265801 156030 268210 156032
rect 166460 156028 166466 156030
rect 265801 156027 265867 156030
rect 200070 155894 217242 155954
rect 166206 154532 166212 154596
rect 166276 154594 166282 154596
rect 200070 154594 200130 155894
rect 217182 155788 217242 155894
rect 231117 155818 231183 155821
rect 228968 155816 231183 155818
rect 228968 155760 231122 155816
rect 231178 155760 231183 155816
rect 228968 155758 231183 155760
rect 231117 155755 231183 155758
rect 265801 155682 265867 155685
rect 268150 155682 268210 155924
rect 265801 155680 268210 155682
rect 265801 155624 265806 155680
rect 265862 155624 268210 155680
rect 265801 155622 268210 155624
rect 265801 155619 265867 155622
rect 213913 155546 213979 155549
rect 283097 155546 283163 155549
rect 213913 155544 217242 155546
rect 213913 155488 213918 155544
rect 213974 155488 217242 155544
rect 279956 155544 283163 155546
rect 213913 155486 217242 155488
rect 213913 155483 213979 155486
rect 217182 155108 217242 155486
rect 230565 155274 230631 155277
rect 228968 155272 230631 155274
rect 228968 155216 230570 155272
rect 230626 155216 230631 155272
rect 228968 155214 230631 155216
rect 230565 155211 230631 155214
rect 231577 155274 231643 155277
rect 251214 155274 251220 155276
rect 231577 155272 251220 155274
rect 231577 155216 231582 155272
rect 231638 155216 251220 155272
rect 231577 155214 251220 155216
rect 231577 155211 231643 155214
rect 251214 155212 251220 155214
rect 251284 155212 251290 155276
rect 265709 155274 265775 155277
rect 268150 155274 268210 155516
rect 279956 155488 283102 155544
rect 283158 155488 283163 155544
rect 279956 155486 283163 155488
rect 283097 155483 283163 155486
rect 265709 155272 268210 155274
rect 265709 155216 265714 155272
rect 265770 155216 268210 155272
rect 265709 155214 268210 155216
rect 265709 155211 265775 155214
rect 231761 154866 231827 154869
rect 228968 154864 231827 154866
rect 228968 154808 231766 154864
rect 231822 154808 231827 154864
rect 228968 154806 231827 154808
rect 231761 154803 231827 154806
rect 265985 154730 266051 154733
rect 268518 154730 268578 155108
rect 281625 154730 281691 154733
rect 265985 154728 268578 154730
rect 265985 154672 265990 154728
rect 266046 154672 268578 154728
rect 265985 154670 268578 154672
rect 279956 154728 281691 154730
rect 279956 154672 281630 154728
rect 281686 154672 281691 154728
rect 279956 154670 281691 154672
rect 265985 154667 266051 154670
rect 281625 154667 281691 154670
rect 166276 154534 200130 154594
rect 266077 154594 266143 154597
rect 266077 154592 267842 154594
rect 266077 154536 266082 154592
rect 266138 154536 267842 154592
rect 266077 154534 267842 154536
rect 166276 154532 166282 154534
rect 266077 154531 266143 154534
rect 214005 153914 214071 153917
rect 217182 153914 217242 154428
rect 229093 154322 229159 154325
rect 228968 154320 229159 154322
rect 228968 154264 229098 154320
rect 229154 154264 229159 154320
rect 228968 154262 229159 154264
rect 267782 154322 267842 154534
rect 268334 154322 268394 154564
rect 267782 154262 268394 154322
rect 229093 154259 229159 154262
rect 237414 153914 237420 153916
rect 214005 153912 217242 153914
rect 214005 153856 214010 153912
rect 214066 153856 217242 153912
rect 214005 153854 217242 153856
rect 228968 153854 237420 153914
rect 214005 153851 214071 153854
rect 237414 153852 237420 153854
rect 237484 153852 237490 153916
rect 265893 153914 265959 153917
rect 268150 153914 268210 154156
rect 281717 154050 281783 154053
rect 279956 154048 281783 154050
rect 279956 153992 281722 154048
rect 281778 153992 281783 154048
rect 279956 153990 281783 153992
rect 281717 153987 281783 153990
rect 265893 153912 268210 153914
rect 265893 153856 265898 153912
rect 265954 153856 268210 153912
rect 265893 153854 268210 153856
rect 265893 153851 265959 153854
rect 213913 153370 213979 153373
rect 217182 153370 217242 153748
rect 265801 153506 265867 153509
rect 268150 153506 268210 153748
rect 265801 153504 268210 153506
rect 265801 153448 265806 153504
rect 265862 153448 268210 153504
rect 265801 153446 268210 153448
rect 265801 153443 265867 153446
rect 231945 153370 232011 153373
rect 213913 153368 217242 153370
rect 213913 153312 213918 153368
rect 213974 153312 217242 153368
rect 213913 153310 217242 153312
rect 228968 153368 232011 153370
rect 228968 153312 231950 153368
rect 232006 153312 232011 153368
rect 228968 153310 232011 153312
rect 213913 153307 213979 153310
rect 231945 153307 232011 153310
rect 232446 153172 232452 153236
rect 232516 153234 232522 153236
rect 241421 153234 241487 153237
rect 232516 153232 241487 153234
rect 232516 153176 241426 153232
rect 241482 153176 241487 153232
rect 232516 153174 241487 153176
rect 232516 153172 232522 153174
rect 241421 153171 241487 153174
rect 265893 153234 265959 153237
rect 265893 153232 267842 153234
rect 265893 153176 265898 153232
rect 265954 153176 267842 153232
rect 265893 153174 267842 153176
rect 265893 153171 265959 153174
rect 267782 153098 267842 153174
rect 268334 153098 268394 153340
rect 282821 153234 282887 153237
rect 279956 153232 282887 153234
rect 279956 153176 282826 153232
rect 282882 153176 282887 153232
rect 279956 153174 282887 153176
rect 282821 153171 282887 153174
rect 214005 152690 214071 152693
rect 217182 152690 217242 153068
rect 267782 153038 268394 153098
rect 231761 152962 231827 152965
rect 228968 152960 231827 152962
rect 228968 152904 231766 152960
rect 231822 152904 231827 152960
rect 228968 152902 231827 152904
rect 231761 152899 231827 152902
rect 214005 152688 217242 152690
rect 214005 152632 214010 152688
rect 214066 152632 217242 152688
rect 214005 152630 217242 152632
rect 265709 152690 265775 152693
rect 268150 152690 268210 152932
rect 265709 152688 268210 152690
rect 265709 152632 265714 152688
rect 265770 152632 268210 152688
rect 265709 152630 268210 152632
rect 579797 152690 579863 152693
rect 583520 152690 584960 152780
rect 579797 152688 584960 152690
rect 579797 152632 579802 152688
rect 579858 152632 584960 152688
rect 579797 152630 584960 152632
rect 214005 152627 214071 152630
rect 265709 152627 265775 152630
rect 579797 152627 579863 152630
rect 231669 152554 231735 152557
rect 228968 152552 231735 152554
rect 213913 152010 213979 152013
rect 217182 152010 217242 152524
rect 228968 152496 231674 152552
rect 231730 152496 231735 152552
rect 583520 152540 584960 152630
rect 228968 152494 231735 152496
rect 231669 152491 231735 152494
rect 264421 152146 264487 152149
rect 268150 152146 268210 152524
rect 282729 152418 282795 152421
rect 279956 152416 282795 152418
rect 279956 152360 282734 152416
rect 282790 152360 282795 152416
rect 279956 152358 282795 152360
rect 282729 152355 282795 152358
rect 264421 152144 268210 152146
rect 264421 152088 264426 152144
rect 264482 152088 268210 152144
rect 264421 152086 268210 152088
rect 264421 152083 264487 152086
rect 231577 152010 231643 152013
rect 213913 152008 217242 152010
rect 213913 151952 213918 152008
rect 213974 151952 217242 152008
rect 213913 151950 217242 151952
rect 228968 152008 231643 152010
rect 228968 151952 231582 152008
rect 231638 151952 231643 152008
rect 228968 151950 231643 151952
rect 213913 151947 213979 151950
rect 231577 151947 231643 151950
rect 215017 151874 215083 151877
rect 265801 151874 265867 151877
rect 215017 151872 217058 151874
rect 215017 151816 215022 151872
rect 215078 151830 217058 151872
rect 265801 151872 267842 151874
rect 217182 151830 217242 151844
rect 215078 151816 217242 151830
rect 215017 151814 217242 151816
rect 215017 151811 215083 151814
rect 216998 151770 217242 151814
rect 265801 151816 265806 151872
rect 265862 151816 267842 151872
rect 265801 151814 267842 151816
rect 265801 151811 265867 151814
rect 267782 151738 267842 151814
rect 268334 151738 268394 151980
rect 280245 151738 280311 151741
rect 267782 151678 268394 151738
rect 279956 151736 280311 151738
rect 279956 151680 280250 151736
rect 280306 151680 280311 151736
rect 279956 151678 280311 151680
rect 280245 151675 280311 151678
rect 231669 151602 231735 151605
rect 228968 151600 231735 151602
rect 228968 151544 231674 151600
rect 231730 151544 231735 151600
rect 228968 151542 231735 151544
rect 231669 151539 231735 151542
rect 265985 151330 266051 151333
rect 268150 151330 268210 151572
rect 265985 151328 268210 151330
rect 265985 151272 265990 151328
rect 266046 151272 268210 151328
rect 265985 151270 268210 151272
rect 265985 151267 266051 151270
rect 214005 150786 214071 150789
rect 217182 150786 217242 151164
rect 231761 151058 231827 151061
rect 228968 151056 231827 151058
rect 228968 151000 231766 151056
rect 231822 151000 231827 151056
rect 228968 150998 231827 151000
rect 231761 150995 231827 150998
rect 233785 151058 233851 151061
rect 252502 151058 252508 151060
rect 233785 151056 252508 151058
rect 233785 151000 233790 151056
rect 233846 151000 252508 151056
rect 233785 150998 252508 151000
rect 233785 150995 233851 150998
rect 252502 150996 252508 150998
rect 252572 150996 252578 151060
rect 265893 150922 265959 150925
rect 268150 150922 268210 151164
rect 282821 150922 282887 150925
rect 265893 150920 268210 150922
rect 265893 150864 265898 150920
rect 265954 150864 268210 150920
rect 265893 150862 268210 150864
rect 279956 150920 282887 150922
rect 279956 150864 282826 150920
rect 282882 150864 282887 150920
rect 279956 150862 282887 150864
rect 265893 150859 265959 150862
rect 282821 150859 282887 150862
rect 214005 150784 217242 150786
rect 214005 150728 214010 150784
rect 214066 150728 217242 150784
rect 214005 150726 217242 150728
rect 214005 150723 214071 150726
rect 213913 150650 213979 150653
rect 231761 150650 231827 150653
rect 213913 150648 217242 150650
rect 213913 150592 213918 150648
rect 213974 150592 217242 150648
rect 213913 150590 217242 150592
rect 228968 150648 231827 150650
rect 228968 150592 231766 150648
rect 231822 150592 231827 150648
rect 228968 150590 231827 150592
rect 213913 150587 213979 150590
rect 217182 150484 217242 150590
rect 231761 150587 231827 150590
rect 265801 150514 265867 150517
rect 268150 150514 268210 150756
rect 265801 150512 268210 150514
rect 265801 150456 265806 150512
rect 265862 150456 268210 150512
rect 265801 150454 268210 150456
rect 265801 150451 265867 150454
rect 214557 150242 214623 150245
rect 214557 150240 217242 150242
rect 214557 150184 214562 150240
rect 214618 150184 217242 150240
rect 214557 150182 217242 150184
rect 214557 150179 214623 150182
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect 217182 149804 217242 150182
rect 231761 150106 231827 150109
rect 228968 150104 231827 150106
rect 228968 150048 231766 150104
rect 231822 150048 231827 150104
rect 228968 150046 231827 150048
rect 231761 150043 231827 150046
rect 265341 150106 265407 150109
rect 268150 150106 268210 150348
rect 282821 150106 282887 150109
rect 265341 150104 268210 150106
rect 265341 150048 265346 150104
rect 265402 150048 268210 150104
rect 265341 150046 268210 150048
rect 279956 150104 282887 150106
rect 279956 150048 282826 150104
rect 282882 150048 282887 150104
rect 279956 150046 282887 150048
rect 265341 150043 265407 150046
rect 282821 150043 282887 150046
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 230933 149698 230999 149701
rect 228968 149696 230999 149698
rect 228968 149640 230938 149696
rect 230994 149640 230999 149696
rect 228968 149638 230999 149640
rect 230933 149635 230999 149638
rect 265893 149698 265959 149701
rect 268150 149698 268210 149940
rect 265893 149696 268210 149698
rect 265893 149640 265898 149696
rect 265954 149640 268210 149696
rect 265893 149638 268210 149640
rect 265893 149635 265959 149638
rect 213913 149562 213979 149565
rect 213913 149560 217242 149562
rect 213913 149504 213918 149560
rect 213974 149504 217242 149560
rect 213913 149502 217242 149504
rect 213913 149499 213979 149502
rect 217182 149124 217242 149502
rect 265801 149290 265867 149293
rect 268150 149290 268210 149532
rect 281533 149426 281599 149429
rect 279956 149424 281599 149426
rect 279956 149368 281538 149424
rect 281594 149368 281599 149424
rect 279956 149366 281599 149368
rect 281533 149363 281599 149366
rect 265801 149288 268210 149290
rect 265801 149232 265806 149288
rect 265862 149232 268210 149288
rect 265801 149230 268210 149232
rect 265801 149227 265867 149230
rect 231669 149154 231735 149157
rect 228968 149152 231735 149154
rect 228968 149096 231674 149152
rect 231730 149096 231735 149152
rect 228968 149094 231735 149096
rect 231669 149091 231735 149094
rect 214741 148882 214807 148885
rect 214741 148880 217242 148882
rect 214741 148824 214746 148880
rect 214802 148824 217242 148880
rect 214741 148822 217242 148824
rect 214741 148819 214807 148822
rect 217182 148444 217242 148822
rect 233366 148746 233372 148748
rect 228968 148686 233372 148746
rect 233366 148684 233372 148686
rect 233436 148684 233442 148748
rect 265433 148746 265499 148749
rect 268150 148746 268210 148988
rect 265433 148744 268210 148746
rect 265433 148688 265438 148744
rect 265494 148688 268210 148744
rect 265433 148686 268210 148688
rect 265433 148683 265499 148686
rect 282821 148610 282887 148613
rect 279956 148608 282887 148610
rect 265157 148338 265223 148341
rect 268150 148338 268210 148580
rect 279956 148552 282826 148608
rect 282882 148552 282887 148608
rect 279956 148550 282887 148552
rect 282821 148547 282887 148550
rect 265157 148336 268210 148338
rect 265157 148280 265162 148336
rect 265218 148280 268210 148336
rect 265157 148278 268210 148280
rect 265157 148275 265223 148278
rect 231761 148202 231827 148205
rect 228968 148200 231827 148202
rect 228968 148144 231766 148200
rect 231822 148144 231827 148200
rect 228968 148142 231827 148144
rect 231761 148139 231827 148142
rect 213913 148066 213979 148069
rect 213913 148064 217242 148066
rect 213913 148008 213918 148064
rect 213974 148008 217242 148064
rect 213913 148006 217242 148008
rect 213913 148003 213979 148006
rect 217182 147900 217242 148006
rect 265801 147930 265867 147933
rect 268518 147932 268578 148172
rect 265801 147928 268210 147930
rect 265801 147872 265806 147928
rect 265862 147872 268210 147928
rect 265801 147870 268210 147872
rect 265801 147867 265867 147870
rect 230473 147794 230539 147797
rect 228968 147792 230539 147794
rect 228968 147736 230478 147792
rect 230534 147736 230539 147792
rect 268150 147764 268210 147870
rect 268510 147868 268516 147932
rect 268580 147868 268586 147932
rect 282269 147794 282335 147797
rect 279956 147792 282335 147794
rect 228968 147734 230539 147736
rect 279956 147736 282274 147792
rect 282330 147736 282335 147792
rect 279956 147734 282335 147736
rect 230473 147731 230539 147734
rect 282269 147731 282335 147734
rect 231761 147250 231827 147253
rect 228968 147248 231827 147250
rect 213913 146706 213979 146709
rect 217182 146706 217242 147220
rect 228968 147192 231766 147248
rect 231822 147192 231827 147248
rect 228968 147190 231827 147192
rect 231761 147187 231827 147190
rect 265525 147114 265591 147117
rect 268150 147114 268210 147356
rect 281717 147114 281783 147117
rect 265525 147112 268210 147114
rect 265525 147056 265530 147112
rect 265586 147056 268210 147112
rect 265525 147054 268210 147056
rect 279956 147112 281783 147114
rect 279956 147056 281722 147112
rect 281778 147056 281783 147112
rect 279956 147054 281783 147056
rect 265525 147051 265591 147054
rect 281717 147051 281783 147054
rect 230933 146842 230999 146845
rect 228968 146840 230999 146842
rect 228968 146784 230938 146840
rect 230994 146784 230999 146840
rect 228968 146782 230999 146784
rect 230933 146779 230999 146782
rect 213913 146704 217242 146706
rect 213913 146648 213918 146704
rect 213974 146648 217242 146704
rect 213913 146646 217242 146648
rect 265801 146706 265867 146709
rect 268150 146706 268210 146948
rect 265801 146704 268210 146706
rect 265801 146648 265806 146704
rect 265862 146648 268210 146704
rect 265801 146646 268210 146648
rect 213913 146643 213979 146646
rect 265801 146643 265867 146646
rect 266077 146570 266143 146573
rect 266077 146568 268210 146570
rect 214557 146434 214623 146437
rect 214557 146432 216874 146434
rect 214557 146376 214562 146432
rect 214618 146376 216874 146432
rect 214557 146374 216874 146376
rect 214557 146371 214623 146374
rect 216814 146298 216874 146374
rect 217366 146298 217426 146540
rect 266077 146512 266082 146568
rect 266138 146512 268210 146568
rect 266077 146510 268210 146512
rect 266077 146507 266143 146510
rect 268150 146404 268210 146510
rect 231761 146298 231827 146301
rect 282821 146298 282887 146301
rect 216814 146238 217426 146298
rect 228968 146296 231827 146298
rect 228968 146240 231766 146296
rect 231822 146240 231827 146296
rect 228968 146238 231827 146240
rect 279956 146296 282887 146298
rect 279956 146240 282826 146296
rect 282882 146240 282887 146296
rect 279956 146238 282887 146240
rect 231761 146235 231827 146238
rect 282821 146235 282887 146238
rect 261569 146162 261635 146165
rect 268510 146162 268516 146164
rect 261569 146160 268516 146162
rect 261569 146104 261574 146160
rect 261630 146104 268516 146160
rect 261569 146102 268516 146104
rect 261569 146099 261635 146102
rect 268510 146100 268516 146102
rect 268580 146100 268586 146164
rect 231669 145890 231735 145893
rect 228968 145888 231735 145890
rect 213913 145346 213979 145349
rect 217182 145346 217242 145860
rect 228968 145832 231674 145888
rect 231730 145832 231735 145888
rect 228968 145830 231735 145832
rect 231669 145827 231735 145830
rect 264513 145754 264579 145757
rect 268150 145754 268210 145996
rect 264513 145752 268210 145754
rect 264513 145696 264518 145752
rect 264574 145696 268210 145752
rect 264513 145694 268210 145696
rect 264513 145691 264579 145694
rect 231761 145618 231827 145621
rect 249742 145618 249748 145620
rect 231761 145616 249748 145618
rect 231761 145560 231766 145616
rect 231822 145560 249748 145616
rect 231761 145558 249748 145560
rect 231761 145555 231827 145558
rect 249742 145556 249748 145558
rect 249812 145556 249818 145620
rect 231025 145346 231091 145349
rect 213913 145344 217242 145346
rect 213913 145288 213918 145344
rect 213974 145288 217242 145344
rect 213913 145286 217242 145288
rect 228968 145344 231091 145346
rect 228968 145288 231030 145344
rect 231086 145288 231091 145344
rect 228968 145286 231091 145288
rect 213913 145283 213979 145286
rect 231025 145283 231091 145286
rect 265801 145346 265867 145349
rect 268150 145346 268210 145588
rect 281993 145482 282059 145485
rect 279956 145480 282059 145482
rect 279956 145424 281998 145480
rect 282054 145424 282059 145480
rect 279956 145422 282059 145424
rect 281993 145419 282059 145422
rect 265801 145344 268210 145346
rect 265801 145288 265806 145344
rect 265862 145288 268210 145344
rect 265801 145286 268210 145288
rect 265801 145283 265867 145286
rect 173014 145012 173020 145076
rect 173084 145074 173090 145076
rect 173084 145014 200130 145074
rect 173084 145012 173090 145014
rect 200070 144938 200130 145014
rect 217366 144938 217426 145180
rect 241830 144938 241836 144940
rect 200070 144878 217426 144938
rect 228968 144878 241836 144938
rect 241830 144876 241836 144878
rect 241900 144876 241906 144940
rect 265525 144938 265591 144941
rect 268334 144938 268394 145180
rect 265525 144936 268394 144938
rect 265525 144880 265530 144936
rect 265586 144880 268394 144936
rect 265525 144878 268394 144880
rect 265525 144875 265591 144878
rect 282545 144802 282611 144805
rect 279956 144800 282611 144802
rect 265433 144530 265499 144533
rect 268150 144530 268210 144772
rect 279956 144744 282550 144800
rect 282606 144744 282611 144800
rect 279956 144742 282611 144744
rect 282545 144739 282611 144742
rect 265433 144528 268210 144530
rect 214005 143986 214071 143989
rect 217182 143986 217242 144500
rect 265433 144472 265438 144528
rect 265494 144472 268210 144528
rect 265433 144470 268210 144472
rect 265433 144467 265499 144470
rect 231761 144394 231827 144397
rect 228968 144392 231827 144394
rect 228968 144336 231766 144392
rect 231822 144336 231827 144392
rect 228968 144334 231827 144336
rect 231761 144331 231827 144334
rect 230974 144060 230980 144124
rect 231044 144122 231050 144124
rect 261477 144122 261543 144125
rect 231044 144120 261543 144122
rect 231044 144064 261482 144120
rect 261538 144064 261543 144120
rect 231044 144062 261543 144064
rect 231044 144060 231050 144062
rect 261477 144059 261543 144062
rect 231577 143986 231643 143989
rect 214005 143984 217242 143986
rect 214005 143928 214010 143984
rect 214066 143928 217242 143984
rect 214005 143926 217242 143928
rect 228968 143984 231643 143986
rect 228968 143928 231582 143984
rect 231638 143928 231643 143984
rect 228968 143926 231643 143928
rect 214005 143923 214071 143926
rect 231577 143923 231643 143926
rect 265801 143986 265867 143989
rect 268150 143986 268210 144364
rect 282821 143986 282887 143989
rect 265801 143984 268210 143986
rect 265801 143928 265806 143984
rect 265862 143928 268210 143984
rect 265801 143926 268210 143928
rect 279956 143984 282887 143986
rect 279956 143928 282826 143984
rect 282882 143928 282887 143984
rect 279956 143926 282887 143928
rect 265801 143923 265867 143926
rect 282821 143923 282887 143926
rect 213913 143578 213979 143581
rect 217366 143578 217426 143820
rect 213913 143576 217426 143578
rect 213913 143520 213918 143576
rect 213974 143520 217426 143576
rect 213913 143518 217426 143520
rect 265893 143578 265959 143581
rect 268150 143578 268210 143820
rect 265893 143576 268210 143578
rect 265893 143520 265898 143576
rect 265954 143520 268210 143576
rect 265893 143518 268210 143520
rect 213913 143515 213979 143518
rect 265893 143515 265959 143518
rect 231761 143442 231827 143445
rect 228968 143440 231827 143442
rect 228968 143384 231766 143440
rect 231822 143384 231827 143440
rect 228968 143382 231827 143384
rect 231761 143379 231827 143382
rect 213913 142762 213979 142765
rect 217182 142762 217242 143276
rect 265709 143170 265775 143173
rect 268150 143170 268210 143412
rect 285622 143170 285628 143172
rect 265709 143168 268210 143170
rect 265709 143112 265714 143168
rect 265770 143112 268210 143168
rect 265709 143110 268210 143112
rect 279956 143110 285628 143170
rect 265709 143107 265775 143110
rect 285622 143108 285628 143110
rect 285692 143108 285698 143172
rect 231669 143034 231735 143037
rect 228968 143032 231735 143034
rect 228968 142976 231674 143032
rect 231730 142976 231735 143032
rect 228968 142974 231735 142976
rect 231669 142971 231735 142974
rect 213913 142760 217242 142762
rect 213913 142704 213918 142760
rect 213974 142704 217242 142760
rect 213913 142702 217242 142704
rect 265341 142762 265407 142765
rect 268150 142762 268210 143004
rect 265341 142760 268210 142762
rect 265341 142704 265346 142760
rect 265402 142704 268210 142760
rect 265341 142702 268210 142704
rect 213913 142699 213979 142702
rect 265341 142699 265407 142702
rect 173198 142156 173204 142220
rect 173268 142218 173274 142220
rect 217182 142218 217242 142596
rect 231117 142490 231183 142493
rect 228968 142488 231183 142490
rect 228968 142432 231122 142488
rect 231178 142432 231183 142488
rect 228968 142430 231183 142432
rect 231117 142427 231183 142430
rect 264605 142354 264671 142357
rect 268518 142356 268578 142596
rect 281625 142490 281691 142493
rect 279956 142488 281691 142490
rect 279956 142432 281630 142488
rect 281686 142432 281691 142488
rect 279956 142430 281691 142432
rect 281625 142427 281691 142430
rect 264605 142352 268210 142354
rect 264605 142296 264610 142352
rect 264666 142296 268210 142352
rect 264605 142294 268210 142296
rect 264605 142291 264671 142294
rect 173268 142158 217242 142218
rect 268150 142188 268210 142294
rect 268510 142292 268516 142356
rect 268580 142292 268586 142356
rect 173268 142156 173274 142158
rect 258390 142082 258396 142084
rect 228968 142022 258396 142082
rect 258390 142020 258396 142022
rect 258460 142020 258466 142084
rect 264329 141946 264395 141949
rect 268510 141946 268516 141948
rect 264329 141944 268516 141946
rect 214005 141402 214071 141405
rect 217182 141402 217242 141916
rect 264329 141888 264334 141944
rect 264390 141888 268516 141944
rect 264329 141886 268516 141888
rect 264329 141883 264395 141886
rect 268510 141884 268516 141886
rect 268580 141884 268586 141948
rect 237598 141674 237604 141676
rect 228968 141614 237604 141674
rect 237598 141612 237604 141614
rect 237668 141612 237674 141676
rect 214005 141400 217242 141402
rect 214005 141344 214010 141400
rect 214066 141344 217242 141400
rect 214005 141342 217242 141344
rect 265985 141402 266051 141405
rect 268518 141402 268578 141780
rect 282821 141674 282887 141677
rect 279956 141672 282887 141674
rect 279956 141616 282826 141672
rect 282882 141616 282887 141672
rect 279956 141614 282887 141616
rect 282821 141611 282887 141614
rect 265985 141400 268578 141402
rect 265985 141344 265990 141400
rect 266046 141344 268578 141400
rect 265985 141342 268578 141344
rect 214005 141339 214071 141342
rect 265985 141339 266051 141342
rect 213913 140994 213979 140997
rect 217182 140994 217242 141236
rect 231761 141130 231827 141133
rect 228968 141128 231827 141130
rect 228968 141072 231766 141128
rect 231822 141072 231827 141128
rect 228968 141070 231827 141072
rect 231761 141067 231827 141070
rect 233734 141068 233740 141132
rect 233804 141130 233810 141132
rect 267774 141130 267780 141132
rect 233804 141070 267780 141130
rect 233804 141068 233810 141070
rect 267774 141068 267780 141070
rect 267844 141068 267850 141132
rect 213913 140992 217242 140994
rect 213913 140936 213918 140992
rect 213974 140936 217242 140992
rect 213913 140934 217242 140936
rect 265801 140994 265867 140997
rect 265801 140992 268210 140994
rect 265801 140936 265806 140992
rect 265862 140936 268210 140992
rect 265801 140934 268210 140936
rect 213913 140931 213979 140934
rect 265801 140931 265867 140934
rect 268150 140828 268210 140934
rect 268326 140932 268332 140996
rect 268396 140994 268402 140996
rect 268518 140994 268578 141236
rect 268396 140934 268578 140994
rect 268396 140932 268402 140934
rect 291326 140858 291332 140860
rect 279956 140798 291332 140858
rect 291326 140796 291332 140798
rect 291396 140796 291402 140860
rect 231761 140722 231827 140725
rect 228968 140720 231827 140722
rect 228968 140664 231766 140720
rect 231822 140664 231827 140720
rect 228968 140662 231827 140664
rect 231761 140659 231827 140662
rect 217182 140042 217242 140556
rect 231669 140178 231735 140181
rect 228968 140176 231735 140178
rect 228968 140120 231674 140176
rect 231730 140120 231735 140176
rect 228968 140118 231735 140120
rect 231669 140115 231735 140118
rect 260465 140178 260531 140181
rect 268150 140178 268210 140420
rect 281901 140178 281967 140181
rect 260465 140176 268210 140178
rect 260465 140120 260470 140176
rect 260526 140120 268210 140176
rect 260465 140118 268210 140120
rect 279956 140176 281967 140178
rect 279956 140120 281906 140176
rect 281962 140120 281967 140176
rect 279956 140118 281967 140120
rect 260465 140115 260531 140118
rect 281901 140115 281967 140118
rect 200070 139982 217242 140042
rect 168230 139436 168236 139500
rect 168300 139498 168306 139500
rect 200070 139498 200130 139982
rect 168300 139438 200130 139498
rect 213913 139498 213979 139501
rect 217182 139498 217242 139876
rect 236494 139844 236500 139908
rect 236564 139906 236570 139908
rect 236564 139846 263610 139906
rect 236564 139844 236570 139846
rect 244774 139770 244780 139772
rect 228968 139710 244780 139770
rect 244774 139708 244780 139710
rect 244844 139708 244850 139772
rect 251766 139708 251772 139772
rect 251836 139770 251842 139772
rect 260465 139770 260531 139773
rect 251836 139768 260531 139770
rect 251836 139712 260470 139768
rect 260526 139712 260531 139768
rect 251836 139710 260531 139712
rect 263550 139770 263610 139846
rect 268334 139770 268394 140012
rect 263550 139710 268394 139770
rect 251836 139708 251842 139710
rect 260465 139707 260531 139710
rect 213913 139496 217242 139498
rect 213913 139440 213918 139496
rect 213974 139440 217242 139496
rect 213913 139438 217242 139440
rect 265433 139498 265499 139501
rect 265433 139496 267842 139498
rect 265433 139440 265438 139496
rect 265494 139440 267842 139496
rect 265433 139438 267842 139440
rect 168300 139436 168306 139438
rect 213913 139435 213979 139438
rect 265433 139435 265499 139438
rect 267782 139362 267842 139438
rect 268334 139362 268394 139604
rect 282821 139362 282887 139365
rect 267782 139302 268394 139362
rect 279956 139360 282887 139362
rect 279956 139304 282826 139360
rect 282882 139304 282887 139360
rect 279956 139302 282887 139304
rect 282821 139299 282887 139302
rect 580257 139362 580323 139365
rect 583520 139362 584960 139452
rect 580257 139360 584960 139362
rect 580257 139304 580262 139360
rect 580318 139304 584960 139360
rect 580257 139302 584960 139304
rect 580257 139299 580323 139302
rect 232446 139226 232452 139228
rect 214005 138818 214071 138821
rect 217182 138818 217242 139196
rect 228968 139166 232452 139226
rect 232446 139164 232452 139166
rect 232516 139164 232522 139228
rect 583520 139212 584960 139302
rect 233182 138818 233188 138820
rect 214005 138816 217242 138818
rect 214005 138760 214010 138816
rect 214066 138760 217242 138816
rect 214005 138758 217242 138760
rect 228968 138758 233188 138818
rect 214005 138755 214071 138758
rect 233182 138756 233188 138758
rect 233252 138756 233258 138820
rect 265433 138818 265499 138821
rect 268150 138818 268210 139196
rect 265433 138816 268210 138818
rect 265433 138760 265438 138816
rect 265494 138760 268210 138816
rect 265433 138758 268210 138760
rect 265433 138755 265499 138758
rect 213913 138138 213979 138141
rect 217182 138138 217242 138652
rect 265157 138410 265223 138413
rect 268150 138410 268210 138652
rect 282729 138546 282795 138549
rect 279956 138544 282795 138546
rect 279956 138488 282734 138544
rect 282790 138488 282795 138544
rect 279956 138486 282795 138488
rect 282729 138483 282795 138486
rect 265157 138408 268210 138410
rect 265157 138352 265162 138408
rect 265218 138352 268210 138408
rect 265157 138350 268210 138352
rect 265157 138347 265223 138350
rect 241646 138274 241652 138276
rect 228968 138214 241652 138274
rect 241646 138212 241652 138214
rect 241716 138212 241722 138276
rect 213913 138136 217242 138138
rect 213913 138080 213918 138136
rect 213974 138080 217242 138136
rect 213913 138078 217242 138080
rect 265617 138138 265683 138141
rect 265617 138136 267842 138138
rect 265617 138080 265622 138136
rect 265678 138080 267842 138136
rect 265617 138078 267842 138080
rect 213913 138075 213979 138078
rect 265617 138075 265683 138078
rect 267782 138002 267842 138078
rect 268334 138002 268394 138244
rect 213913 137458 213979 137461
rect 217182 137458 217242 137972
rect 267782 137942 268394 138002
rect 238518 137866 238524 137868
rect 228968 137806 238524 137866
rect 238518 137804 238524 137806
rect 238588 137804 238594 137868
rect 282821 137866 282887 137869
rect 279956 137864 282887 137866
rect 265617 137594 265683 137597
rect 268150 137594 268210 137836
rect 279956 137808 282826 137864
rect 282882 137808 282887 137864
rect 279956 137806 282887 137808
rect 282821 137803 282887 137806
rect 265617 137592 268210 137594
rect 265617 137536 265622 137592
rect 265678 137536 268210 137592
rect 265617 137534 268210 137536
rect 265617 137531 265683 137534
rect 213913 137456 217242 137458
rect 213913 137400 213918 137456
rect 213974 137400 217242 137456
rect 213913 137398 217242 137400
rect 213913 137395 213979 137398
rect 231393 137322 231459 137325
rect 228968 137320 231459 137322
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 166206 136716 166212 136780
rect 166276 136778 166282 136780
rect 217182 136778 217242 137292
rect 228968 137264 231398 137320
rect 231454 137264 231459 137320
rect 228968 137262 231459 137264
rect 231393 137259 231459 137262
rect 232446 137124 232452 137188
rect 232516 137186 232522 137188
rect 268150 137186 268210 137428
rect 232516 137126 268210 137186
rect 232516 137124 232522 137126
rect 282177 137050 282243 137053
rect 279956 137048 282243 137050
rect 231761 136914 231827 136917
rect 228968 136912 231827 136914
rect 228968 136856 231766 136912
rect 231822 136856 231827 136912
rect 228968 136854 231827 136856
rect 231761 136851 231827 136854
rect 166276 136718 217242 136778
rect 265525 136778 265591 136781
rect 268150 136778 268210 137020
rect 279956 136992 282182 137048
rect 282238 136992 282243 137048
rect 279956 136990 282243 136992
rect 282177 136987 282243 136990
rect 265525 136776 268210 136778
rect 265525 136720 265530 136776
rect 265586 136720 268210 136776
rect 265525 136718 268210 136720
rect 166276 136716 166282 136718
rect 265525 136715 265591 136718
rect 213177 136098 213243 136101
rect 217182 136098 217242 136612
rect 240358 136370 240364 136372
rect 228968 136310 240364 136370
rect 240358 136308 240364 136310
rect 240428 136308 240434 136372
rect 265617 136370 265683 136373
rect 268150 136370 268210 136612
rect 280153 136370 280219 136373
rect 265617 136368 268210 136370
rect 265617 136312 265622 136368
rect 265678 136312 268210 136368
rect 265617 136310 268210 136312
rect 279956 136368 280219 136370
rect 279956 136312 280158 136368
rect 280214 136312 280219 136368
rect 279956 136310 280219 136312
rect 265617 136307 265683 136310
rect 280153 136307 280219 136310
rect 213177 136096 217242 136098
rect 213177 136040 213182 136096
rect 213238 136040 217242 136096
rect 213177 136038 217242 136040
rect 213177 136035 213243 136038
rect 231393 135962 231459 135965
rect 228968 135960 231459 135962
rect 214741 135554 214807 135557
rect 217182 135554 217242 135932
rect 228968 135904 231398 135960
rect 231454 135904 231459 135960
rect 228968 135902 231459 135904
rect 231393 135899 231459 135902
rect 265341 135962 265407 135965
rect 268150 135962 268210 136204
rect 265341 135960 268210 135962
rect 265341 135904 265346 135960
rect 265402 135904 268210 135960
rect 265341 135902 268210 135904
rect 265341 135899 265407 135902
rect 266077 135826 266143 135829
rect 266077 135824 268210 135826
rect 266077 135768 266082 135824
rect 266138 135768 268210 135824
rect 266077 135766 268210 135768
rect 266077 135763 266143 135766
rect 268150 135660 268210 135766
rect 214741 135552 217242 135554
rect 214741 135496 214746 135552
rect 214802 135496 217242 135552
rect 214741 135494 217242 135496
rect 214741 135491 214807 135494
rect 231761 135418 231827 135421
rect 200070 135358 217242 135418
rect 228968 135416 231827 135418
rect 228968 135360 231766 135416
rect 231822 135360 231827 135416
rect 228968 135358 231827 135360
rect 170254 135220 170260 135284
rect 170324 135282 170330 135284
rect 200070 135282 200130 135358
rect 170324 135222 200130 135282
rect 217182 135252 217242 135358
rect 231761 135355 231827 135358
rect 265893 135418 265959 135421
rect 265893 135416 268210 135418
rect 265893 135360 265898 135416
rect 265954 135360 268210 135416
rect 265893 135358 268210 135360
rect 265893 135355 265959 135358
rect 238017 135282 238083 135285
rect 231718 135280 238083 135282
rect 231718 135224 238022 135280
rect 238078 135224 238083 135280
rect 268150 135252 268210 135358
rect 279926 135282 279986 135524
rect 296478 135282 296484 135284
rect 231718 135222 238083 135224
rect 279926 135222 296484 135282
rect 170324 135220 170330 135222
rect 231718 135010 231778 135222
rect 238017 135219 238083 135222
rect 296478 135220 296484 135222
rect 296548 135220 296554 135284
rect 228968 134950 231778 135010
rect 265525 134602 265591 134605
rect 268150 134602 268210 134844
rect 265525 134600 268210 134602
rect 214649 134194 214715 134197
rect 217182 134194 217242 134572
rect 265525 134544 265530 134600
rect 265586 134544 268210 134600
rect 265525 134542 268210 134544
rect 265525 134539 265591 134542
rect 231485 134466 231551 134469
rect 228968 134464 231551 134466
rect 228968 134408 231490 134464
rect 231546 134408 231551 134464
rect 228968 134406 231551 134408
rect 231485 134403 231551 134406
rect 214649 134192 217242 134194
rect 214649 134136 214654 134192
rect 214710 134136 217242 134192
rect 214649 134134 217242 134136
rect 265893 134194 265959 134197
rect 268150 134194 268210 134436
rect 265893 134192 268210 134194
rect 265893 134136 265898 134192
rect 265954 134136 268210 134192
rect 265893 134134 268210 134136
rect 279926 134194 279986 134708
rect 290590 134194 290596 134196
rect 279926 134134 290596 134194
rect 214649 134131 214715 134134
rect 265893 134131 265959 134134
rect 290590 134132 290596 134134
rect 290660 134132 290666 134196
rect 213913 134058 213979 134061
rect 231025 134058 231091 134061
rect 282821 134058 282887 134061
rect 213913 134056 217242 134058
rect 213913 134000 213918 134056
rect 213974 134000 217242 134056
rect 213913 133998 217242 134000
rect 228968 134056 231091 134058
rect 228968 134000 231030 134056
rect 231086 134000 231091 134056
rect 279956 134056 282887 134058
rect 228968 133998 231091 134000
rect 213913 133995 213979 133998
rect 217182 133892 217242 133998
rect 231025 133995 231091 133998
rect 265893 133922 265959 133925
rect 265893 133920 267842 133922
rect 265893 133864 265898 133920
rect 265954 133864 267842 133920
rect 265893 133862 267842 133864
rect 265893 133859 265959 133862
rect 267782 133786 267842 133862
rect 268334 133786 268394 134028
rect 279956 134000 282826 134056
rect 282882 134000 282887 134056
rect 279956 133998 282887 134000
rect 282821 133995 282887 133998
rect 267782 133726 268394 133786
rect 231577 133514 231643 133517
rect 228968 133512 231643 133514
rect 228968 133456 231582 133512
rect 231638 133456 231643 133512
rect 228968 133454 231643 133456
rect 231577 133451 231643 133454
rect 214005 132834 214071 132837
rect 217182 132834 217242 133348
rect 258758 133180 258764 133244
rect 258828 133242 258834 133244
rect 268150 133242 268210 133620
rect 282821 133242 282887 133245
rect 258828 133182 268210 133242
rect 279956 133240 282887 133242
rect 279956 133184 282826 133240
rect 282882 133184 282887 133240
rect 279956 133182 282887 133184
rect 258828 133180 258834 133182
rect 282821 133179 282887 133182
rect 230933 133106 230999 133109
rect 228968 133104 230999 133106
rect 228968 133048 230938 133104
rect 230994 133048 230999 133104
rect 228968 133046 230999 133048
rect 230933 133043 230999 133046
rect 214005 132832 217242 132834
rect 214005 132776 214010 132832
rect 214066 132776 217242 132832
rect 214005 132774 217242 132776
rect 265617 132834 265683 132837
rect 268150 132834 268210 133076
rect 265617 132832 268210 132834
rect 265617 132776 265622 132832
rect 265678 132776 268210 132832
rect 265617 132774 268210 132776
rect 214005 132771 214071 132774
rect 265617 132771 265683 132774
rect 213913 132562 213979 132565
rect 213913 132560 216874 132562
rect 213913 132504 213918 132560
rect 213974 132510 216874 132560
rect 217366 132510 217426 132668
rect 231669 132562 231735 132565
rect 213974 132504 217426 132510
rect 213913 132502 217426 132504
rect 228968 132560 231735 132562
rect 228968 132504 231674 132560
rect 231730 132504 231735 132560
rect 228968 132502 231735 132504
rect 213913 132499 213979 132502
rect 216814 132450 217426 132502
rect 231669 132499 231735 132502
rect 265893 132562 265959 132565
rect 265893 132560 267842 132562
rect 265893 132504 265898 132560
rect 265954 132504 267842 132560
rect 265893 132502 267842 132504
rect 265893 132499 265959 132502
rect 267782 132426 267842 132502
rect 268334 132426 268394 132668
rect 282821 132426 282887 132429
rect 267782 132366 268394 132426
rect 279956 132424 282887 132426
rect 279956 132368 282826 132424
rect 282882 132368 282887 132424
rect 279956 132366 282887 132368
rect 282821 132363 282887 132366
rect 231761 132154 231827 132157
rect 228968 132152 231827 132154
rect 228968 132096 231766 132152
rect 231822 132096 231827 132152
rect 228968 132094 231827 132096
rect 231761 132091 231827 132094
rect 265893 132018 265959 132021
rect 268150 132018 268210 132260
rect 265893 132016 268210 132018
rect 214005 131474 214071 131477
rect 217182 131474 217242 131988
rect 265893 131960 265898 132016
rect 265954 131960 268210 132016
rect 265893 131958 268210 131960
rect 265893 131955 265959 131958
rect 231301 131610 231367 131613
rect 228968 131608 231367 131610
rect 228968 131552 231306 131608
rect 231362 131552 231367 131608
rect 228968 131550 231367 131552
rect 231301 131547 231367 131550
rect 265157 131610 265223 131613
rect 268150 131610 268210 131852
rect 265157 131608 268210 131610
rect 265157 131552 265162 131608
rect 265218 131552 268210 131608
rect 265157 131550 268210 131552
rect 265157 131547 265223 131550
rect 214005 131472 217242 131474
rect 214005 131416 214010 131472
rect 214066 131416 217242 131472
rect 214005 131414 217242 131416
rect 214005 131411 214071 131414
rect 213913 131202 213979 131205
rect 213913 131200 216874 131202
rect 213913 131144 213918 131200
rect 213974 131144 216874 131200
rect 213913 131142 216874 131144
rect 213913 131139 213979 131142
rect 216814 131066 216874 131142
rect 217366 131066 217426 131308
rect 231669 131202 231735 131205
rect 228968 131200 231735 131202
rect 228968 131144 231674 131200
rect 231730 131144 231735 131200
rect 228968 131142 231735 131144
rect 231669 131139 231735 131142
rect 265617 131202 265683 131205
rect 268334 131202 268394 131444
rect 265617 131200 268394 131202
rect 265617 131144 265622 131200
rect 265678 131144 268394 131200
rect 265617 131142 268394 131144
rect 279926 131202 279986 131716
rect 288566 131202 288572 131204
rect 279926 131142 288572 131202
rect 265617 131139 265683 131142
rect 288566 131140 288572 131142
rect 288636 131140 288642 131204
rect 216814 131006 217426 131066
rect 231761 130658 231827 130661
rect 228968 130656 231827 130658
rect 214005 130114 214071 130117
rect 217182 130114 217242 130628
rect 228968 130600 231766 130656
rect 231822 130600 231827 130656
rect 228968 130598 231827 130600
rect 231761 130595 231827 130598
rect 265525 130658 265591 130661
rect 268150 130658 268210 131036
rect 282821 130930 282887 130933
rect 279956 130928 282887 130930
rect 279956 130872 282826 130928
rect 282882 130872 282887 130928
rect 279956 130870 282887 130872
rect 282821 130867 282887 130870
rect 265525 130656 268210 130658
rect 265525 130600 265530 130656
rect 265586 130600 268210 130656
rect 265525 130598 268210 130600
rect 265525 130595 265591 130598
rect 231393 130250 231459 130253
rect 228968 130248 231459 130250
rect 228968 130192 231398 130248
rect 231454 130192 231459 130248
rect 228968 130190 231459 130192
rect 231393 130187 231459 130190
rect 250294 130188 250300 130252
rect 250364 130250 250370 130252
rect 268150 130250 268210 130492
rect 250364 130190 268210 130250
rect 250364 130188 250370 130190
rect 282269 130114 282335 130117
rect 214005 130112 217242 130114
rect 214005 130056 214010 130112
rect 214066 130056 217242 130112
rect 279956 130112 282335 130114
rect 214005 130054 217242 130056
rect 214005 130051 214071 130054
rect 213913 129842 213979 129845
rect 213913 129840 216874 129842
rect 213913 129784 213918 129840
rect 213974 129784 216874 129840
rect 213913 129782 216874 129784
rect 213913 129779 213979 129782
rect 216814 129706 216874 129782
rect 217366 129706 217426 129948
rect 231669 129842 231735 129845
rect 228968 129840 231735 129842
rect 228968 129784 231674 129840
rect 231730 129784 231735 129840
rect 228968 129782 231735 129784
rect 231669 129779 231735 129782
rect 260046 129780 260052 129844
rect 260116 129842 260122 129844
rect 268150 129842 268210 130084
rect 279956 130056 282274 130112
rect 282330 130056 282335 130112
rect 279956 130054 282335 130056
rect 282269 130051 282335 130054
rect 260116 129782 268210 129842
rect 260116 129780 260122 129782
rect 216814 129646 217426 129706
rect 265893 129434 265959 129437
rect 268150 129434 268210 129676
rect 265893 129432 268210 129434
rect 265893 129376 265898 129432
rect 265954 129376 268210 129432
rect 265893 129374 268210 129376
rect 265893 129371 265959 129374
rect 66069 129298 66135 129301
rect 68142 129298 68816 129304
rect 231301 129298 231367 129301
rect 66069 129296 68816 129298
rect 66069 129240 66074 129296
rect 66130 129244 68816 129296
rect 228968 129296 231367 129298
rect 66130 129240 68202 129244
rect 66069 129238 68202 129240
rect 66069 129235 66135 129238
rect 217182 128890 217242 129268
rect 228968 129240 231306 129296
rect 231362 129240 231367 129296
rect 228968 129238 231367 129240
rect 231301 129235 231367 129238
rect 265617 129026 265683 129029
rect 268150 129026 268210 129268
rect 265617 129024 268210 129026
rect 265617 128968 265622 129024
rect 265678 128968 268210 129024
rect 265617 128966 268210 128968
rect 265617 128963 265683 128966
rect 231485 128890 231551 128893
rect 200070 128830 217242 128890
rect 228968 128888 231551 128890
rect 228968 128832 231490 128888
rect 231546 128832 231551 128888
rect 228968 128830 231551 128832
rect 168966 128420 168972 128484
rect 169036 128482 169042 128484
rect 200070 128482 200130 128830
rect 231485 128827 231551 128830
rect 169036 128422 200130 128482
rect 213913 128482 213979 128485
rect 217182 128482 217242 128724
rect 268518 128620 268578 128860
rect 279926 128754 279986 129404
rect 287278 128754 287284 128756
rect 279926 128694 287284 128754
rect 287278 128692 287284 128694
rect 287348 128692 287354 128756
rect 258030 128558 268210 128618
rect 213913 128480 217242 128482
rect 213913 128424 213918 128480
rect 213974 128424 217242 128480
rect 213913 128422 217242 128424
rect 169036 128420 169042 128422
rect 213913 128419 213979 128422
rect 255814 128420 255820 128484
rect 255884 128482 255890 128484
rect 258030 128482 258090 128558
rect 255884 128422 258090 128482
rect 268150 128452 268210 128558
rect 268510 128556 268516 128620
rect 268580 128556 268586 128620
rect 282821 128618 282887 128621
rect 279956 128616 282887 128618
rect 279956 128560 282826 128616
rect 282882 128560 282887 128616
rect 279956 128558 282887 128560
rect 282821 128555 282887 128558
rect 255884 128420 255890 128422
rect 231761 128346 231827 128349
rect 228968 128344 231827 128346
rect 228968 128288 231766 128344
rect 231822 128288 231827 128344
rect 228968 128286 231827 128288
rect 231761 128283 231827 128286
rect 262806 128148 262812 128212
rect 262876 128210 262882 128212
rect 268510 128210 268516 128212
rect 262876 128150 268516 128210
rect 262876 128148 262882 128150
rect 268510 128148 268516 128150
rect 268580 128148 268586 128212
rect 66161 128074 66227 128077
rect 68142 128074 68816 128080
rect 66161 128072 68816 128074
rect 66161 128016 66166 128072
rect 66222 128020 68816 128072
rect 66222 128016 68202 128020
rect 66161 128014 68202 128016
rect 66161 128011 66227 128014
rect 217182 127530 217242 128044
rect 231669 127938 231735 127941
rect 228968 127936 231735 127938
rect 228968 127880 231674 127936
rect 231730 127880 231735 127936
rect 228968 127878 231735 127880
rect 231669 127875 231735 127878
rect 265341 127666 265407 127669
rect 268150 127666 268210 127908
rect 281717 127802 281783 127805
rect 279956 127800 281783 127802
rect 279956 127744 281722 127800
rect 281778 127744 281783 127800
rect 279956 127742 281783 127744
rect 281717 127739 281783 127742
rect 265341 127664 268210 127666
rect 265341 127608 265346 127664
rect 265402 127608 268210 127664
rect 265341 127606 268210 127608
rect 265341 127603 265407 127606
rect 200070 127470 217242 127530
rect 169150 127060 169156 127124
rect 169220 127122 169226 127124
rect 200070 127122 200130 127470
rect 231669 127394 231735 127397
rect 228968 127392 231735 127394
rect 169220 127062 200130 127122
rect 213913 127122 213979 127125
rect 217182 127122 217242 127364
rect 228968 127336 231674 127392
rect 231730 127336 231735 127392
rect 228968 127334 231735 127336
rect 231669 127331 231735 127334
rect 265893 127258 265959 127261
rect 268518 127260 268578 127500
rect 265893 127256 268210 127258
rect 265893 127200 265898 127256
rect 265954 127200 268210 127256
rect 265893 127198 268210 127200
rect 265893 127195 265959 127198
rect 213913 127120 217242 127122
rect 213913 127064 213918 127120
rect 213974 127064 217242 127120
rect 268150 127092 268210 127198
rect 268510 127196 268516 127260
rect 268580 127196 268586 127260
rect 287094 127122 287100 127124
rect 213913 127062 217242 127064
rect 279956 127062 287100 127122
rect 169220 127060 169226 127062
rect 213913 127059 213979 127062
rect 287094 127060 287100 127062
rect 287164 127060 287170 127124
rect 231761 126986 231827 126989
rect 228968 126984 231827 126986
rect 228968 126928 231766 126984
rect 231822 126928 231827 126984
rect 228968 126926 231827 126928
rect 231761 126923 231827 126926
rect 264094 126788 264100 126852
rect 264164 126850 264170 126852
rect 268510 126850 268516 126852
rect 264164 126790 268516 126850
rect 264164 126788 264170 126790
rect 268510 126788 268516 126790
rect 268580 126788 268586 126852
rect 65149 126306 65215 126309
rect 68142 126306 68816 126312
rect 65149 126304 68816 126306
rect 65149 126248 65154 126304
rect 65210 126252 68816 126304
rect 65210 126248 68202 126252
rect 65149 126246 68202 126248
rect 65149 126243 65215 126246
rect 214005 126170 214071 126173
rect 217182 126170 217242 126684
rect 231117 126442 231183 126445
rect 228968 126440 231183 126442
rect 228968 126384 231122 126440
rect 231178 126384 231183 126440
rect 228968 126382 231183 126384
rect 231117 126379 231183 126382
rect 265893 126442 265959 126445
rect 268150 126442 268210 126684
rect 265893 126440 268210 126442
rect 265893 126384 265898 126440
rect 265954 126384 268210 126440
rect 265893 126382 268210 126384
rect 265893 126379 265959 126382
rect 282821 126306 282887 126309
rect 279956 126304 282887 126306
rect 214005 126168 217242 126170
rect 214005 126112 214010 126168
rect 214066 126112 217242 126168
rect 214005 126110 217242 126112
rect 214005 126107 214071 126110
rect 231025 126034 231091 126037
rect 228968 126032 231091 126034
rect 213913 125762 213979 125765
rect 217182 125762 217242 126004
rect 228968 125976 231030 126032
rect 231086 125976 231091 126032
rect 228968 125974 231091 125976
rect 231025 125971 231091 125974
rect 265249 126034 265315 126037
rect 268150 126034 268210 126276
rect 279956 126248 282826 126304
rect 282882 126248 282887 126304
rect 279956 126246 282887 126248
rect 282821 126243 282887 126246
rect 265249 126032 268210 126034
rect 265249 125976 265254 126032
rect 265310 125976 268210 126032
rect 265249 125974 268210 125976
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 265249 125971 265315 125974
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 213913 125760 217242 125762
rect 213913 125704 213918 125760
rect 213974 125704 217242 125760
rect 213913 125702 217242 125704
rect 213913 125699 213979 125702
rect 266169 125626 266235 125629
rect 268150 125626 268210 125868
rect 266169 125624 268210 125626
rect 266169 125568 266174 125624
rect 266230 125568 268210 125624
rect 266169 125566 268210 125568
rect 266169 125563 266235 125566
rect 230974 125490 230980 125492
rect 228968 125430 230980 125490
rect 230974 125428 230980 125430
rect 231044 125428 231050 125492
rect 282821 125490 282887 125493
rect 279956 125488 282887 125490
rect 279956 125432 282826 125488
rect 282882 125432 282887 125488
rect 279956 125430 282887 125432
rect 282821 125427 282887 125430
rect 67633 125218 67699 125221
rect 68142 125218 68816 125224
rect 67633 125216 68816 125218
rect 67633 125160 67638 125216
rect 67694 125164 68816 125216
rect 67694 125160 68202 125164
rect 67633 125158 68202 125160
rect 67633 125155 67699 125158
rect 214005 124810 214071 124813
rect 217182 124810 217242 125324
rect 231761 125082 231827 125085
rect 228968 125080 231827 125082
rect 228968 125024 231766 125080
rect 231822 125024 231827 125080
rect 228968 125022 231827 125024
rect 231761 125019 231827 125022
rect 265893 125082 265959 125085
rect 268150 125082 268210 125324
rect 265893 125080 268210 125082
rect 265893 125024 265898 125080
rect 265954 125024 268210 125080
rect 265893 125022 268210 125024
rect 265893 125019 265959 125022
rect 214005 124808 217242 124810
rect 214005 124752 214010 124808
rect 214066 124752 217242 124808
rect 214005 124750 217242 124752
rect 214005 124747 214071 124750
rect 265525 124674 265591 124677
rect 268150 124674 268210 124916
rect 282085 124810 282151 124813
rect 279956 124808 282151 124810
rect 279956 124752 282090 124808
rect 282146 124752 282151 124808
rect 279956 124750 282151 124752
rect 282085 124747 282151 124750
rect 265525 124672 268210 124674
rect 213913 124402 213979 124405
rect 217182 124402 217242 124644
rect 265525 124616 265530 124672
rect 265586 124616 268210 124672
rect 265525 124614 268210 124616
rect 265525 124611 265591 124614
rect 231301 124538 231367 124541
rect 228968 124536 231367 124538
rect 228968 124480 231306 124536
rect 231362 124480 231367 124536
rect 228968 124478 231367 124480
rect 231301 124475 231367 124478
rect 213913 124400 217242 124402
rect 213913 124344 213918 124400
rect 213974 124344 217242 124400
rect 213913 124342 217242 124344
rect 213913 124339 213979 124342
rect 265985 124266 266051 124269
rect 268334 124266 268394 124508
rect 265985 124264 268394 124266
rect 265985 124208 265990 124264
rect 266046 124208 268394 124264
rect 265985 124206 268394 124208
rect 265985 124203 266051 124206
rect 231577 124130 231643 124133
rect 228968 124128 231643 124130
rect -960 123572 480 123812
rect 65977 123586 66043 123589
rect 68142 123586 68816 123592
rect 65977 123584 68816 123586
rect 65977 123528 65982 123584
rect 66038 123532 68816 123584
rect 214005 123586 214071 123589
rect 217182 123586 217242 124100
rect 228968 124072 231582 124128
rect 231638 124072 231643 124128
rect 228968 124070 231643 124072
rect 231577 124067 231643 124070
rect 264329 123858 264395 123861
rect 268150 123858 268210 124100
rect 282821 123994 282887 123997
rect 279956 123992 282887 123994
rect 279956 123936 282826 123992
rect 282882 123936 282887 123992
rect 279956 123934 282887 123936
rect 282821 123931 282887 123934
rect 264329 123856 268210 123858
rect 264329 123800 264334 123856
rect 264390 123800 268210 123856
rect 264329 123798 268210 123800
rect 264329 123795 264395 123798
rect 231577 123586 231643 123589
rect 214005 123584 217242 123586
rect 66038 123528 68202 123532
rect 65977 123526 68202 123528
rect 214005 123528 214010 123584
rect 214066 123528 217242 123584
rect 214005 123526 217242 123528
rect 228968 123584 231643 123586
rect 228968 123528 231582 123584
rect 231638 123528 231643 123584
rect 228968 123526 231643 123528
rect 65977 123523 66043 123526
rect 214005 123523 214071 123526
rect 231577 123523 231643 123526
rect 265525 123450 265591 123453
rect 268150 123450 268210 123692
rect 265525 123448 268210 123450
rect 213913 123178 213979 123181
rect 217182 123178 217242 123420
rect 265525 123392 265530 123448
rect 265586 123392 268210 123448
rect 265525 123390 268210 123392
rect 265525 123387 265591 123390
rect 231761 123178 231827 123181
rect 213913 123176 217242 123178
rect 213913 123120 213918 123176
rect 213974 123120 217242 123176
rect 213913 123118 217242 123120
rect 228968 123176 231827 123178
rect 228968 123120 231766 123176
rect 231822 123120 231827 123176
rect 228968 123118 231827 123120
rect 213913 123115 213979 123118
rect 231761 123115 231827 123118
rect 265065 123042 265131 123045
rect 268150 123042 268210 123284
rect 282729 123178 282795 123181
rect 279956 123176 282795 123178
rect 279956 123120 282734 123176
rect 282790 123120 282795 123176
rect 279956 123118 282795 123120
rect 282729 123115 282795 123118
rect 265065 123040 268210 123042
rect 265065 122984 265070 123040
rect 265126 122984 268210 123040
rect 265065 122982 268210 122984
rect 265065 122979 265131 122982
rect 266261 122906 266327 122909
rect 266261 122904 267842 122906
rect 266261 122848 266266 122904
rect 266322 122848 267842 122904
rect 266261 122846 267842 122848
rect 266261 122843 266327 122846
rect 67541 122634 67607 122637
rect 68142 122634 68816 122640
rect 67541 122632 68816 122634
rect 67541 122576 67546 122632
rect 67602 122580 68816 122632
rect 67602 122576 68202 122580
rect 67541 122574 68202 122576
rect 67541 122571 67607 122574
rect 213913 122226 213979 122229
rect 217182 122226 217242 122740
rect 231485 122634 231551 122637
rect 228968 122632 231551 122634
rect 228968 122576 231490 122632
rect 231546 122576 231551 122632
rect 228968 122574 231551 122576
rect 267782 122634 267842 122846
rect 268334 122634 268394 122876
rect 267782 122574 268394 122634
rect 231485 122571 231551 122574
rect 282085 122498 282151 122501
rect 279956 122496 282151 122498
rect 279956 122440 282090 122496
rect 282146 122440 282151 122496
rect 279956 122438 282151 122440
rect 282085 122435 282151 122438
rect 231301 122226 231367 122229
rect 213913 122224 217242 122226
rect 213913 122168 213918 122224
rect 213974 122168 217242 122224
rect 213913 122166 217242 122168
rect 228968 122224 231367 122226
rect 228968 122168 231306 122224
rect 231362 122168 231367 122224
rect 228968 122166 231367 122168
rect 213913 122163 213979 122166
rect 231301 122163 231367 122166
rect 265985 122090 266051 122093
rect 268150 122090 268210 122332
rect 265985 122088 268210 122090
rect 214465 121682 214531 121685
rect 217182 121682 217242 122060
rect 265985 122032 265990 122088
rect 266046 122032 268210 122088
rect 265985 122030 268210 122032
rect 265985 122027 266051 122030
rect 230841 121682 230907 121685
rect 214465 121680 217242 121682
rect 214465 121624 214470 121680
rect 214526 121624 217242 121680
rect 214465 121622 217242 121624
rect 228968 121680 230907 121682
rect 228968 121624 230846 121680
rect 230902 121624 230907 121680
rect 228968 121622 230907 121624
rect 214465 121619 214531 121622
rect 230841 121619 230907 121622
rect 265893 121682 265959 121685
rect 268518 121684 268578 121924
rect 265893 121680 268210 121682
rect 265893 121624 265898 121680
rect 265954 121624 268210 121680
rect 265893 121622 268210 121624
rect 265893 121619 265959 121622
rect 268150 121516 268210 121622
rect 268510 121620 268516 121684
rect 268580 121620 268586 121684
rect 279956 121622 287070 121682
rect 287010 121546 287070 121622
rect 294270 121546 294276 121548
rect 287010 121486 294276 121546
rect 294270 121484 294276 121486
rect 294340 121484 294346 121548
rect 67449 120866 67515 120869
rect 68142 120866 68816 120872
rect 67449 120864 68816 120866
rect 67449 120808 67454 120864
rect 67510 120812 68816 120864
rect 214005 120866 214071 120869
rect 217182 120866 217242 121380
rect 231761 121274 231827 121277
rect 228968 121272 231827 121274
rect 228968 121216 231766 121272
rect 231822 121216 231827 121272
rect 228968 121214 231827 121216
rect 231761 121211 231827 121214
rect 214005 120864 217242 120866
rect 67510 120808 68202 120812
rect 67449 120806 68202 120808
rect 214005 120808 214010 120864
rect 214066 120808 217242 120864
rect 214005 120806 217242 120808
rect 265985 120866 266051 120869
rect 268150 120866 268210 121108
rect 281717 120866 281783 120869
rect 265985 120864 268210 120866
rect 265985 120808 265990 120864
rect 266046 120808 268210 120864
rect 265985 120806 268210 120808
rect 279956 120864 281783 120866
rect 279956 120808 281722 120864
rect 281778 120808 281783 120864
rect 279956 120806 281783 120808
rect 67449 120803 67515 120806
rect 214005 120803 214071 120806
rect 265985 120803 266051 120806
rect 281717 120803 281783 120806
rect 230933 120730 230999 120733
rect 228968 120728 230999 120730
rect 213913 120458 213979 120461
rect 217182 120458 217242 120700
rect 228968 120672 230938 120728
rect 230994 120672 230999 120728
rect 228968 120670 230999 120672
rect 230933 120667 230999 120670
rect 213913 120456 217242 120458
rect 213913 120400 213918 120456
rect 213974 120400 217242 120456
rect 213913 120398 217242 120400
rect 213913 120395 213979 120398
rect 264278 120396 264284 120460
rect 264348 120458 264354 120460
rect 268150 120458 268210 120700
rect 264348 120398 268210 120458
rect 264348 120396 264354 120398
rect 231117 120322 231183 120325
rect 228968 120320 231183 120322
rect 228968 120264 231122 120320
rect 231178 120264 231183 120320
rect 228968 120262 231183 120264
rect 231117 120259 231183 120262
rect 265893 120186 265959 120189
rect 265893 120184 267842 120186
rect 265893 120128 265898 120184
rect 265954 120128 267842 120184
rect 265893 120126 267842 120128
rect 265893 120123 265959 120126
rect 267782 120050 267842 120126
rect 268334 120050 268394 120292
rect 282453 120186 282519 120189
rect 279956 120184 282519 120186
rect 279956 120128 282458 120184
rect 282514 120128 282519 120184
rect 279956 120126 282519 120128
rect 282453 120123 282519 120126
rect 214005 119642 214071 119645
rect 217182 119642 217242 120020
rect 267782 119990 268394 120050
rect 261661 119914 261727 119917
rect 268510 119914 268516 119916
rect 261661 119912 268516 119914
rect 261661 119856 261666 119912
rect 261722 119856 268516 119912
rect 261661 119854 268516 119856
rect 261661 119851 261727 119854
rect 268510 119852 268516 119854
rect 268580 119852 268586 119916
rect 230933 119778 230999 119781
rect 228968 119776 230999 119778
rect 228968 119720 230938 119776
rect 230994 119720 230999 119776
rect 228968 119718 230999 119720
rect 230933 119715 230999 119718
rect 214005 119640 217242 119642
rect 214005 119584 214010 119640
rect 214066 119584 217242 119640
rect 214005 119582 217242 119584
rect 214005 119579 214071 119582
rect 265709 119506 265775 119509
rect 268150 119506 268210 119748
rect 265709 119504 268210 119506
rect 213269 119098 213335 119101
rect 217182 119098 217242 119476
rect 265709 119448 265714 119504
rect 265770 119448 268210 119504
rect 265709 119446 268210 119448
rect 265709 119443 265775 119446
rect 231761 119370 231827 119373
rect 282085 119370 282151 119373
rect 228968 119368 231827 119370
rect 228968 119312 231766 119368
rect 231822 119312 231827 119368
rect 279956 119368 282151 119370
rect 228968 119310 231827 119312
rect 231761 119307 231827 119310
rect 213269 119096 217242 119098
rect 213269 119040 213274 119096
rect 213330 119040 217242 119096
rect 213269 119038 217242 119040
rect 265249 119098 265315 119101
rect 268150 119098 268210 119340
rect 279956 119312 282090 119368
rect 282146 119312 282151 119368
rect 279956 119310 282151 119312
rect 282085 119307 282151 119310
rect 265249 119096 268210 119098
rect 265249 119040 265254 119096
rect 265310 119040 268210 119096
rect 265249 119038 268210 119040
rect 213269 119035 213335 119038
rect 265249 119035 265315 119038
rect 213913 118962 213979 118965
rect 231485 118962 231551 118965
rect 213913 118960 217242 118962
rect 213913 118904 213918 118960
rect 213974 118904 217242 118960
rect 213913 118902 217242 118904
rect 228968 118960 231551 118962
rect 228968 118904 231490 118960
rect 231546 118904 231551 118960
rect 228968 118902 231551 118904
rect 213913 118899 213979 118902
rect 217182 118796 217242 118902
rect 231485 118899 231551 118902
rect 258574 118764 258580 118828
rect 258644 118826 258650 118828
rect 258644 118766 267842 118826
rect 258644 118764 258650 118766
rect 267782 118690 267842 118766
rect 268334 118690 268394 118932
rect 267782 118630 268394 118690
rect 282821 118554 282887 118557
rect 279956 118552 282887 118554
rect 230657 118418 230723 118421
rect 228968 118416 230723 118418
rect 228968 118360 230662 118416
rect 230718 118360 230723 118416
rect 228968 118358 230723 118360
rect 230657 118355 230723 118358
rect 265525 118282 265591 118285
rect 268150 118282 268210 118524
rect 279956 118496 282826 118552
rect 282882 118496 282887 118552
rect 279956 118494 282887 118496
rect 282821 118491 282887 118494
rect 265525 118280 268210 118282
rect 265525 118224 265530 118280
rect 265586 118224 268210 118280
rect 265525 118222 268210 118224
rect 265525 118219 265591 118222
rect 214005 117602 214071 117605
rect 217182 117602 217242 118116
rect 231761 118010 231827 118013
rect 228968 118008 231827 118010
rect 228968 117952 231766 118008
rect 231822 117952 231827 118008
rect 228968 117950 231827 117952
rect 231761 117947 231827 117950
rect 265157 117874 265223 117877
rect 268150 117874 268210 118116
rect 282729 117874 282795 117877
rect 265157 117872 268210 117874
rect 265157 117816 265162 117872
rect 265218 117816 268210 117872
rect 265157 117814 268210 117816
rect 279956 117872 282795 117874
rect 279956 117816 282734 117872
rect 282790 117816 282795 117872
rect 279956 117814 282795 117816
rect 265157 117811 265223 117814
rect 282729 117811 282795 117814
rect 214005 117600 217242 117602
rect 214005 117544 214010 117600
rect 214066 117544 217242 117600
rect 214005 117542 217242 117544
rect 214005 117539 214071 117542
rect 230933 117466 230999 117469
rect 228968 117464 230999 117466
rect 213913 117330 213979 117333
rect 213913 117328 216874 117330
rect 213913 117272 213918 117328
rect 213974 117272 216874 117328
rect 213913 117270 216874 117272
rect 213913 117267 213979 117270
rect 216814 117194 216874 117270
rect 217366 117194 217426 117436
rect 228968 117408 230938 117464
rect 230994 117408 230999 117464
rect 228968 117406 230999 117408
rect 230933 117403 230999 117406
rect 265709 117466 265775 117469
rect 268150 117466 268210 117708
rect 265709 117464 268210 117466
rect 265709 117408 265714 117464
rect 265770 117408 268210 117464
rect 265709 117406 268210 117408
rect 265709 117403 265775 117406
rect 216814 117134 217426 117194
rect 230657 117058 230723 117061
rect 228968 117056 230723 117058
rect 228968 117000 230662 117056
rect 230718 117000 230723 117056
rect 228968 116998 230723 117000
rect 230657 116995 230723 116998
rect 266169 116922 266235 116925
rect 268150 116922 268210 117164
rect 282821 117058 282887 117061
rect 279956 117056 282887 117058
rect 279956 117000 282826 117056
rect 282882 117000 282887 117056
rect 279956 116998 282887 117000
rect 282821 116995 282887 116998
rect 266169 116920 268210 116922
rect 266169 116864 266174 116920
rect 266230 116864 268210 116920
rect 266169 116862 268210 116864
rect 266169 116859 266235 116862
rect 213913 116242 213979 116245
rect 217182 116242 217242 116756
rect 230565 116514 230631 116517
rect 228968 116512 230631 116514
rect 228968 116456 230570 116512
rect 230626 116456 230631 116512
rect 228968 116454 230631 116456
rect 230565 116451 230631 116454
rect 266077 116514 266143 116517
rect 268150 116514 268210 116756
rect 266077 116512 268210 116514
rect 266077 116456 266082 116512
rect 266138 116456 268210 116512
rect 266077 116454 268210 116456
rect 266077 116451 266143 116454
rect 282729 116378 282795 116381
rect 279956 116376 282795 116378
rect 213913 116240 217242 116242
rect 213913 116184 213918 116240
rect 213974 116184 217242 116240
rect 213913 116182 217242 116184
rect 213913 116179 213979 116182
rect 230749 116106 230815 116109
rect 228968 116104 230815 116106
rect 213361 115970 213427 115973
rect 213361 115968 216874 115970
rect 213361 115912 213366 115968
rect 213422 115912 216874 115968
rect 213361 115910 216874 115912
rect 213361 115907 213427 115910
rect 216814 115834 216874 115910
rect 217366 115834 217426 116076
rect 228968 116048 230754 116104
rect 230810 116048 230815 116104
rect 228968 116046 230815 116048
rect 230749 116043 230815 116046
rect 260230 116044 260236 116108
rect 260300 116106 260306 116108
rect 260300 116046 268210 116106
rect 260300 116044 260306 116046
rect 264513 115970 264579 115973
rect 267774 115970 267780 115972
rect 264513 115968 267780 115970
rect 264513 115912 264518 115968
rect 264574 115912 267780 115968
rect 264513 115910 267780 115912
rect 264513 115907 264579 115910
rect 267774 115908 267780 115910
rect 267844 115908 267850 115972
rect 268150 115940 268210 116046
rect 268326 116044 268332 116108
rect 268396 116106 268402 116108
rect 268518 116106 268578 116348
rect 279956 116320 282734 116376
rect 282790 116320 282795 116376
rect 279956 116318 282795 116320
rect 282729 116315 282795 116318
rect 268396 116046 268578 116106
rect 268396 116044 268402 116046
rect 216814 115774 217426 115834
rect 231761 115562 231827 115565
rect 282085 115562 282151 115565
rect 228968 115560 231827 115562
rect 228968 115504 231766 115560
rect 231822 115504 231827 115560
rect 279956 115560 282151 115562
rect 228968 115502 231827 115504
rect 231761 115499 231827 115502
rect 214005 115018 214071 115021
rect 217182 115018 217242 115396
rect 268150 115290 268210 115532
rect 279956 115504 282090 115560
rect 282146 115504 282151 115560
rect 279956 115502 282151 115504
rect 282085 115499 282151 115502
rect 258030 115230 268210 115290
rect 231761 115154 231827 115157
rect 228968 115152 231827 115154
rect 228968 115096 231766 115152
rect 231822 115096 231827 115152
rect 228968 115094 231827 115096
rect 231761 115091 231827 115094
rect 214005 115016 217242 115018
rect 214005 114960 214010 115016
rect 214066 114960 217242 115016
rect 214005 114958 217242 114960
rect 214005 114955 214071 114958
rect 213913 114610 213979 114613
rect 217182 114610 217242 114852
rect 249006 114820 249012 114884
rect 249076 114882 249082 114884
rect 258030 114882 258090 115230
rect 249076 114822 258090 114882
rect 265249 114882 265315 114885
rect 268150 114882 268210 115124
rect 265249 114880 268210 114882
rect 265249 114824 265254 114880
rect 265310 114824 268210 114880
rect 265249 114822 268210 114824
rect 249076 114820 249082 114822
rect 265249 114819 265315 114822
rect 262990 114684 262996 114748
rect 263060 114746 263066 114748
rect 281717 114746 281783 114749
rect 263060 114686 268210 114746
rect 279956 114744 281783 114746
rect 279956 114688 281722 114744
rect 281778 114688 281783 114744
rect 279956 114686 281783 114688
rect 263060 114684 263066 114686
rect 231669 114610 231735 114613
rect 213913 114608 217242 114610
rect 213913 114552 213918 114608
rect 213974 114552 217242 114608
rect 213913 114550 217242 114552
rect 228968 114608 231735 114610
rect 228968 114552 231674 114608
rect 231730 114552 231735 114608
rect 268150 114580 268210 114686
rect 281717 114683 281783 114686
rect 228968 114550 231735 114552
rect 213913 114547 213979 114550
rect 231669 114547 231735 114550
rect 230657 114202 230723 114205
rect 228968 114200 230723 114202
rect 214005 113658 214071 113661
rect 217182 113658 217242 114172
rect 228968 114144 230662 114200
rect 230718 114144 230723 114200
rect 228968 114142 230723 114144
rect 230657 114139 230723 114142
rect 265709 113930 265775 113933
rect 268150 113930 268210 114172
rect 282821 114066 282887 114069
rect 279956 114064 282887 114066
rect 279956 114008 282826 114064
rect 282882 114008 282887 114064
rect 279956 114006 282887 114008
rect 282821 114003 282887 114006
rect 265709 113928 268210 113930
rect 265709 113872 265714 113928
rect 265770 113872 268210 113928
rect 265709 113870 268210 113872
rect 265709 113867 265775 113870
rect 231485 113658 231551 113661
rect 214005 113656 217242 113658
rect 214005 113600 214010 113656
rect 214066 113600 217242 113656
rect 214005 113598 217242 113600
rect 228968 113656 231551 113658
rect 228968 113600 231490 113656
rect 231546 113600 231551 113656
rect 228968 113598 231551 113600
rect 214005 113595 214071 113598
rect 231485 113595 231551 113598
rect 265249 113522 265315 113525
rect 268150 113522 268210 113764
rect 265249 113520 268210 113522
rect 213913 113250 213979 113253
rect 217366 113250 217426 113492
rect 265249 113464 265254 113520
rect 265310 113464 268210 113520
rect 265249 113462 268210 113464
rect 265249 113459 265315 113462
rect 230565 113250 230631 113253
rect 213913 113248 217426 113250
rect 213913 113192 213918 113248
rect 213974 113192 217426 113248
rect 213913 113190 217426 113192
rect 228968 113248 230631 113250
rect 228968 113192 230570 113248
rect 230626 113192 230631 113248
rect 228968 113190 230631 113192
rect 213913 113187 213979 113190
rect 230565 113187 230631 113190
rect 265433 113250 265499 113253
rect 265433 113248 267842 113250
rect 265433 113192 265438 113248
rect 265494 113192 267842 113248
rect 265433 113190 267842 113192
rect 265433 113187 265499 113190
rect 267782 113114 267842 113190
rect 268334 113114 268394 113356
rect 292614 113250 292620 113252
rect 279956 113190 292620 113250
rect 292614 113188 292620 113190
rect 292684 113188 292690 113252
rect 267782 113054 268394 113114
rect 214005 112298 214071 112301
rect 217182 112298 217242 112812
rect 230933 112706 230999 112709
rect 228968 112704 230999 112706
rect 228968 112648 230938 112704
rect 230994 112648 230999 112704
rect 228968 112646 230999 112648
rect 230933 112643 230999 112646
rect 265525 112706 265591 112709
rect 268150 112706 268210 112948
rect 582833 112842 582899 112845
rect 583520 112842 584960 112932
rect 582833 112840 584960 112842
rect 582833 112784 582838 112840
rect 582894 112784 584960 112840
rect 582833 112782 584960 112784
rect 582833 112779 582899 112782
rect 265525 112704 268210 112706
rect 265525 112648 265530 112704
rect 265586 112648 268210 112704
rect 583520 112692 584960 112782
rect 265525 112646 268210 112648
rect 265525 112643 265591 112646
rect 231669 112298 231735 112301
rect 214005 112296 217242 112298
rect 214005 112240 214010 112296
rect 214066 112240 217242 112296
rect 214005 112238 217242 112240
rect 228968 112296 231735 112298
rect 228968 112240 231674 112296
rect 231730 112240 231735 112296
rect 228968 112238 231735 112240
rect 214005 112235 214071 112238
rect 231669 112235 231735 112238
rect 265709 112298 265775 112301
rect 268150 112298 268210 112540
rect 282085 112434 282151 112437
rect 279956 112432 282151 112434
rect 279956 112376 282090 112432
rect 282146 112376 282151 112432
rect 279956 112374 282151 112376
rect 282085 112371 282151 112374
rect 265709 112296 268210 112298
rect 265709 112240 265714 112296
rect 265770 112240 268210 112296
rect 265709 112238 268210 112240
rect 265709 112235 265775 112238
rect 266077 112162 266143 112165
rect 266077 112160 268210 112162
rect 213913 111890 213979 111893
rect 217182 111890 217242 112132
rect 266077 112104 266082 112160
rect 266138 112104 268210 112160
rect 266077 112102 268210 112104
rect 266077 112099 266143 112102
rect 268150 111996 268210 112102
rect 213913 111888 217242 111890
rect 213913 111832 213918 111888
rect 213974 111832 217242 111888
rect 213913 111830 217242 111832
rect 213913 111827 213979 111830
rect 167913 111754 167979 111757
rect 231761 111754 231827 111757
rect 282821 111754 282887 111757
rect 164694 111752 167979 111754
rect 164694 111696 167918 111752
rect 167974 111696 167979 111752
rect 164694 111694 167979 111696
rect 228968 111752 231827 111754
rect 228968 111696 231766 111752
rect 231822 111696 231827 111752
rect 228968 111694 231827 111696
rect 279956 111752 282887 111754
rect 279956 111696 282826 111752
rect 282882 111696 282887 111752
rect 279956 111694 282887 111696
rect 167913 111691 167979 111694
rect 231761 111691 231827 111694
rect 282821 111691 282887 111694
rect 214005 110938 214071 110941
rect 217182 110938 217242 111452
rect 231669 111346 231735 111349
rect 228968 111344 231735 111346
rect 228968 111288 231674 111344
rect 231730 111288 231735 111344
rect 228968 111286 231735 111288
rect 231669 111283 231735 111286
rect 265525 111346 265591 111349
rect 268150 111346 268210 111588
rect 265525 111344 268210 111346
rect 265525 111288 265530 111344
rect 265586 111288 268210 111344
rect 265525 111286 268210 111288
rect 265525 111283 265591 111286
rect 214005 110936 217242 110938
rect 214005 110880 214010 110936
rect 214066 110880 217242 110936
rect 214005 110878 217242 110880
rect 265157 110938 265223 110941
rect 268150 110938 268210 111180
rect 280153 110938 280219 110941
rect 265157 110936 268210 110938
rect 265157 110880 265162 110936
rect 265218 110880 268210 110936
rect 265157 110878 268210 110880
rect 279956 110936 280219 110938
rect 279956 110880 280158 110936
rect 280214 110880 280219 110936
rect 279956 110878 280219 110880
rect 214005 110875 214071 110878
rect 265157 110875 265223 110878
rect 280153 110875 280219 110878
rect 231577 110802 231643 110805
rect 228968 110800 231643 110802
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 213913 110530 213979 110533
rect 217366 110530 217426 110772
rect 228968 110744 231582 110800
rect 231638 110744 231643 110800
rect 228968 110742 231643 110744
rect 231577 110739 231643 110742
rect 213913 110528 217426 110530
rect 213913 110472 213918 110528
rect 213974 110472 217426 110528
rect 213913 110470 217426 110472
rect 265709 110530 265775 110533
rect 268150 110530 268210 110772
rect 265709 110528 268210 110530
rect 265709 110472 265714 110528
rect 265770 110472 268210 110528
rect 265709 110470 268210 110472
rect 213913 110467 213979 110470
rect 265709 110467 265775 110470
rect 231761 110394 231827 110397
rect 228968 110392 231827 110394
rect 228968 110336 231766 110392
rect 231822 110336 231827 110392
rect 228968 110334 231827 110336
rect 231761 110331 231827 110334
rect 167453 110122 167519 110125
rect 164694 110120 167519 110122
rect 164694 110064 167458 110120
rect 167514 110064 167519 110120
rect 164694 110062 167519 110064
rect 167453 110059 167519 110062
rect 214005 109714 214071 109717
rect 217182 109714 217242 110228
rect 264513 110122 264579 110125
rect 268150 110122 268210 110364
rect 264513 110120 268210 110122
rect 264513 110064 264518 110120
rect 264574 110064 268210 110120
rect 264513 110062 268210 110064
rect 264513 110059 264579 110062
rect 231117 109850 231183 109853
rect 228968 109848 231183 109850
rect 228968 109792 231122 109848
rect 231178 109792 231183 109848
rect 228968 109790 231183 109792
rect 231117 109787 231183 109790
rect 214005 109712 217242 109714
rect 214005 109656 214010 109712
rect 214066 109656 217242 109712
rect 214005 109654 217242 109656
rect 265525 109714 265591 109717
rect 268150 109714 268210 109956
rect 265525 109712 268210 109714
rect 265525 109656 265530 109712
rect 265586 109656 268210 109712
rect 265525 109654 268210 109656
rect 214005 109651 214071 109654
rect 265525 109651 265591 109654
rect 279926 109578 279986 110092
rect 291142 109578 291148 109580
rect 213913 109170 213979 109173
rect 217182 109170 217242 109548
rect 231485 109442 231551 109445
rect 228968 109440 231551 109442
rect 228968 109384 231490 109440
rect 231546 109384 231551 109440
rect 228968 109382 231551 109384
rect 231485 109379 231551 109382
rect 265709 109306 265775 109309
rect 268150 109306 268210 109548
rect 279926 109518 291148 109578
rect 291142 109516 291148 109518
rect 291212 109516 291218 109580
rect 265709 109304 268210 109306
rect 265709 109248 265714 109304
rect 265770 109248 268210 109304
rect 265709 109246 268210 109248
rect 265709 109243 265775 109246
rect 213913 109168 217242 109170
rect 213913 109112 213918 109168
rect 213974 109112 217242 109168
rect 213913 109110 217242 109112
rect 279926 109170 279986 109412
rect 295374 109170 295380 109172
rect 279926 109110 295380 109170
rect 213913 109107 213979 109110
rect 295374 109108 295380 109110
rect 295444 109108 295450 109172
rect 231761 108898 231827 108901
rect 228968 108896 231827 108898
rect 167913 108762 167979 108765
rect 164694 108760 167979 108762
rect 164694 108704 167918 108760
rect 167974 108704 167979 108760
rect 164694 108702 167979 108704
rect 167913 108699 167979 108702
rect 214741 108490 214807 108493
rect 200070 108488 214807 108490
rect 200070 108432 214746 108488
rect 214802 108432 214807 108488
rect 200070 108430 214807 108432
rect 170438 108292 170444 108356
rect 170508 108354 170514 108356
rect 200070 108354 200130 108430
rect 214741 108427 214807 108430
rect 170508 108294 200130 108354
rect 214005 108354 214071 108357
rect 217182 108354 217242 108868
rect 228968 108840 231766 108896
rect 231822 108840 231827 108896
rect 228968 108838 231827 108840
rect 231761 108835 231827 108838
rect 265709 108762 265775 108765
rect 268150 108762 268210 109004
rect 265709 108760 268210 108762
rect 265709 108704 265714 108760
rect 265770 108704 268210 108760
rect 265709 108702 268210 108704
rect 265709 108699 265775 108702
rect 282821 108626 282887 108629
rect 279956 108624 282887 108626
rect 231117 108490 231183 108493
rect 228968 108488 231183 108490
rect 228968 108432 231122 108488
rect 231178 108432 231183 108488
rect 228968 108430 231183 108432
rect 231117 108427 231183 108430
rect 214005 108352 217242 108354
rect 214005 108296 214010 108352
rect 214066 108296 217242 108352
rect 214005 108294 217242 108296
rect 265433 108354 265499 108357
rect 268150 108354 268210 108596
rect 279956 108568 282826 108624
rect 282882 108568 282887 108624
rect 279956 108566 282887 108568
rect 282821 108563 282887 108566
rect 265433 108352 268210 108354
rect 265433 108296 265438 108352
rect 265494 108296 268210 108352
rect 265433 108294 268210 108296
rect 170508 108292 170514 108294
rect 214005 108291 214071 108294
rect 265433 108291 265499 108294
rect 213913 107946 213979 107949
rect 217182 107946 217242 108188
rect 231669 107946 231735 107949
rect 213913 107944 217242 107946
rect 213913 107888 213918 107944
rect 213974 107888 217242 107944
rect 213913 107886 217242 107888
rect 228968 107944 231735 107946
rect 228968 107888 231674 107944
rect 231730 107888 231735 107944
rect 228968 107886 231735 107888
rect 213913 107883 213979 107886
rect 231669 107883 231735 107886
rect 265341 107946 265407 107949
rect 268334 107948 268394 108188
rect 265341 107944 268210 107946
rect 265341 107888 265346 107944
rect 265402 107888 268210 107944
rect 265341 107886 268210 107888
rect 265341 107883 265407 107886
rect 268150 107780 268210 107886
rect 268326 107884 268332 107948
rect 268396 107884 268402 107948
rect 281533 107810 281599 107813
rect 279956 107808 281599 107810
rect 279956 107752 281538 107808
rect 281594 107752 281599 107808
rect 279956 107750 281599 107752
rect 281533 107747 281599 107750
rect 231761 107538 231827 107541
rect 228968 107536 231827 107538
rect 214005 106994 214071 106997
rect 217182 106994 217242 107508
rect 228968 107480 231766 107536
rect 231822 107480 231827 107536
rect 228968 107478 231827 107480
rect 231761 107475 231827 107478
rect 264237 107538 264303 107541
rect 268326 107538 268332 107540
rect 264237 107536 268332 107538
rect 264237 107480 264242 107536
rect 264298 107480 268332 107536
rect 264237 107478 268332 107480
rect 264237 107475 264303 107478
rect 268326 107476 268332 107478
rect 268396 107476 268402 107540
rect 231577 107130 231643 107133
rect 228968 107128 231643 107130
rect 228968 107072 231582 107128
rect 231638 107072 231643 107128
rect 228968 107070 231643 107072
rect 231577 107067 231643 107070
rect 265525 107130 265591 107133
rect 268150 107130 268210 107372
rect 280245 107130 280311 107133
rect 265525 107128 268210 107130
rect 265525 107072 265530 107128
rect 265586 107072 268210 107128
rect 265525 107070 268210 107072
rect 279956 107128 280311 107130
rect 279956 107072 280250 107128
rect 280306 107072 280311 107128
rect 279956 107070 280311 107072
rect 265525 107067 265591 107070
rect 280245 107067 280311 107070
rect 214005 106992 217242 106994
rect 214005 106936 214010 106992
rect 214066 106936 217242 106992
rect 214005 106934 217242 106936
rect 214005 106931 214071 106934
rect 213913 106586 213979 106589
rect 217182 106586 217242 106828
rect 265801 106722 265867 106725
rect 268150 106722 268210 106964
rect 265801 106720 268210 106722
rect 265801 106664 265806 106720
rect 265862 106664 268210 106720
rect 265801 106662 268210 106664
rect 265801 106659 265867 106662
rect 230565 106586 230631 106589
rect 213913 106584 217242 106586
rect 213913 106528 213918 106584
rect 213974 106528 217242 106584
rect 213913 106526 217242 106528
rect 228968 106584 230631 106586
rect 228968 106528 230570 106584
rect 230626 106528 230631 106584
rect 228968 106526 230631 106528
rect 213913 106523 213979 106526
rect 230565 106523 230631 106526
rect 265709 106586 265775 106589
rect 265709 106584 268210 106586
rect 265709 106528 265714 106584
rect 265770 106528 268210 106584
rect 265709 106526 268210 106528
rect 265709 106523 265775 106526
rect 268150 106420 268210 106526
rect 282453 106314 282519 106317
rect 279956 106312 282519 106314
rect 279956 106256 282458 106312
rect 282514 106256 282519 106312
rect 279956 106254 282519 106256
rect 282453 106251 282519 106254
rect 231669 106178 231735 106181
rect 228968 106176 231735 106178
rect 214005 105770 214071 105773
rect 217182 105770 217242 106148
rect 228968 106120 231674 106176
rect 231730 106120 231735 106176
rect 228968 106118 231735 106120
rect 231669 106115 231735 106118
rect 214005 105768 217242 105770
rect 214005 105712 214010 105768
rect 214066 105712 217242 105768
rect 214005 105710 217242 105712
rect 265709 105770 265775 105773
rect 268150 105770 268210 106012
rect 265709 105768 268210 105770
rect 265709 105712 265714 105768
rect 265770 105712 268210 105768
rect 265709 105710 268210 105712
rect 214005 105707 214071 105710
rect 265709 105707 265775 105710
rect 231761 105634 231827 105637
rect 228968 105632 231827 105634
rect 213913 105362 213979 105365
rect 217182 105362 217242 105604
rect 228968 105576 231766 105632
rect 231822 105576 231827 105632
rect 228968 105574 231827 105576
rect 231761 105571 231827 105574
rect 213913 105360 217242 105362
rect 213913 105304 213918 105360
rect 213974 105304 217242 105360
rect 213913 105302 217242 105304
rect 265801 105362 265867 105365
rect 268150 105362 268210 105604
rect 282821 105498 282887 105501
rect 279956 105496 282887 105498
rect 279956 105440 282826 105496
rect 282882 105440 282887 105496
rect 279956 105438 282887 105440
rect 282821 105435 282887 105438
rect 265801 105360 268210 105362
rect 265801 105304 265806 105360
rect 265862 105304 268210 105360
rect 265801 105302 268210 105304
rect 213913 105299 213979 105302
rect 265801 105299 265867 105302
rect 213453 105226 213519 105229
rect 230841 105226 230907 105229
rect 213453 105224 217426 105226
rect 213453 105168 213458 105224
rect 213514 105168 217426 105224
rect 213453 105166 217426 105168
rect 228968 105224 230907 105226
rect 228968 105168 230846 105224
rect 230902 105168 230907 105224
rect 228968 105166 230907 105168
rect 213453 105163 213519 105166
rect 217366 104924 217426 105166
rect 230841 105163 230907 105166
rect 266077 104954 266143 104957
rect 268334 104954 268394 105196
rect 266077 104952 268394 104954
rect 266077 104896 266082 104952
rect 266138 104896 268394 104952
rect 266077 104894 268394 104896
rect 282453 104954 282519 104957
rect 288382 104954 288388 104956
rect 282453 104952 288388 104954
rect 282453 104896 282458 104952
rect 282514 104896 288388 104952
rect 282453 104894 288388 104896
rect 266077 104891 266143 104894
rect 282453 104891 282519 104894
rect 288382 104892 288388 104894
rect 288452 104892 288458 104956
rect 280337 104818 280403 104821
rect 279956 104816 280403 104818
rect 231577 104682 231643 104685
rect 228968 104680 231643 104682
rect 228968 104624 231582 104680
rect 231638 104624 231643 104680
rect 228968 104622 231643 104624
rect 231577 104619 231643 104622
rect 264421 104546 264487 104549
rect 268150 104546 268210 104788
rect 279956 104760 280342 104816
rect 280398 104760 280403 104816
rect 279956 104758 280403 104760
rect 280337 104755 280403 104758
rect 264421 104544 268210 104546
rect 264421 104488 264426 104544
rect 264482 104488 268210 104544
rect 264421 104486 268210 104488
rect 264421 104483 264487 104486
rect 231761 104274 231827 104277
rect 228968 104272 231827 104274
rect 213913 103730 213979 103733
rect 217182 103730 217242 104244
rect 228968 104216 231766 104272
rect 231822 104216 231827 104272
rect 228968 104214 231827 104216
rect 231761 104211 231827 104214
rect 266077 104002 266143 104005
rect 268150 104002 268210 104380
rect 284334 104002 284340 104004
rect 266077 104000 268210 104002
rect 266077 103944 266082 104000
rect 266138 103944 268210 104000
rect 266077 103942 268210 103944
rect 279956 103942 284340 104002
rect 266077 103939 266143 103942
rect 284334 103940 284340 103942
rect 284404 103940 284410 104004
rect 231025 103730 231091 103733
rect 213913 103728 217242 103730
rect 213913 103672 213918 103728
rect 213974 103672 217242 103728
rect 213913 103670 217242 103672
rect 228968 103728 231091 103730
rect 228968 103672 231030 103728
rect 231086 103672 231091 103728
rect 228968 103670 231091 103672
rect 213913 103667 213979 103670
rect 231025 103667 231091 103670
rect 214414 103532 214420 103596
rect 214484 103594 214490 103596
rect 265801 103594 265867 103597
rect 268150 103594 268210 103836
rect 214484 103534 217058 103594
rect 265801 103592 268210 103594
rect 214484 103532 214490 103534
rect 216998 103530 217058 103534
rect 217182 103530 217242 103564
rect 265801 103536 265806 103592
rect 265862 103536 268210 103592
rect 265801 103534 268210 103536
rect 265801 103531 265867 103534
rect 216998 103470 217242 103530
rect 231577 103322 231643 103325
rect 228968 103320 231643 103322
rect 228968 103264 231582 103320
rect 231638 103264 231643 103320
rect 228968 103262 231643 103264
rect 231577 103259 231643 103262
rect 265709 103186 265775 103189
rect 268150 103186 268210 103428
rect 282821 103186 282887 103189
rect 265709 103184 268210 103186
rect 265709 103128 265714 103184
rect 265770 103128 268210 103184
rect 265709 103126 268210 103128
rect 279956 103184 282887 103186
rect 279956 103128 282826 103184
rect 282882 103128 282887 103184
rect 279956 103126 282887 103128
rect 265709 103123 265775 103126
rect 282821 103123 282887 103126
rect 217182 102642 217242 102884
rect 231761 102778 231827 102781
rect 228968 102776 231827 102778
rect 228968 102720 231766 102776
rect 231822 102720 231827 102776
rect 228968 102718 231827 102720
rect 231761 102715 231827 102718
rect 262070 102716 262076 102780
rect 262140 102778 262146 102780
rect 268150 102778 268210 103020
rect 262140 102718 268210 102778
rect 262140 102716 262146 102718
rect 268326 102716 268332 102780
rect 268396 102716 268402 102780
rect 200070 102582 217242 102642
rect 268334 102612 268394 102716
rect 68142 102316 68816 102376
rect 64781 102234 64847 102237
rect 68142 102234 68202 102316
rect 172094 102308 172100 102372
rect 172164 102370 172170 102372
rect 200070 102370 200130 102582
rect 214741 102506 214807 102509
rect 214741 102504 217426 102506
rect 214741 102448 214746 102504
rect 214802 102448 217426 102504
rect 214741 102446 217426 102448
rect 214741 102443 214807 102446
rect 172164 102310 200130 102370
rect 172164 102308 172170 102310
rect 64781 102232 68202 102234
rect 64781 102176 64786 102232
rect 64842 102176 68202 102232
rect 217366 102204 217426 102446
rect 253054 102444 253060 102508
rect 253124 102506 253130 102508
rect 267774 102506 267780 102508
rect 253124 102446 267780 102506
rect 253124 102444 253130 102446
rect 267774 102444 267780 102446
rect 267844 102444 267850 102508
rect 282453 102506 282519 102509
rect 279956 102504 282519 102506
rect 279956 102448 282458 102504
rect 282514 102448 282519 102504
rect 279956 102446 282519 102448
rect 282453 102443 282519 102446
rect 231301 102370 231367 102373
rect 228968 102368 231367 102370
rect 228968 102312 231306 102368
rect 231362 102312 231367 102368
rect 228968 102310 231367 102312
rect 231301 102307 231367 102310
rect 265801 102370 265867 102373
rect 265801 102368 268210 102370
rect 265801 102312 265806 102368
rect 265862 102312 268210 102368
rect 265801 102310 268210 102312
rect 265801 102307 265867 102310
rect 268150 102204 268210 102310
rect 64781 102174 68202 102176
rect 64781 102171 64847 102174
rect 265525 101962 265591 101965
rect 265525 101960 268210 101962
rect 265525 101904 265530 101960
rect 265586 101904 268210 101960
rect 265525 101902 268210 101904
rect 265525 101899 265591 101902
rect 229921 101826 229987 101829
rect 228968 101824 229987 101826
rect 228968 101768 229926 101824
rect 229982 101768 229987 101824
rect 268150 101796 268210 101902
rect 228968 101766 229987 101768
rect 229921 101763 229987 101766
rect 281625 101690 281691 101693
rect 279956 101688 281691 101690
rect 279956 101632 281630 101688
rect 281686 101632 281691 101688
rect 279956 101630 281691 101632
rect 281625 101627 281691 101630
rect 265709 101554 265775 101557
rect 265709 101552 268394 101554
rect 214005 101282 214071 101285
rect 217182 101282 217242 101524
rect 265709 101496 265714 101552
rect 265770 101496 268394 101552
rect 265709 101494 268394 101496
rect 265709 101491 265775 101494
rect 231117 101418 231183 101421
rect 228968 101416 231183 101418
rect 228968 101360 231122 101416
rect 231178 101360 231183 101416
rect 228968 101358 231183 101360
rect 231117 101355 231183 101358
rect 214005 101280 217242 101282
rect 214005 101224 214010 101280
rect 214066 101224 217242 101280
rect 268334 101252 268394 101494
rect 214005 101222 217242 101224
rect 214005 101219 214071 101222
rect 213913 101146 213979 101149
rect 213913 101144 217242 101146
rect 213913 101088 213918 101144
rect 213974 101088 217242 101144
rect 213913 101086 217242 101088
rect 213913 101083 213979 101086
rect 217182 100980 217242 101086
rect 265801 101010 265867 101013
rect 265801 101008 268210 101010
rect 265801 100952 265806 101008
rect 265862 100952 268210 101008
rect 265801 100950 268210 100952
rect 265801 100947 265867 100950
rect 230565 100874 230631 100877
rect 228968 100872 230631 100874
rect 228968 100816 230570 100872
rect 230626 100816 230631 100872
rect 268150 100844 268210 100950
rect 281809 100874 281875 100877
rect 279956 100872 281875 100874
rect 228968 100814 230631 100816
rect 279956 100816 281814 100872
rect 281870 100816 281875 100872
rect 279956 100814 281875 100816
rect 230565 100811 230631 100814
rect 281809 100811 281875 100814
rect 67725 100738 67791 100741
rect 68142 100738 68816 100744
rect 67725 100736 68816 100738
rect 67725 100680 67730 100736
rect 67786 100684 68816 100736
rect 67786 100680 68202 100684
rect 67725 100678 68202 100680
rect 67725 100675 67791 100678
rect 231761 100466 231827 100469
rect 228968 100464 231827 100466
rect 228968 100408 231766 100464
rect 231822 100408 231827 100464
rect 228968 100406 231827 100408
rect 231761 100403 231827 100406
rect 213913 99786 213979 99789
rect 217182 99786 217242 100300
rect 265709 100194 265775 100197
rect 268150 100194 268210 100436
rect 281533 100194 281599 100197
rect 265709 100192 268210 100194
rect 265709 100136 265714 100192
rect 265770 100136 268210 100192
rect 265709 100134 268210 100136
rect 279956 100192 281599 100194
rect 279956 100136 281538 100192
rect 281594 100136 281599 100192
rect 279956 100134 281599 100136
rect 265709 100131 265775 100134
rect 281533 100131 281599 100134
rect 231669 99922 231735 99925
rect 228968 99920 231735 99922
rect 228968 99864 231674 99920
rect 231730 99864 231735 99920
rect 228968 99862 231735 99864
rect 231669 99859 231735 99862
rect 213913 99784 217242 99786
rect 213913 99728 213918 99784
rect 213974 99728 217242 99784
rect 213913 99726 217242 99728
rect 265801 99786 265867 99789
rect 268150 99786 268210 100028
rect 265801 99784 268210 99786
rect 265801 99728 265806 99784
rect 265862 99728 268210 99784
rect 265801 99726 268210 99728
rect 213913 99723 213979 99726
rect 265801 99723 265867 99726
rect 214097 99514 214163 99517
rect 214097 99512 216874 99514
rect 214097 99456 214102 99512
rect 214158 99456 216874 99512
rect 214097 99454 216874 99456
rect 214097 99451 214163 99454
rect 216814 99378 216874 99454
rect 217366 99378 217426 99620
rect 231393 99514 231459 99517
rect 228968 99512 231459 99514
rect 228968 99456 231398 99512
rect 231454 99456 231459 99512
rect 228968 99454 231459 99456
rect 231393 99451 231459 99454
rect 265525 99514 265591 99517
rect 265525 99512 267842 99514
rect 265525 99456 265530 99512
rect 265586 99456 267842 99512
rect 265525 99454 267842 99456
rect 265525 99451 265591 99454
rect 216814 99318 217426 99378
rect 267782 99378 267842 99454
rect 268334 99378 268394 99620
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 282821 99378 282887 99381
rect 267782 99318 268394 99378
rect 279956 99376 282887 99378
rect 279956 99320 282826 99376
rect 282882 99320 282887 99376
rect 583520 99364 584960 99454
rect 279956 99318 282887 99320
rect 282821 99315 282887 99318
rect 230657 98970 230723 98973
rect 228968 98968 230723 98970
rect 214005 98426 214071 98429
rect 217182 98426 217242 98940
rect 228968 98912 230662 98968
rect 230718 98912 230723 98968
rect 228968 98910 230723 98912
rect 230657 98907 230723 98910
rect 266854 98772 266860 98836
rect 266924 98834 266930 98836
rect 268150 98834 268210 99212
rect 266924 98774 268210 98834
rect 266924 98772 266930 98774
rect 231485 98562 231551 98565
rect 228968 98560 231551 98562
rect 228968 98504 231490 98560
rect 231546 98504 231551 98560
rect 228968 98502 231551 98504
rect 231485 98499 231551 98502
rect 214005 98424 217242 98426
rect 214005 98368 214010 98424
rect 214066 98368 217242 98424
rect 214005 98366 217242 98368
rect 265801 98426 265867 98429
rect 268150 98426 268210 98668
rect 265801 98424 268210 98426
rect 265801 98368 265806 98424
rect 265862 98368 268210 98424
rect 265801 98366 268210 98368
rect 214005 98363 214071 98366
rect 265801 98363 265867 98366
rect 213913 98018 213979 98021
rect 217366 98018 217426 98260
rect 233734 98018 233740 98020
rect 213913 98016 217426 98018
rect 213913 97960 213918 98016
rect 213974 97960 217426 98016
rect 213913 97958 217426 97960
rect 228968 97958 233740 98018
rect 213913 97955 213979 97958
rect 233734 97956 233740 97958
rect 233804 97956 233810 98020
rect 265433 98018 265499 98021
rect 268334 98018 268394 98260
rect 279374 98157 279434 98532
rect 279374 98152 279483 98157
rect 279374 98096 279422 98152
rect 279478 98096 279483 98152
rect 279374 98094 279483 98096
rect 279417 98091 279483 98094
rect 265433 98016 268394 98018
rect 265433 97960 265438 98016
rect 265494 97960 268394 98016
rect 265433 97958 268394 97960
rect 265433 97955 265499 97958
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect 230473 97610 230539 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect 228968 97608 230539 97610
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 213913 97066 213979 97069
rect 217182 97066 217242 97580
rect 228968 97552 230478 97608
rect 230534 97552 230539 97608
rect 228968 97550 230539 97552
rect 230473 97547 230539 97550
rect 265801 97610 265867 97613
rect 268150 97610 268210 97852
rect 265801 97608 268210 97610
rect 265801 97552 265806 97608
rect 265862 97552 268210 97608
rect 265801 97550 268210 97552
rect 265801 97547 265867 97550
rect 265157 97202 265223 97205
rect 268150 97202 268210 97444
rect 279558 97341 279618 97852
rect 279509 97336 279618 97341
rect 279509 97280 279514 97336
rect 279570 97280 279618 97336
rect 279509 97278 279618 97280
rect 279509 97275 279575 97278
rect 265157 97200 268210 97202
rect 265157 97144 265162 97200
rect 265218 97144 268210 97200
rect 265157 97142 268210 97144
rect 265157 97139 265223 97142
rect 229134 97066 229140 97068
rect 213913 97064 217242 97066
rect 213913 97008 213918 97064
rect 213974 97008 217242 97064
rect 213913 97006 217242 97008
rect 228968 97006 229140 97066
rect 213913 97003 213979 97006
rect 229134 97004 229140 97006
rect 229204 97066 229210 97068
rect 230473 97066 230539 97069
rect 229204 97064 230539 97066
rect 229204 97008 230478 97064
rect 230534 97008 230539 97064
rect 229204 97006 230539 97008
rect 229204 97004 229210 97006
rect 230473 97003 230539 97006
rect 214833 96658 214899 96661
rect 217182 96658 217242 96900
rect 263550 96734 268210 96794
rect 231117 96658 231183 96661
rect 214833 96656 217242 96658
rect 214833 96600 214838 96656
rect 214894 96600 217242 96656
rect 214833 96598 217242 96600
rect 228968 96656 231183 96658
rect 228968 96600 231122 96656
rect 231178 96600 231183 96656
rect 228968 96598 231183 96600
rect 214833 96595 214899 96598
rect 231117 96595 231183 96598
rect 253238 96596 253244 96660
rect 253308 96658 253314 96660
rect 263550 96658 263610 96734
rect 253308 96598 263610 96658
rect 253308 96596 253314 96598
rect 265750 96596 265756 96660
rect 265820 96658 265826 96660
rect 267774 96658 267780 96660
rect 265820 96598 267780 96658
rect 265820 96596 265826 96598
rect 267774 96596 267780 96598
rect 267844 96596 267850 96660
rect 268150 96628 268210 96734
rect 268326 96732 268332 96796
rect 268396 96794 268402 96796
rect 268518 96794 268578 97036
rect 268396 96734 268578 96794
rect 268396 96732 268402 96734
rect 279374 96661 279434 97036
rect 279325 96656 279434 96661
rect 279325 96600 279330 96656
rect 279386 96600 279434 96656
rect 279325 96598 279434 96600
rect 279325 96595 279391 96598
rect 265801 96386 265867 96389
rect 265801 96384 268210 96386
rect 166942 95780 166948 95844
rect 167012 95842 167018 95844
rect 214097 95842 214163 95845
rect 167012 95840 214163 95842
rect 167012 95784 214102 95840
rect 214158 95784 214163 95840
rect 167012 95782 214163 95784
rect 167012 95780 167018 95782
rect 214097 95779 214163 95782
rect 214557 95842 214623 95845
rect 217182 95842 217242 96356
rect 265801 96328 265806 96384
rect 265862 96328 268210 96384
rect 265801 96326 268210 96328
rect 265801 96323 265867 96326
rect 268150 96220 268210 96326
rect 214557 95840 217242 95842
rect 214557 95784 214562 95840
rect 214618 95784 217242 95840
rect 214557 95782 217242 95784
rect 214557 95779 214623 95782
rect 228774 95706 228834 96220
rect 267181 95978 267247 95981
rect 279325 95978 279391 95981
rect 267181 95976 279391 95978
rect 267181 95920 267186 95976
rect 267242 95920 279330 95976
rect 279386 95920 279391 95976
rect 267181 95918 279391 95920
rect 267181 95915 267247 95918
rect 279325 95915 279391 95918
rect 279926 95842 279986 96356
rect 280061 95842 280127 95845
rect 279926 95840 280127 95842
rect 279926 95784 280066 95840
rect 280122 95784 280127 95840
rect 279926 95782 280127 95784
rect 280061 95779 280127 95782
rect 230473 95706 230539 95709
rect 228774 95704 230539 95706
rect 228774 95648 230478 95704
rect 230534 95648 230539 95704
rect 228774 95646 230539 95648
rect 230473 95643 230539 95646
rect 227662 95236 227668 95300
rect 227732 95298 227738 95300
rect 228950 95298 228956 95300
rect 227732 95238 228956 95298
rect 227732 95236 227738 95238
rect 228950 95236 228956 95238
rect 229020 95236 229026 95300
rect 195830 95100 195836 95164
rect 195900 95162 195906 95164
rect 279417 95162 279483 95165
rect 195900 95160 279483 95162
rect 195900 95104 279422 95160
rect 279478 95104 279483 95160
rect 195900 95102 279483 95104
rect 195900 95100 195906 95102
rect 279417 95099 279483 95102
rect 66069 94890 66135 94893
rect 204989 94890 205055 94893
rect 66069 94888 205055 94890
rect 66069 94832 66074 94888
rect 66130 94832 204994 94888
rect 205050 94832 205055 94888
rect 66069 94830 205055 94832
rect 66069 94827 66135 94830
rect 204989 94827 205055 94830
rect 105721 94756 105787 94757
rect 112345 94756 112411 94757
rect 105656 94692 105662 94756
rect 105726 94754 105787 94756
rect 105726 94752 105818 94754
rect 105782 94696 105818 94752
rect 105726 94694 105818 94696
rect 105726 94692 105787 94694
rect 112320 94692 112326 94756
rect 112390 94754 112411 94756
rect 128077 94756 128143 94757
rect 151721 94756 151787 94757
rect 128077 94754 128102 94756
rect 112390 94752 112482 94754
rect 112406 94696 112482 94752
rect 112390 94694 112482 94696
rect 128010 94752 128102 94754
rect 128010 94696 128082 94752
rect 128010 94694 128102 94696
rect 112390 94692 112411 94694
rect 105721 94691 105787 94692
rect 112345 94691 112411 94692
rect 128077 94692 128102 94694
rect 128166 94692 128172 94756
rect 151721 94754 151766 94756
rect 151674 94752 151766 94754
rect 151674 94696 151726 94752
rect 151674 94694 151766 94696
rect 151721 94692 151766 94694
rect 151830 94692 151836 94756
rect 128077 94691 128143 94692
rect 151721 94691 151787 94692
rect 106457 94076 106523 94077
rect 106406 94012 106412 94076
rect 106476 94074 106523 94076
rect 106476 94072 106568 94074
rect 106518 94016 106568 94072
rect 106476 94014 106568 94016
rect 106476 94012 106523 94014
rect 106457 94011 106523 94012
rect 66161 93802 66227 93805
rect 213453 93802 213519 93805
rect 66161 93800 213519 93802
rect 66161 93744 66166 93800
rect 66222 93744 213458 93800
rect 213514 93744 213519 93800
rect 66161 93742 213519 93744
rect 66161 93739 66227 93742
rect 213453 93739 213519 93742
rect 121729 93668 121795 93669
rect 121678 93666 121684 93668
rect 121638 93606 121684 93666
rect 121748 93664 121795 93668
rect 171961 93666 172027 93669
rect 121790 93608 121795 93664
rect 121678 93604 121684 93606
rect 121748 93604 121795 93608
rect 121729 93603 121795 93604
rect 122790 93664 172027 93666
rect 122790 93608 171966 93664
rect 172022 93608 172027 93664
rect 122790 93606 172027 93608
rect 88977 93532 89043 93533
rect 111241 93532 111307 93533
rect 88926 93530 88932 93532
rect 88886 93470 88932 93530
rect 88996 93528 89043 93532
rect 111190 93530 111196 93532
rect 89038 93472 89043 93528
rect 88926 93468 88932 93470
rect 88996 93468 89043 93472
rect 111150 93470 111196 93530
rect 111260 93528 111307 93532
rect 111302 93472 111307 93528
rect 111190 93468 111196 93470
rect 111260 93468 111307 93472
rect 119286 93468 119292 93532
rect 119356 93530 119362 93532
rect 122790 93530 122850 93606
rect 171961 93603 172027 93606
rect 195646 93604 195652 93668
rect 195716 93666 195722 93668
rect 280061 93666 280127 93669
rect 195716 93664 280127 93666
rect 195716 93608 280066 93664
rect 280122 93608 280127 93664
rect 195716 93606 280127 93608
rect 195716 93604 195722 93606
rect 280061 93603 280127 93606
rect 134425 93532 134491 93533
rect 134374 93530 134380 93532
rect 119356 93470 122850 93530
rect 134334 93470 134380 93530
rect 134444 93528 134491 93532
rect 134486 93472 134491 93528
rect 119356 93468 119362 93470
rect 134374 93468 134380 93470
rect 134444 93468 134491 93472
rect 197118 93468 197124 93532
rect 197188 93530 197194 93532
rect 280245 93530 280311 93533
rect 197188 93528 280311 93530
rect 197188 93472 280250 93528
rect 280306 93472 280311 93528
rect 197188 93470 280311 93472
rect 197188 93468 197194 93470
rect 88977 93467 89043 93468
rect 111241 93467 111307 93468
rect 134425 93467 134491 93468
rect 280245 93467 280311 93470
rect 103278 93196 103284 93260
rect 103348 93258 103354 93260
rect 103421 93258 103487 93261
rect 110137 93260 110203 93261
rect 110086 93258 110092 93260
rect 103348 93256 103487 93258
rect 103348 93200 103426 93256
rect 103482 93200 103487 93256
rect 103348 93198 103487 93200
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 110198 93200 110203 93256
rect 103348 93196 103354 93198
rect 103421 93195 103487 93198
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 110137 93195 110203 93196
rect 85798 92380 85804 92444
rect 85868 92442 85874 92444
rect 86585 92442 86651 92445
rect 98545 92444 98611 92445
rect 98494 92442 98500 92444
rect 85868 92440 86651 92442
rect 85868 92384 86590 92440
rect 86646 92384 86651 92440
rect 85868 92382 86651 92384
rect 98454 92382 98500 92442
rect 98564 92440 98611 92444
rect 98606 92384 98611 92440
rect 85868 92380 85874 92382
rect 86585 92379 86651 92382
rect 98494 92380 98500 92382
rect 98564 92380 98611 92384
rect 104198 92380 104204 92444
rect 104268 92442 104274 92444
rect 104341 92442 104407 92445
rect 104617 92444 104683 92445
rect 106641 92444 106707 92445
rect 110689 92444 110755 92445
rect 118049 92444 118115 92445
rect 126697 92444 126763 92445
rect 133137 92444 133203 92445
rect 151537 92444 151603 92445
rect 104566 92442 104572 92444
rect 104268 92440 104407 92442
rect 104268 92384 104346 92440
rect 104402 92384 104407 92440
rect 104268 92382 104407 92384
rect 104526 92382 104572 92442
rect 104636 92440 104683 92444
rect 106590 92442 106596 92444
rect 104678 92384 104683 92440
rect 104268 92380 104274 92382
rect 98545 92379 98611 92380
rect 104341 92379 104407 92382
rect 104566 92380 104572 92382
rect 104636 92380 104683 92384
rect 106550 92382 106596 92442
rect 106660 92440 106707 92444
rect 110638 92442 110644 92444
rect 106702 92384 106707 92440
rect 106590 92380 106596 92382
rect 106660 92380 106707 92384
rect 110598 92382 110644 92442
rect 110708 92440 110755 92444
rect 117998 92442 118004 92444
rect 110750 92384 110755 92440
rect 110638 92380 110644 92382
rect 110708 92380 110755 92384
rect 117958 92382 118004 92442
rect 118068 92440 118115 92444
rect 126646 92442 126652 92444
rect 118110 92384 118115 92440
rect 117998 92380 118004 92382
rect 118068 92380 118115 92384
rect 126606 92382 126652 92442
rect 126716 92440 126763 92444
rect 133086 92442 133092 92444
rect 126758 92384 126763 92440
rect 126646 92380 126652 92382
rect 126716 92380 126763 92384
rect 133046 92382 133092 92442
rect 133156 92440 133203 92444
rect 151486 92442 151492 92444
rect 133198 92384 133203 92440
rect 133086 92380 133092 92382
rect 133156 92380 133203 92384
rect 151446 92382 151492 92442
rect 151556 92440 151603 92444
rect 151598 92384 151603 92440
rect 151486 92380 151492 92382
rect 151556 92380 151603 92384
rect 104617 92379 104683 92380
rect 106641 92379 106707 92380
rect 110689 92379 110755 92380
rect 118049 92379 118115 92380
rect 126697 92379 126763 92380
rect 133137 92379 133203 92380
rect 151537 92379 151603 92380
rect 113030 92244 113036 92308
rect 113100 92306 113106 92308
rect 170438 92306 170444 92308
rect 113100 92246 170444 92306
rect 113100 92244 113106 92246
rect 170438 92244 170444 92246
rect 170508 92244 170514 92308
rect 88006 92108 88012 92172
rect 88076 92170 88082 92172
rect 166942 92170 166948 92172
rect 88076 92110 166948 92170
rect 88076 92108 88082 92110
rect 166942 92108 166948 92110
rect 167012 92108 167018 92172
rect 115473 92036 115539 92037
rect 126513 92036 126579 92037
rect 151353 92036 151419 92037
rect 115422 92034 115428 92036
rect 115382 91974 115428 92034
rect 115492 92032 115539 92036
rect 126462 92034 126468 92036
rect 115534 91976 115539 92032
rect 115422 91972 115428 91974
rect 115492 91972 115539 91976
rect 126422 91974 126468 92034
rect 126532 92032 126579 92036
rect 151302 92034 151308 92036
rect 126574 91976 126579 92032
rect 126462 91972 126468 91974
rect 126532 91972 126579 91976
rect 151262 91974 151308 92034
rect 151372 92032 151419 92036
rect 151414 91976 151419 92032
rect 151302 91972 151308 91974
rect 151372 91972 151419 91976
rect 115473 91971 115539 91972
rect 126513 91971 126579 91972
rect 151353 91971 151419 91972
rect 90214 91700 90220 91764
rect 90284 91762 90290 91764
rect 90357 91762 90423 91765
rect 90284 91760 90423 91762
rect 90284 91704 90362 91760
rect 90418 91704 90423 91760
rect 90284 91702 90423 91704
rect 90284 91700 90290 91702
rect 90357 91699 90423 91702
rect 119654 91700 119660 91764
rect 119724 91762 119730 91764
rect 119889 91762 119955 91765
rect 119724 91760 119955 91762
rect 119724 91704 119894 91760
rect 119950 91704 119955 91760
rect 119724 91702 119955 91704
rect 119724 91700 119730 91702
rect 119889 91699 119955 91702
rect 105486 91564 105492 91628
rect 105556 91626 105562 91628
rect 105997 91626 106063 91629
rect 132401 91628 132467 91629
rect 132350 91626 132356 91628
rect 105556 91624 106063 91626
rect 105556 91568 106002 91624
rect 106058 91568 106063 91624
rect 105556 91566 106063 91568
rect 132310 91566 132356 91626
rect 132420 91624 132467 91628
rect 132462 91568 132467 91624
rect 105556 91564 105562 91566
rect 105997 91563 106063 91566
rect 132350 91564 132356 91566
rect 132420 91564 132467 91568
rect 132401 91563 132467 91564
rect 101857 91492 101923 91493
rect 101806 91490 101812 91492
rect 101766 91430 101812 91490
rect 101876 91488 101923 91492
rect 101918 91432 101923 91488
rect 101806 91428 101812 91430
rect 101876 91428 101923 91432
rect 109166 91428 109172 91492
rect 109236 91490 109242 91492
rect 109493 91490 109559 91493
rect 109236 91488 109559 91490
rect 109236 91432 109498 91488
rect 109554 91432 109559 91488
rect 109236 91430 109559 91432
rect 109236 91428 109242 91430
rect 101857 91427 101923 91428
rect 109493 91427 109559 91430
rect 122782 91428 122788 91492
rect 122852 91490 122858 91492
rect 124121 91490 124187 91493
rect 122852 91488 124187 91490
rect 122852 91432 124126 91488
rect 124182 91432 124187 91488
rect 122852 91430 124187 91432
rect 122852 91428 122858 91430
rect 124121 91427 124187 91430
rect 93894 91292 93900 91356
rect 93964 91354 93970 91356
rect 95049 91354 95115 91357
rect 93964 91352 95115 91354
rect 93964 91296 95054 91352
rect 95110 91296 95115 91352
rect 93964 91294 95115 91296
rect 93964 91292 93970 91294
rect 95049 91291 95115 91294
rect 98126 91292 98132 91356
rect 98196 91354 98202 91356
rect 99189 91354 99255 91357
rect 100569 91356 100635 91357
rect 100518 91354 100524 91356
rect 98196 91352 99255 91354
rect 98196 91296 99194 91352
rect 99250 91296 99255 91352
rect 98196 91294 99255 91296
rect 100478 91294 100524 91354
rect 100588 91352 100635 91356
rect 100630 91296 100635 91352
rect 98196 91292 98202 91294
rect 99189 91291 99255 91294
rect 100518 91292 100524 91294
rect 100588 91292 100635 91296
rect 100886 91292 100892 91356
rect 100956 91354 100962 91356
rect 101949 91354 102015 91357
rect 100956 91352 102015 91354
rect 100956 91296 101954 91352
rect 102010 91296 102015 91352
rect 100956 91294 102015 91296
rect 100956 91292 100962 91294
rect 100569 91291 100635 91292
rect 101949 91291 102015 91294
rect 107694 91292 107700 91356
rect 107764 91354 107770 91356
rect 108849 91354 108915 91357
rect 114369 91356 114435 91357
rect 117129 91356 117195 91357
rect 114318 91354 114324 91356
rect 107764 91352 108915 91354
rect 107764 91296 108854 91352
rect 108910 91296 108915 91352
rect 107764 91294 108915 91296
rect 114278 91294 114324 91354
rect 114388 91352 114435 91356
rect 117078 91354 117084 91356
rect 114430 91296 114435 91352
rect 107764 91292 107770 91294
rect 108849 91291 108915 91294
rect 114318 91292 114324 91294
rect 114388 91292 114435 91296
rect 117038 91294 117084 91354
rect 117148 91352 117195 91356
rect 117190 91296 117195 91352
rect 117078 91292 117084 91294
rect 117148 91292 117195 91296
rect 120574 91292 120580 91356
rect 120644 91354 120650 91356
rect 120809 91354 120875 91357
rect 125409 91356 125475 91357
rect 125358 91354 125364 91356
rect 120644 91352 120875 91354
rect 120644 91296 120814 91352
rect 120870 91296 120875 91352
rect 120644 91294 120875 91296
rect 125318 91294 125364 91354
rect 125428 91352 125475 91356
rect 125470 91296 125475 91352
rect 120644 91292 120650 91294
rect 114369 91291 114435 91292
rect 117129 91291 117195 91292
rect 120809 91291 120875 91294
rect 125358 91292 125364 91294
rect 125428 91292 125475 91296
rect 125409 91291 125475 91292
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75821 91218 75887 91221
rect 74828 91216 75887 91218
rect 74828 91160 75826 91216
rect 75882 91160 75887 91216
rect 74828 91158 75887 91160
rect 74828 91156 74834 91158
rect 75821 91155 75887 91158
rect 84326 91156 84332 91220
rect 84396 91218 84402 91220
rect 84653 91218 84719 91221
rect 84396 91216 84719 91218
rect 84396 91160 84658 91216
rect 84714 91160 84719 91216
rect 84396 91158 84719 91160
rect 84396 91156 84402 91158
rect 84653 91155 84719 91158
rect 86718 91156 86724 91220
rect 86788 91218 86794 91220
rect 86861 91218 86927 91221
rect 86788 91216 86927 91218
rect 86788 91160 86866 91216
rect 86922 91160 86927 91216
rect 86788 91158 86927 91160
rect 86788 91156 86794 91158
rect 86861 91155 86927 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 92289 91218 92355 91221
rect 91388 91216 92355 91218
rect 91388 91160 92294 91216
rect 92350 91160 92355 91216
rect 91388 91158 92355 91160
rect 91388 91156 91394 91158
rect 92289 91155 92355 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 94998 91156 95004 91220
rect 95068 91218 95074 91220
rect 95141 91218 95207 91221
rect 95068 91216 95207 91218
rect 95068 91160 95146 91216
rect 95202 91160 95207 91216
rect 95068 91158 95207 91160
rect 95068 91156 95074 91158
rect 95141 91155 95207 91158
rect 96286 91156 96292 91220
rect 96356 91218 96362 91220
rect 96521 91218 96587 91221
rect 96356 91216 96587 91218
rect 96356 91160 96526 91216
rect 96582 91160 96587 91216
rect 96356 91158 96587 91160
rect 96356 91156 96362 91158
rect 96521 91155 96587 91158
rect 96654 91156 96660 91220
rect 96724 91218 96730 91220
rect 97073 91218 97139 91221
rect 96724 91216 97139 91218
rect 96724 91160 97078 91216
rect 97134 91160 97139 91216
rect 96724 91158 97139 91160
rect 96724 91156 96730 91158
rect 97073 91155 97139 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97901 91218 97967 91221
rect 97276 91216 97967 91218
rect 97276 91160 97906 91216
rect 97962 91160 97967 91216
rect 97276 91158 97967 91160
rect 97276 91156 97282 91158
rect 97901 91155 97967 91158
rect 99046 91156 99052 91220
rect 99116 91218 99122 91220
rect 99281 91218 99347 91221
rect 99116 91216 99347 91218
rect 99116 91160 99286 91216
rect 99342 91160 99347 91216
rect 99116 91158 99347 91160
rect 99116 91156 99122 91158
rect 99281 91155 99347 91158
rect 99966 91156 99972 91220
rect 100036 91218 100042 91220
rect 100661 91218 100727 91221
rect 102041 91220 102107 91221
rect 101990 91218 101996 91220
rect 100036 91216 100727 91218
rect 100036 91160 100666 91216
rect 100722 91160 100727 91216
rect 100036 91158 100727 91160
rect 101950 91158 101996 91218
rect 102060 91216 102107 91220
rect 102102 91160 102107 91216
rect 100036 91156 100042 91158
rect 100661 91155 100727 91158
rect 101990 91156 101996 91158
rect 102060 91156 102107 91160
rect 102726 91156 102732 91220
rect 102796 91218 102802 91220
rect 103053 91218 103119 91221
rect 102796 91216 103119 91218
rect 102796 91160 103058 91216
rect 103114 91160 103119 91216
rect 102796 91158 103119 91160
rect 102796 91156 102802 91158
rect 102041 91155 102107 91156
rect 103053 91155 103119 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108941 91218 109007 91221
rect 108132 91216 109007 91218
rect 108132 91160 108946 91216
rect 109002 91160 109007 91216
rect 108132 91158 109007 91160
rect 108132 91156 108138 91158
rect 108941 91155 109007 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110321 91218 110387 91221
rect 109604 91216 110387 91218
rect 109604 91160 110326 91216
rect 110382 91160 110387 91216
rect 109604 91158 110387 91160
rect 109604 91156 109610 91158
rect 110321 91155 110387 91158
rect 111926 91156 111932 91220
rect 111996 91218 112002 91220
rect 113081 91218 113147 91221
rect 111996 91216 113147 91218
rect 111996 91160 113086 91216
rect 113142 91160 113147 91216
rect 111996 91158 113147 91160
rect 111996 91156 112002 91158
rect 113081 91155 113147 91158
rect 113214 91156 113220 91220
rect 113284 91218 113290 91220
rect 114461 91218 114527 91221
rect 113284 91216 114527 91218
rect 113284 91160 114466 91216
rect 114522 91160 114527 91216
rect 113284 91158 114527 91160
rect 113284 91156 113290 91158
rect 114461 91155 114527 91158
rect 114870 91156 114876 91220
rect 114940 91218 114946 91220
rect 115565 91218 115631 91221
rect 115841 91220 115907 91221
rect 115790 91218 115796 91220
rect 114940 91216 115631 91218
rect 114940 91160 115570 91216
rect 115626 91160 115631 91216
rect 114940 91158 115631 91160
rect 115750 91158 115796 91218
rect 115860 91216 115907 91220
rect 115902 91160 115907 91216
rect 114940 91156 114946 91158
rect 115565 91155 115631 91158
rect 115790 91156 115796 91158
rect 115860 91156 115907 91160
rect 116710 91156 116716 91220
rect 116780 91218 116786 91220
rect 117221 91218 117287 91221
rect 116780 91216 117287 91218
rect 116780 91160 117226 91216
rect 117282 91160 117287 91216
rect 116780 91158 117287 91160
rect 116780 91156 116786 91158
rect 115841 91155 115907 91156
rect 117221 91155 117287 91158
rect 118182 91156 118188 91220
rect 118252 91218 118258 91220
rect 118601 91218 118667 91221
rect 118252 91216 118667 91218
rect 118252 91160 118606 91216
rect 118662 91160 118667 91216
rect 118252 91158 118667 91160
rect 118252 91156 118258 91158
rect 118601 91155 118667 91158
rect 120206 91156 120212 91220
rect 120276 91218 120282 91220
rect 121361 91218 121427 91221
rect 120276 91216 121427 91218
rect 120276 91160 121366 91216
rect 121422 91160 121427 91216
rect 120276 91158 121427 91160
rect 120276 91156 120282 91158
rect 121361 91155 121427 91158
rect 123150 91156 123156 91220
rect 123220 91218 123226 91220
rect 123753 91218 123819 91221
rect 123220 91216 123819 91218
rect 123220 91160 123758 91216
rect 123814 91160 123819 91216
rect 123220 91158 123819 91160
rect 123220 91156 123226 91158
rect 123753 91155 123819 91158
rect 124029 91220 124095 91221
rect 124029 91216 124076 91220
rect 124140 91218 124146 91220
rect 124029 91160 124034 91216
rect 124029 91156 124076 91160
rect 124140 91158 124186 91218
rect 124140 91156 124146 91158
rect 124438 91156 124444 91220
rect 124508 91218 124514 91220
rect 125501 91218 125567 91221
rect 124508 91216 125567 91218
rect 124508 91160 125506 91216
rect 125562 91160 125567 91216
rect 124508 91158 125567 91160
rect 124508 91156 124514 91158
rect 124029 91155 124095 91156
rect 125501 91155 125567 91158
rect 125726 91156 125732 91220
rect 125796 91218 125802 91220
rect 126697 91218 126763 91221
rect 125796 91216 126763 91218
rect 125796 91160 126702 91216
rect 126758 91160 126763 91216
rect 125796 91158 126763 91160
rect 125796 91156 125802 91158
rect 126697 91155 126763 91158
rect 129406 91156 129412 91220
rect 129476 91218 129482 91220
rect 129641 91218 129707 91221
rect 130745 91220 130811 91221
rect 130694 91218 130700 91220
rect 129476 91216 129707 91218
rect 129476 91160 129646 91216
rect 129702 91160 129707 91216
rect 129476 91158 129707 91160
rect 130654 91158 130700 91218
rect 130764 91216 130811 91220
rect 130806 91160 130811 91216
rect 129476 91156 129482 91158
rect 129641 91155 129707 91158
rect 130694 91156 130700 91158
rect 130764 91156 130811 91160
rect 136030 91156 136036 91220
rect 136100 91218 136106 91220
rect 136541 91218 136607 91221
rect 136100 91216 136607 91218
rect 136100 91160 136546 91216
rect 136602 91160 136607 91216
rect 136100 91158 136607 91160
rect 136100 91156 136106 91158
rect 130745 91155 130811 91156
rect 136541 91155 136607 91158
rect 152038 91156 152044 91220
rect 152108 91218 152114 91220
rect 152641 91218 152707 91221
rect 152108 91216 152707 91218
rect 152108 91160 152646 91216
rect 152702 91160 152707 91216
rect 152108 91158 152707 91160
rect 152108 91156 152114 91158
rect 152641 91155 152707 91158
rect 67633 91082 67699 91085
rect 214414 91082 214420 91084
rect 67633 91080 214420 91082
rect 67633 91024 67638 91080
rect 67694 91024 214420 91080
rect 67633 91022 214420 91024
rect 67633 91019 67699 91022
rect 214414 91020 214420 91022
rect 214484 91020 214490 91084
rect 65977 90946 66043 90949
rect 172094 90946 172100 90948
rect 65977 90944 172100 90946
rect 65977 90888 65982 90944
rect 66038 90888 172100 90944
rect 65977 90886 172100 90888
rect 65977 90883 66043 90886
rect 172094 90884 172100 90886
rect 172164 90884 172170 90948
rect 122046 90748 122052 90812
rect 122116 90810 122122 90812
rect 168230 90810 168236 90812
rect 122116 90750 168236 90810
rect 122116 90748 122122 90750
rect 168230 90748 168236 90750
rect 168300 90748 168306 90812
rect 115473 89722 115539 89725
rect 166206 89722 166212 89724
rect 115473 89720 166212 89722
rect 115473 89664 115478 89720
rect 115534 89664 166212 89720
rect 115473 89662 166212 89664
rect 115473 89659 115539 89662
rect 166206 89660 166212 89662
rect 166276 89660 166282 89724
rect 67725 88226 67791 88229
rect 214833 88226 214899 88229
rect 67725 88224 214899 88226
rect 67725 88168 67730 88224
rect 67786 88168 214838 88224
rect 214894 88168 214899 88224
rect 67725 88166 214899 88168
rect 67725 88163 67791 88166
rect 214833 88163 214899 88166
rect 126697 86866 126763 86869
rect 173198 86866 173204 86868
rect 126697 86864 173204 86866
rect 126697 86808 126702 86864
rect 126758 86808 173204 86864
rect 126697 86806 173204 86808
rect 126697 86803 126763 86806
rect 173198 86804 173204 86806
rect 173268 86804 173274 86868
rect 582373 86186 582439 86189
rect 583520 86186 584960 86276
rect 582373 86184 584960 86186
rect 582373 86128 582378 86184
rect 582434 86128 584960 86184
rect 582373 86126 584960 86128
rect 582373 86123 582439 86126
rect 583520 86036 584960 86126
rect 130745 85506 130811 85509
rect 173014 85506 173020 85508
rect 130745 85504 173020 85506
rect 130745 85448 130750 85504
rect 130806 85448 173020 85504
rect 130745 85446 173020 85448
rect 130745 85443 130811 85446
rect 173014 85444 173020 85446
rect 173084 85444 173090 85508
rect -960 84690 480 84780
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 99189 82786 99255 82789
rect 169150 82786 169156 82788
rect 99189 82784 169156 82786
rect 99189 82728 99194 82784
rect 99250 82728 169156 82784
rect 99189 82726 169156 82728
rect 99189 82723 99255 82726
rect 169150 82724 169156 82726
rect 169220 82724 169226 82788
rect 101949 81426 102015 81429
rect 168966 81426 168972 81428
rect 101949 81424 168972 81426
rect 101949 81368 101954 81424
rect 102010 81368 168972 81424
rect 101949 81366 168972 81368
rect 101949 81363 102015 81366
rect 168966 81364 168972 81366
rect 169036 81364 169042 81428
rect 113081 81290 113147 81293
rect 170254 81290 170260 81292
rect 113081 81288 170260 81290
rect 113081 81232 113086 81288
rect 113142 81232 170260 81288
rect 113081 81230 170260 81232
rect 113081 81227 113147 81230
rect 170254 81228 170260 81230
rect 170324 81228 170330 81292
rect 582741 72994 582807 72997
rect 583520 72994 584960 73084
rect 582741 72992 584960 72994
rect 582741 72936 582746 72992
rect 582802 72936 584960 72992
rect 582741 72934 584960 72936
rect 582741 72931 582807 72934
rect 583520 72844 584960 72934
rect 70393 72450 70459 72453
rect 258758 72450 258764 72452
rect 70393 72448 258764 72450
rect 70393 72392 70398 72448
rect 70454 72392 258764 72448
rect 70393 72390 258764 72392
rect 70393 72387 70459 72390
rect 258758 72388 258764 72390
rect 258828 72388 258834 72452
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 27613 71090 27679 71093
rect 262990 71090 262996 71092
rect 27613 71088 262996 71090
rect 27613 71032 27618 71088
rect 27674 71032 262996 71088
rect 27613 71030 262996 71032
rect 27613 71027 27679 71030
rect 262990 71028 262996 71030
rect 263060 71028 263066 71092
rect 124213 62794 124279 62797
rect 236494 62794 236500 62796
rect 124213 62792 236500 62794
rect 124213 62736 124218 62792
rect 124274 62736 236500 62792
rect 124213 62734 236500 62736
rect 124213 62731 124279 62734
rect 236494 62732 236500 62734
rect 236564 62732 236570 62796
rect 583520 59666 584960 59756
rect 567150 59606 584960 59666
rect 298686 59332 298692 59396
rect 298756 59394 298762 59396
rect 567150 59394 567210 59606
rect 583520 59516 584960 59606
rect 298756 59334 567210 59394
rect 298756 59332 298762 59334
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 40033 57218 40099 57221
rect 253054 57218 253060 57220
rect 40033 57216 253060 57218
rect 40033 57160 40038 57216
rect 40094 57160 253060 57216
rect 40033 57158 253060 57160
rect 40033 57155 40099 57158
rect 253054 57156 253060 57158
rect 253124 57156 253130 57220
rect 2773 55858 2839 55861
rect 253238 55858 253244 55860
rect 2773 55856 253244 55858
rect 2773 55800 2778 55856
rect 2834 55800 253244 55856
rect 2773 55798 253244 55800
rect 2773 55795 2839 55798
rect 253238 55796 253244 55798
rect 253308 55796 253314 55860
rect 62113 51778 62179 51781
rect 258574 51778 258580 51780
rect 62113 51776 258580 51778
rect 62113 51720 62118 51776
rect 62174 51720 258580 51776
rect 62113 51718 258580 51720
rect 62113 51715 62179 51718
rect 258574 51716 258580 51718
rect 258644 51716 258650 51780
rect 77293 47562 77359 47565
rect 264278 47562 264284 47564
rect 77293 47560 264284 47562
rect 77293 47504 77298 47560
rect 77354 47504 264284 47560
rect 77293 47502 264284 47504
rect 77293 47499 77359 47502
rect 264278 47500 264284 47502
rect 264348 47500 264354 47564
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 42793 46202 42859 46205
rect 260046 46202 260052 46204
rect 42793 46200 260052 46202
rect 42793 46144 42798 46200
rect 42854 46144 260052 46200
rect 42793 46142 260052 46144
rect 42793 46139 42859 46142
rect 260046 46140 260052 46142
rect 260116 46140 260122 46204
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2865 45522 2931 45525
rect -960 45520 2931 45522
rect -960 45464 2870 45520
rect 2926 45464 2931 45520
rect -960 45462 2931 45464
rect -960 45372 480 45462
rect 2865 45459 2931 45462
rect 1393 44842 1459 44845
rect 227662 44842 227668 44844
rect 1393 44840 227668 44842
rect 1393 44784 1398 44840
rect 1454 44784 227668 44840
rect 1393 44782 227668 44784
rect 1393 44779 1459 44782
rect 227662 44780 227668 44782
rect 227732 44780 227738 44844
rect 31753 43482 31819 43485
rect 262806 43482 262812 43484
rect 31753 43480 262812 43482
rect 31753 43424 31758 43480
rect 31814 43424 262812 43480
rect 31753 43422 262812 43424
rect 31753 43419 31819 43422
rect 262806 43420 262812 43422
rect 262876 43420 262882 43484
rect 27705 40626 27771 40629
rect 255814 40626 255820 40628
rect 27705 40624 255820 40626
rect 27705 40568 27710 40624
rect 27766 40568 255820 40624
rect 27705 40566 255820 40568
rect 27705 40563 27771 40566
rect 255814 40564 255820 40566
rect 255884 40564 255890 40628
rect 19425 36546 19491 36549
rect 264094 36546 264100 36548
rect 19425 36544 264100 36546
rect 19425 36488 19430 36544
rect 19486 36488 264100 36544
rect 19425 36486 264100 36488
rect 19425 36483 19491 36486
rect 264094 36484 264100 36486
rect 264164 36484 264170 36548
rect 37273 33826 37339 33829
rect 260230 33826 260236 33828
rect 37273 33824 260236 33826
rect 37273 33768 37278 33824
rect 37334 33768 260236 33824
rect 37273 33766 260236 33768
rect 37273 33763 37339 33766
rect 260230 33764 260236 33766
rect 260300 33764 260306 33828
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 44173 22674 44239 22677
rect 262070 22674 262076 22676
rect 44173 22672 262076 22674
rect 44173 22616 44178 22672
rect 44234 22616 262076 22672
rect 44173 22614 262076 22616
rect 44173 22611 44239 22614
rect 262070 22612 262076 22614
rect 262140 22612 262146 22676
rect 582649 19818 582715 19821
rect 583520 19818 584960 19908
rect 582649 19816 584960 19818
rect 582649 19760 582654 19816
rect 582710 19760 584960 19816
rect 582649 19758 584960 19760
rect 582649 19755 582715 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 45553 17234 45619 17237
rect 250294 17234 250300 17236
rect 45553 17232 250300 17234
rect 45553 17176 45558 17232
rect 45614 17176 250300 17232
rect 45553 17174 250300 17176
rect 45553 17171 45619 17174
rect 250294 17172 250300 17174
rect 250364 17172 250370 17236
rect 7649 11658 7715 11661
rect 266854 11658 266860 11660
rect 7649 11656 266860 11658
rect 7649 11600 7654 11656
rect 7710 11600 266860 11656
rect 7649 11598 266860 11600
rect 7649 11595 7715 11598
rect 266854 11596 266860 11598
rect 266924 11596 266930 11660
rect 103329 10434 103395 10437
rect 232446 10434 232452 10436
rect 103329 10432 232452 10434
rect 103329 10376 103334 10432
rect 103390 10376 232452 10432
rect 103329 10374 232452 10376
rect 103329 10371 103395 10374
rect 232446 10372 232452 10374
rect 232516 10372 232522 10436
rect 2865 10298 2931 10301
rect 251766 10298 251772 10300
rect 2865 10296 251772 10298
rect 2865 10240 2870 10296
rect 2926 10240 251772 10296
rect 2865 10238 251772 10240
rect 2865 10235 2931 10238
rect 251766 10236 251772 10238
rect 251836 10236 251842 10300
rect 34789 7578 34855 7581
rect 249006 7578 249012 7580
rect 34789 7576 249012 7578
rect 34789 7520 34794 7576
rect 34850 7520 249012 7576
rect 34789 7518 249012 7520
rect 34789 7515 34855 7518
rect 249006 7516 249012 7518
rect 249076 7516 249082 7580
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 6453 4858 6519 4861
rect 265750 4858 265756 4860
rect 6453 4856 265756 4858
rect 6453 4800 6458 4856
rect 6514 4800 265756 4856
rect 6453 4798 265756 4800
rect 6453 4795 6519 4798
rect 265750 4796 265756 4798
rect 265820 4796 265826 4860
<< via3 >>
rect 191604 697444 191668 697508
rect 255820 576812 255884 576876
rect 187556 456860 187620 456924
rect 190500 397428 190564 397492
rect 291148 299508 291212 299572
rect 295564 298148 295628 298212
rect 258396 296924 258460 296988
rect 295380 296788 295444 296852
rect 249012 294204 249076 294268
rect 288388 294068 288452 294132
rect 200252 293932 200316 293996
rect 288572 292572 288636 292636
rect 200068 291544 200132 291548
rect 200068 291488 200118 291544
rect 200118 291488 200132 291544
rect 200068 291484 200132 291488
rect 200068 290668 200132 290732
rect 195836 289852 195900 289916
rect 253060 285092 253124 285156
rect 195652 283732 195716 283796
rect 250300 281692 250364 281756
rect 278820 278972 278884 279036
rect 251220 274892 251284 274956
rect 199884 273804 199948 273868
rect 249748 269180 249812 269244
rect 249564 268364 249628 268428
rect 197124 252316 197188 252380
rect 252508 246332 252572 246396
rect 200620 245924 200684 245988
rect 191604 242932 191668 242996
rect 192340 242116 192404 242180
rect 187556 241572 187620 241636
rect 190500 240136 190564 240140
rect 190500 240080 190550 240136
rect 190550 240080 190564 240136
rect 190500 240076 190564 240080
rect 236500 239668 236564 239732
rect 238524 239668 238588 239732
rect 237420 239532 237484 239596
rect 241652 239396 241716 239460
rect 255820 238580 255884 238644
rect 192340 238444 192404 238508
rect 200620 236540 200684 236604
rect 244780 235180 244844 235244
rect 298692 228244 298756 228308
rect 287100 197916 287164 197980
rect 285628 193836 285692 193900
rect 290596 191116 290660 191180
rect 294276 190980 294340 191044
rect 233372 186900 233436 186964
rect 276612 185540 276676 185604
rect 287284 184180 287348 184244
rect 228772 181460 228836 181524
rect 284340 181460 284404 181524
rect 292620 181324 292684 181388
rect 241652 180100 241716 180164
rect 166212 179420 166276 179484
rect 234660 178740 234724 178804
rect 105676 177652 105740 177716
rect 108068 177712 108132 177716
rect 108068 177656 108118 177712
rect 108118 177656 108132 177712
rect 108068 177652 108132 177656
rect 114324 177652 114388 177716
rect 119476 177712 119540 177716
rect 119476 177656 119526 177712
rect 119526 177656 119540 177712
rect 119476 177652 119540 177656
rect 124444 177652 124508 177716
rect 127020 177712 127084 177716
rect 127020 177656 127070 177712
rect 127070 177656 127084 177712
rect 127020 177652 127084 177656
rect 130700 177712 130764 177716
rect 130700 177656 130750 177712
rect 130750 177656 130764 177712
rect 130700 177652 130764 177656
rect 132356 177712 132420 177716
rect 132356 177656 132406 177712
rect 132406 177656 132420 177712
rect 132356 177652 132420 177656
rect 276612 177516 276676 177580
rect 233188 177380 233252 177444
rect 291332 177380 291396 177444
rect 237604 177244 237668 177308
rect 253060 177244 253124 177308
rect 113220 177108 113284 177172
rect 123156 177108 123220 177172
rect 129412 177168 129476 177172
rect 129412 177112 129462 177168
rect 129462 177112 129476 177168
rect 129412 177108 129476 177112
rect 97028 176972 97092 177036
rect 98316 176972 98380 177036
rect 101996 176972 102060 177036
rect 100708 176836 100772 176900
rect 166396 176836 166460 176900
rect 104572 176760 104636 176764
rect 104572 176704 104622 176760
rect 104622 176704 104636 176760
rect 104572 176700 104636 176704
rect 106964 176760 107028 176764
rect 106964 176704 107014 176760
rect 107014 176704 107028 176760
rect 106964 176700 107028 176704
rect 109540 176760 109604 176764
rect 109540 176704 109590 176760
rect 109590 176704 109604 176760
rect 109540 176700 109604 176704
rect 110644 176760 110708 176764
rect 110644 176704 110694 176760
rect 110694 176704 110708 176760
rect 110644 176700 110708 176704
rect 112116 176700 112180 176764
rect 118372 176760 118436 176764
rect 118372 176704 118422 176760
rect 118422 176704 118436 176760
rect 118372 176700 118436 176704
rect 125732 176700 125796 176764
rect 133092 176760 133156 176764
rect 133092 176704 133142 176760
rect 133142 176704 133156 176760
rect 133092 176700 133156 176704
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 158852 176700 158916 176764
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 128124 176428 128188 176492
rect 240364 175884 240428 175948
rect 281580 175884 281644 175948
rect 116900 175400 116964 175404
rect 116900 175344 116950 175400
rect 116950 175344 116964 175400
rect 116900 175340 116964 175344
rect 120764 175400 120828 175404
rect 120764 175344 120814 175400
rect 120814 175344 120828 175400
rect 120764 175340 120828 175344
rect 121868 175400 121932 175404
rect 121868 175344 121918 175400
rect 121918 175344 121932 175400
rect 121868 175340 121932 175344
rect 134380 175400 134444 175404
rect 134380 175344 134430 175400
rect 134430 175344 134444 175400
rect 134380 175340 134444 175344
rect 115726 174992 115790 174996
rect 115726 174936 115754 174992
rect 115754 174936 115790 174992
rect 279372 175068 279436 175132
rect 115726 174932 115790 174936
rect 229140 174252 229204 174316
rect 214420 173164 214484 173228
rect 295564 171124 295628 171188
rect 296668 171184 296732 171188
rect 296668 171128 296682 171184
rect 296682 171128 296732 171184
rect 296668 171124 296732 171128
rect 268516 168540 268580 168604
rect 268516 168132 268580 168196
rect 268516 167180 268580 167244
rect 268516 166772 268580 166836
rect 236500 163780 236564 163844
rect 234660 163372 234724 163436
rect 268516 161604 268580 161668
rect 214420 160788 214484 160852
rect 250300 159972 250364 160036
rect 166396 156028 166460 156092
rect 268516 157252 268580 157316
rect 281580 156980 281644 157044
rect 166212 154532 166276 154596
rect 251220 155212 251284 155276
rect 237420 153852 237484 153916
rect 232452 153172 232516 153236
rect 252508 150996 252572 151060
rect 233372 148684 233436 148748
rect 268516 147868 268580 147932
rect 268516 146100 268580 146164
rect 249748 145556 249812 145620
rect 173020 145012 173084 145076
rect 241836 144876 241900 144940
rect 230980 144060 231044 144124
rect 285628 143108 285692 143172
rect 173204 142156 173268 142220
rect 268516 142292 268580 142356
rect 258396 142020 258460 142084
rect 268516 141884 268580 141948
rect 237604 141612 237668 141676
rect 233740 141068 233804 141132
rect 267780 141068 267844 141132
rect 268332 140932 268396 140996
rect 291332 140796 291396 140860
rect 168236 139436 168300 139500
rect 236500 139844 236564 139908
rect 244780 139708 244844 139772
rect 251772 139708 251836 139772
rect 232452 139164 232516 139228
rect 233188 138756 233252 138820
rect 241652 138212 241716 138276
rect 238524 137804 238588 137868
rect 166212 136716 166276 136780
rect 232452 137124 232516 137188
rect 240364 136308 240428 136372
rect 170260 135220 170324 135284
rect 296484 135220 296548 135284
rect 290596 134132 290660 134196
rect 258764 133180 258828 133244
rect 288572 131140 288636 131204
rect 250300 130188 250364 130252
rect 260052 129780 260116 129844
rect 168972 128420 169036 128484
rect 287284 128692 287348 128756
rect 255820 128420 255884 128484
rect 268516 128556 268580 128620
rect 262812 128148 262876 128212
rect 268516 128148 268580 128212
rect 169156 127060 169220 127124
rect 268516 127196 268580 127260
rect 287100 127060 287164 127124
rect 264100 126788 264164 126852
rect 268516 126788 268580 126852
rect 230980 125428 231044 125492
rect 268516 121620 268580 121684
rect 294276 121484 294340 121548
rect 264284 120396 264348 120460
rect 268516 119852 268580 119916
rect 258580 118764 258644 118828
rect 260236 116044 260300 116108
rect 267780 115908 267844 115972
rect 268332 116044 268396 116108
rect 249012 114820 249076 114884
rect 262996 114684 263060 114748
rect 292620 113188 292684 113252
rect 291148 109516 291212 109580
rect 295380 109108 295444 109172
rect 170444 108292 170508 108356
rect 268332 107884 268396 107948
rect 268332 107476 268396 107540
rect 288388 104892 288452 104956
rect 284340 103940 284404 104004
rect 214420 103532 214484 103596
rect 262076 102716 262140 102780
rect 268332 102716 268396 102780
rect 172100 102308 172164 102372
rect 253060 102444 253124 102508
rect 267780 102444 267844 102508
rect 266860 98772 266924 98836
rect 233740 97956 233804 98020
rect 229140 97004 229204 97068
rect 253244 96596 253308 96660
rect 265756 96596 265820 96660
rect 267780 96596 267844 96660
rect 268332 96732 268396 96796
rect 166948 95780 167012 95844
rect 227668 95236 227732 95300
rect 228956 95236 229020 95300
rect 195836 95100 195900 95164
rect 105662 94692 105726 94756
rect 112326 94752 112390 94756
rect 112326 94696 112350 94752
rect 112350 94696 112390 94752
rect 112326 94692 112390 94696
rect 128102 94752 128166 94756
rect 128102 94696 128138 94752
rect 128138 94696 128166 94752
rect 128102 94692 128166 94696
rect 151766 94752 151830 94756
rect 151766 94696 151782 94752
rect 151782 94696 151830 94752
rect 151766 94692 151830 94696
rect 106412 94072 106476 94076
rect 106412 94016 106462 94072
rect 106462 94016 106476 94072
rect 106412 94012 106476 94016
rect 121684 93664 121748 93668
rect 121684 93608 121734 93664
rect 121734 93608 121748 93664
rect 121684 93604 121748 93608
rect 88932 93528 88996 93532
rect 88932 93472 88982 93528
rect 88982 93472 88996 93528
rect 88932 93468 88996 93472
rect 111196 93528 111260 93532
rect 111196 93472 111246 93528
rect 111246 93472 111260 93528
rect 111196 93468 111260 93472
rect 119292 93468 119356 93532
rect 195652 93604 195716 93668
rect 134380 93528 134444 93532
rect 134380 93472 134430 93528
rect 134430 93472 134444 93528
rect 134380 93468 134444 93472
rect 197124 93468 197188 93532
rect 103284 93196 103348 93260
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 85804 92380 85868 92444
rect 98500 92440 98564 92444
rect 98500 92384 98550 92440
rect 98550 92384 98564 92440
rect 98500 92380 98564 92384
rect 104204 92380 104268 92444
rect 104572 92440 104636 92444
rect 104572 92384 104622 92440
rect 104622 92384 104636 92440
rect 104572 92380 104636 92384
rect 106596 92440 106660 92444
rect 106596 92384 106646 92440
rect 106646 92384 106660 92440
rect 106596 92380 106660 92384
rect 110644 92440 110708 92444
rect 110644 92384 110694 92440
rect 110694 92384 110708 92440
rect 110644 92380 110708 92384
rect 118004 92440 118068 92444
rect 118004 92384 118054 92440
rect 118054 92384 118068 92440
rect 118004 92380 118068 92384
rect 126652 92440 126716 92444
rect 126652 92384 126702 92440
rect 126702 92384 126716 92440
rect 126652 92380 126716 92384
rect 133092 92440 133156 92444
rect 133092 92384 133142 92440
rect 133142 92384 133156 92440
rect 133092 92380 133156 92384
rect 151492 92440 151556 92444
rect 151492 92384 151542 92440
rect 151542 92384 151556 92440
rect 151492 92380 151556 92384
rect 113036 92244 113100 92308
rect 170444 92244 170508 92308
rect 88012 92108 88076 92172
rect 166948 92108 167012 92172
rect 115428 92032 115492 92036
rect 115428 91976 115478 92032
rect 115478 91976 115492 92032
rect 115428 91972 115492 91976
rect 126468 92032 126532 92036
rect 126468 91976 126518 92032
rect 126518 91976 126532 92032
rect 126468 91972 126532 91976
rect 151308 92032 151372 92036
rect 151308 91976 151358 92032
rect 151358 91976 151372 92032
rect 151308 91972 151372 91976
rect 90220 91700 90284 91764
rect 119660 91700 119724 91764
rect 105492 91564 105556 91628
rect 132356 91624 132420 91628
rect 132356 91568 132406 91624
rect 132406 91568 132420 91624
rect 132356 91564 132420 91568
rect 101812 91488 101876 91492
rect 101812 91432 101862 91488
rect 101862 91432 101876 91488
rect 101812 91428 101876 91432
rect 109172 91428 109236 91492
rect 122788 91428 122852 91492
rect 93900 91292 93964 91356
rect 98132 91292 98196 91356
rect 100524 91352 100588 91356
rect 100524 91296 100574 91352
rect 100574 91296 100588 91352
rect 100524 91292 100588 91296
rect 100892 91292 100956 91356
rect 107700 91292 107764 91356
rect 114324 91352 114388 91356
rect 114324 91296 114374 91352
rect 114374 91296 114388 91352
rect 114324 91292 114388 91296
rect 117084 91352 117148 91356
rect 117084 91296 117134 91352
rect 117134 91296 117148 91352
rect 117084 91292 117148 91296
rect 120580 91292 120644 91356
rect 125364 91352 125428 91356
rect 125364 91296 125414 91352
rect 125414 91296 125428 91352
rect 125364 91292 125428 91296
rect 74764 91156 74828 91220
rect 84332 91156 84396 91220
rect 86724 91156 86788 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 95004 91156 95068 91220
rect 96292 91156 96356 91220
rect 96660 91156 96724 91220
rect 97212 91156 97276 91220
rect 99052 91156 99116 91220
rect 99972 91156 100036 91220
rect 101996 91216 102060 91220
rect 101996 91160 102046 91216
rect 102046 91160 102060 91216
rect 101996 91156 102060 91160
rect 102732 91156 102796 91220
rect 108068 91156 108132 91220
rect 109540 91156 109604 91220
rect 111932 91156 111996 91220
rect 113220 91156 113284 91220
rect 114876 91156 114940 91220
rect 115796 91216 115860 91220
rect 115796 91160 115846 91216
rect 115846 91160 115860 91216
rect 115796 91156 115860 91160
rect 116716 91156 116780 91220
rect 118188 91156 118252 91220
rect 120212 91156 120276 91220
rect 123156 91156 123220 91220
rect 124076 91216 124140 91220
rect 124076 91160 124090 91216
rect 124090 91160 124140 91216
rect 124076 91156 124140 91160
rect 124444 91156 124508 91220
rect 125732 91156 125796 91220
rect 129412 91156 129476 91220
rect 130700 91216 130764 91220
rect 130700 91160 130750 91216
rect 130750 91160 130764 91216
rect 130700 91156 130764 91160
rect 136036 91156 136100 91220
rect 152044 91156 152108 91220
rect 214420 91020 214484 91084
rect 172100 90884 172164 90948
rect 122052 90748 122116 90812
rect 168236 90748 168300 90812
rect 166212 89660 166276 89724
rect 173204 86804 173268 86868
rect 173020 85444 173084 85508
rect 169156 82724 169220 82788
rect 168972 81364 169036 81428
rect 170260 81228 170324 81292
rect 258764 72388 258828 72452
rect 262996 71028 263060 71092
rect 236500 62732 236564 62796
rect 298692 59332 298756 59396
rect 253060 57156 253124 57220
rect 253244 55796 253308 55860
rect 258580 51716 258644 51780
rect 264284 47500 264348 47564
rect 260052 46140 260116 46204
rect 227668 44780 227732 44844
rect 262812 43420 262876 43484
rect 255820 40564 255884 40628
rect 264100 36484 264164 36548
rect 260236 33764 260300 33828
rect 262076 22612 262140 22676
rect 250300 17172 250364 17236
rect 266860 11596 266924 11660
rect 232452 10372 232516 10436
rect 251772 10236 251836 10300
rect 249012 7516 249076 7580
rect 265756 4796 265820 4860
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176600 67574 212058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 177036 97093 177037
rect 97027 176972 97028 177036
rect 97092 176972 97093 177036
rect 97027 176971 97093 176972
rect 98315 177036 98381 177037
rect 98315 176972 98316 177036
rect 98380 176972 98381 177036
rect 98315 176971 98381 176972
rect 97030 175130 97090 176971
rect 96960 175070 97090 175130
rect 98318 175130 98378 176971
rect 99234 176600 99854 208338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 101995 177036 102061 177037
rect 101995 176972 101996 177036
rect 102060 176972 102061 177036
rect 101995 176971 102061 176972
rect 100707 176900 100773 176901
rect 100707 176836 100708 176900
rect 100772 176836 100773 176900
rect 100707 176835 100773 176836
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 176835
rect 101998 175130 102058 176971
rect 102954 176600 103574 212058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 105675 177716 105741 177717
rect 105675 177652 105676 177716
rect 105740 177652 105741 177716
rect 105675 177651 105741 177652
rect 108067 177716 108133 177717
rect 108067 177652 108068 177716
rect 108132 177652 108133 177716
rect 108067 177651 108133 177652
rect 104571 176764 104637 176765
rect 104571 176700 104572 176764
rect 104636 176700 104637 176764
rect 104571 176699 104637 176700
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 176699
rect 105678 175130 105738 177651
rect 106963 176764 107029 176765
rect 106963 176700 106964 176764
rect 107028 176700 107029 176764
rect 106963 176699 107029 176700
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 176699
rect 108070 175130 108130 177651
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 109542 175130 109602 176699
rect 109794 176600 110414 182898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113219 177172 113285 177173
rect 113219 177108 113220 177172
rect 113284 177108 113285 177172
rect 113219 177107 113285 177108
rect 110643 176764 110709 176765
rect 110643 176700 110644 176764
rect 110708 176700 110709 176764
rect 110643 176699 110709 176700
rect 112115 176764 112181 176765
rect 112115 176700 112116 176764
rect 112180 176700 112181 176764
rect 112115 176699 112181 176700
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 176699
rect 112118 175130 112178 176699
rect 113222 175130 113282 177107
rect 113514 176600 114134 186618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 114323 177716 114389 177717
rect 114323 177652 114324 177716
rect 114388 177652 114389 177716
rect 114323 177651 114389 177652
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 177651
rect 117234 176600 117854 190338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 119475 177716 119541 177717
rect 119475 177652 119476 177716
rect 119540 177652 119541 177716
rect 119475 177651 119541 177652
rect 118371 176764 118437 176765
rect 118371 176700 118372 176764
rect 118436 176700 118437 176764
rect 118371 176699 118437 176700
rect 116899 175404 116965 175405
rect 116899 175340 116900 175404
rect 116964 175340 116965 175404
rect 116899 175339 116965 175340
rect 116902 175130 116962 175339
rect 118374 175130 118434 176699
rect 119478 175130 119538 177651
rect 120954 176600 121574 194058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 124443 177716 124509 177717
rect 124443 177652 124444 177716
rect 124508 177652 124509 177716
rect 124443 177651 124509 177652
rect 127019 177716 127085 177717
rect 127019 177652 127020 177716
rect 127084 177652 127085 177716
rect 127019 177651 127085 177652
rect 123155 177172 123221 177173
rect 123155 177108 123156 177172
rect 123220 177108 123221 177172
rect 123155 177107 123221 177108
rect 120763 175404 120829 175405
rect 120763 175340 120764 175404
rect 120828 175340 120829 175404
rect 120763 175339 120829 175340
rect 121867 175404 121933 175405
rect 121867 175340 121868 175404
rect 121932 175340 121933 175404
rect 121867 175339 121933 175340
rect 120766 175130 120826 175339
rect 121870 175130 121930 175339
rect 123158 175130 123218 177107
rect 124446 175130 124506 177651
rect 125731 176764 125797 176765
rect 125731 176700 125732 176764
rect 125796 176700 125797 176764
rect 125731 176699 125797 176700
rect 125734 175130 125794 176699
rect 127022 175130 127082 177651
rect 127794 176600 128414 200898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 130699 177716 130765 177717
rect 130699 177652 130700 177716
rect 130764 177652 130765 177716
rect 130699 177651 130765 177652
rect 129411 177172 129477 177173
rect 129411 177108 129412 177172
rect 129476 177108 129477 177172
rect 129411 177107 129477 177108
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 114326 175070 114428 175130
rect 116902 175070 117012 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115725 174996 115791 174997
rect 115725 174932 115726 174996
rect 115790 174932 115791 174996
rect 115725 174931 115791 174932
rect 115728 174494 115788 174931
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 177107
rect 130702 175130 130762 177651
rect 131514 176600 132134 204618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 132355 177716 132421 177717
rect 132355 177652 132356 177716
rect 132420 177652 132421 177716
rect 132355 177651 132421 177652
rect 132358 175130 132418 177651
rect 133091 176764 133157 176765
rect 133091 176700 133092 176764
rect 133156 176700 133157 176764
rect 133091 176699 133157 176700
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 176699
rect 135234 176600 135854 208338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 134379 175404 134445 175405
rect 134379 175340 134380 175404
rect 134444 175340 134445 175404
rect 134379 175339 134445 175340
rect 134382 175130 134442 175339
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135720 175070 136098 175130
rect 148182 175130 148242 176699
rect 149514 176600 150134 186618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 163794 176600 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 166211 179484 166277 179485
rect 166211 179420 166212 179484
rect 166276 179420 166277 179484
rect 166211 179419 166277 179420
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 166214 154597 166274 179419
rect 166395 176900 166461 176901
rect 166395 176836 166396 176900
rect 166460 176836 166461 176900
rect 166395 176835 166461 176836
rect 166398 156093 166458 176835
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 166395 156092 166461 156093
rect 166395 156028 166396 156092
rect 166460 156028 166461 156092
rect 166395 156027 166461 156028
rect 166211 154596 166277 154597
rect 166211 154532 166212 154596
rect 166276 154532 166277 154596
rect 166211 154531 166277 154532
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 166211 136780 166277 136781
rect 166211 136716 166212 136780
rect 166276 136716 166277 136780
rect 166211 136715 166277 136716
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85866 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 91221 84394 94830
rect 84331 91220 84397 91221
rect 84331 91156 84332 91220
rect 84396 91156 84397 91220
rect 84331 91155 84397 91156
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 85806 92445 85866 94830
rect 85803 92444 85869 92445
rect 85803 92380 85804 92444
rect 85868 92380 85869 92444
rect 85803 92379 85869 92380
rect 86726 91221 86786 94830
rect 88014 92173 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 93533 88994 94830
rect 88931 93532 88997 93533
rect 88931 93468 88932 93532
rect 88996 93468 88997 93532
rect 88931 93467 88997 93468
rect 88011 92172 88077 92173
rect 88011 92108 88012 92172
rect 88076 92108 88077 92172
rect 88011 92107 88077 92108
rect 90222 91765 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 90219 91764 90285 91765
rect 90219 91700 90220 91764
rect 90284 91700 90285 91764
rect 90219 91699 90285 91700
rect 91326 91221 91386 94830
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91357 93962 94830
rect 93899 91356 93965 91357
rect 93899 91292 93900 91356
rect 93964 91292 93965 91356
rect 93899 91291 93965 91292
rect 95006 91221 95066 94830
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91221 96722 94830
rect 97214 91221 97274 94830
rect 98134 91357 98194 94830
rect 98502 92445 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 99544 94830 100034 94890
rect 98499 92444 98565 92445
rect 98499 92380 98500 92444
rect 98564 92380 98565 92444
rect 98499 92379 98565 92380
rect 98131 91356 98197 91357
rect 98131 91292 98132 91356
rect 98196 91292 98197 91356
rect 98131 91291 98197 91292
rect 99054 91221 99114 94830
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 96659 91220 96725 91221
rect 96659 91156 96660 91220
rect 96724 91156 96725 91220
rect 96659 91155 96725 91156
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 99051 91220 99117 91221
rect 99051 91156 99052 91220
rect 99116 91156 99117 91220
rect 99051 91155 99117 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 91221 100034 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 100526 91357 100586 94830
rect 100894 91357 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 101814 91493 101874 94830
rect 101811 91492 101877 91493
rect 101811 91428 101812 91492
rect 101876 91428 101877 91492
rect 101811 91427 101877 91428
rect 100523 91356 100589 91357
rect 100523 91292 100524 91356
rect 100588 91292 100589 91356
rect 100523 91291 100589 91292
rect 100891 91356 100957 91357
rect 100891 91292 100892 91356
rect 100956 91292 100957 91356
rect 100891 91291 100957 91292
rect 101998 91221 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 102918 93870 102978 94830
rect 102734 93810 102978 93870
rect 102734 91221 102794 93810
rect 103286 93261 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 103283 93260 103349 93261
rect 103283 93196 103284 93260
rect 103348 93196 103349 93260
rect 103283 93195 103349 93196
rect 99971 91220 100037 91221
rect 99971 91156 99972 91220
rect 100036 91156 100037 91220
rect 99971 91155 100037 91156
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 102731 91220 102797 91221
rect 102731 91156 102732 91220
rect 102796 91156 102797 91220
rect 102731 91155 102797 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 92445 104266 94830
rect 104574 92445 104634 94830
rect 104203 92444 104269 92445
rect 104203 92380 104204 92444
rect 104268 92380 104269 92444
rect 104203 92379 104269 92380
rect 104571 92444 104637 92445
rect 104571 92380 104572 92444
rect 104636 92380 104637 92444
rect 104571 92379 104637 92380
rect 105494 91629 105554 94830
rect 105664 94757 105724 95200
rect 106480 94890 106540 95200
rect 106414 94830 106540 94890
rect 105661 94756 105727 94757
rect 105661 94692 105662 94756
rect 105726 94692 105727 94756
rect 105661 94691 105727 94692
rect 106414 94077 106474 94830
rect 106616 94210 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106598 94150 106676 94210
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 106411 94076 106477 94077
rect 106411 94012 106412 94076
rect 106476 94012 106477 94076
rect 106411 94011 106477 94012
rect 106598 92445 106658 94150
rect 106595 92444 106661 92445
rect 106595 92380 106596 92444
rect 106660 92380 106661 92444
rect 106595 92379 106661 92380
rect 105491 91628 105557 91629
rect 105491 91564 105492 91628
rect 105556 91564 105557 91628
rect 105491 91563 105557 91564
rect 107702 91357 107762 94830
rect 107699 91356 107765 91357
rect 107699 91292 107700 91356
rect 107764 91292 107765 91356
rect 107699 91291 107765 91292
rect 108070 91221 108130 94830
rect 109174 91493 109234 94830
rect 109171 91492 109237 91493
rect 109171 91428 109172 91492
rect 109236 91428 109237 91492
rect 109171 91427 109237 91428
rect 109542 91221 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 111920 94830 111994 94890
rect 110094 93261 110154 94830
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 92445 110706 94830
rect 111198 93533 111258 94830
rect 111195 93532 111261 93533
rect 111195 93468 111196 93532
rect 111260 93468 111261 93532
rect 111195 93467 111261 93468
rect 110643 92444 110709 92445
rect 110643 92380 110644 92444
rect 110708 92380 110709 92444
rect 110643 92379 110709 92380
rect 111934 91221 111994 94830
rect 112328 94757 112388 95200
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 113038 94830 113204 94890
rect 113406 94830 113748 94890
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 112325 94756 112391 94757
rect 112325 94692 112326 94756
rect 112390 94692 112391 94756
rect 112325 94691 112391 94692
rect 113038 92309 113098 94830
rect 113406 93870 113466 94830
rect 113222 93810 113466 93870
rect 113035 92308 113101 92309
rect 113035 92244 113036 92308
rect 113100 92244 113101 92308
rect 113035 92243 113101 92244
rect 113222 91221 113282 93810
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 113219 91220 113285 91221
rect 113219 91156 113220 91220
rect 113284 91156 113285 91220
rect 113219 91155 113285 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91357 114386 94830
rect 114323 91356 114389 91357
rect 114323 91292 114324 91356
rect 114388 91292 114389 91356
rect 114323 91291 114389 91292
rect 114878 91221 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115430 92037 115490 94830
rect 115427 92036 115493 92037
rect 115427 91972 115428 92036
rect 115492 91972 115493 92036
rect 115427 91971 115493 91972
rect 115798 91221 115858 94830
rect 116718 91221 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 117086 91357 117146 94830
rect 117083 91356 117149 91357
rect 117083 91292 117084 91356
rect 117148 91292 117149 91356
rect 117083 91291 117149 91292
rect 114875 91220 114941 91221
rect 114875 91156 114876 91220
rect 114940 91156 114941 91220
rect 114875 91155 114941 91156
rect 115795 91220 115861 91221
rect 115795 91156 115796 91220
rect 115860 91156 115861 91220
rect 115795 91155 115861 91156
rect 116715 91220 116781 91221
rect 116715 91156 116716 91220
rect 116780 91156 116781 91220
rect 116715 91155 116781 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 92445 118066 94830
rect 118003 92444 118069 92445
rect 118003 92380 118004 92444
rect 118068 92380 118069 92444
rect 118003 92379 118069 92380
rect 118190 91221 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 119294 93533 119354 94830
rect 119291 93532 119357 93533
rect 119291 93468 119292 93532
rect 119356 93468 119357 93532
rect 119291 93467 119357 93468
rect 119662 91765 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 119659 91764 119725 91765
rect 119659 91700 119660 91764
rect 119724 91700 119725 91764
rect 119659 91699 119725 91700
rect 120214 91221 120274 94830
rect 120582 91357 120642 94830
rect 121686 93669 121746 94830
rect 121683 93668 121749 93669
rect 121683 93604 121684 93668
rect 121748 93604 121749 93668
rect 121683 93603 121749 93604
rect 120579 91356 120645 91357
rect 120579 91292 120580 91356
rect 120644 91292 120645 91356
rect 120579 91291 120645 91292
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 120211 91220 120277 91221
rect 120211 91156 120212 91220
rect 120276 91156 120277 91220
rect 120211 91155 120277 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 122054 90813 122114 94830
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122606 91490 122666 93810
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 123158 91221 123218 94830
rect 124078 91221 124138 94830
rect 124446 91221 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 125366 91357 125426 94830
rect 125363 91356 125429 91357
rect 125363 91292 125364 91356
rect 125428 91292 125429 91356
rect 125363 91291 125429 91292
rect 125734 91221 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 126608 94830 126714 94890
rect 126470 92037 126530 94830
rect 126654 92445 126714 94830
rect 128104 94757 128164 95200
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 128101 94756 128167 94757
rect 128101 94692 128102 94756
rect 128166 94692 128167 94756
rect 128101 94691 128167 94692
rect 126651 92444 126717 92445
rect 126651 92380 126652 92444
rect 126716 92380 126717 92444
rect 126651 92379 126717 92380
rect 126467 92036 126533 92037
rect 126467 91972 126468 92036
rect 126532 91972 126533 92036
rect 126467 91971 126533 91972
rect 123155 91220 123221 91221
rect 123155 91156 123156 91220
rect 123220 91156 123221 91220
rect 123155 91155 123221 91156
rect 124075 91220 124141 91221
rect 124075 91156 124076 91220
rect 124140 91156 124141 91220
rect 124075 91155 124141 91156
rect 124443 91220 124509 91221
rect 124443 91156 124444 91220
rect 124508 91156 124509 91220
rect 124443 91155 124509 91156
rect 125731 91220 125797 91221
rect 125731 91156 125732 91220
rect 125796 91156 125797 91220
rect 125731 91155 125797 91156
rect 122051 90812 122117 90813
rect 122051 90748 122052 90812
rect 122116 90748 122117 90812
rect 122051 90747 122117 90748
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 129414 91221 129474 94830
rect 130702 91221 130762 94830
rect 129411 91220 129477 91221
rect 129411 91156 129412 91220
rect 129476 91156 129477 91220
rect 129411 91155 129477 91156
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 91629 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 133094 92445 133154 94830
rect 134382 93533 134442 94830
rect 134379 93532 134445 93533
rect 134379 93468 134380 93532
rect 134444 93468 134445 93532
rect 134379 93467 134445 93468
rect 133091 92444 133157 92445
rect 133091 92380 133092 92444
rect 133156 92380 133157 92444
rect 133091 92379 133157 92380
rect 132355 91628 132421 91629
rect 132355 91564 132356 91628
rect 132420 91564 132421 91628
rect 132355 91563 132421 91564
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 91221 136098 94830
rect 151310 94830 151556 94890
rect 136035 91220 136101 91221
rect 136035 91156 136036 91220
rect 136100 91156 136101 91220
rect 136035 91155 136101 91156
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151310 92037 151370 94830
rect 151632 94754 151692 95200
rect 151768 94757 151828 95200
rect 151494 94694 151692 94754
rect 151765 94756 151831 94757
rect 151494 92445 151554 94694
rect 151765 94692 151766 94756
rect 151830 94692 151831 94756
rect 151904 94754 151964 95200
rect 151904 94694 152106 94754
rect 151765 94691 151831 94692
rect 151491 92444 151557 92445
rect 151491 92380 151492 92444
rect 151556 92380 151557 92444
rect 151491 92379 151557 92380
rect 151307 92036 151373 92037
rect 151307 91972 151308 92036
rect 151372 91972 151373 92036
rect 151307 91971 151373 91972
rect 152046 91221 152106 94694
rect 152043 91220 152109 91221
rect 152043 91156 152044 91220
rect 152108 91156 152109 91220
rect 152043 91155 152109 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 89725 166274 136715
rect 167514 133174 168134 168618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 168235 139500 168301 139501
rect 168235 139436 168236 139500
rect 168300 139436 168301 139500
rect 168235 139435 168301 139436
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166947 95844 167013 95845
rect 166947 95780 166948 95844
rect 167012 95780 167013 95844
rect 166947 95779 167013 95780
rect 166950 92173 167010 95779
rect 166947 92172 167013 92173
rect 166947 92108 166948 92172
rect 167012 92108 167013 92172
rect 166947 92107 167013 92108
rect 166211 89724 166277 89725
rect 166211 89660 166212 89724
rect 166276 89660 166277 89724
rect 166211 89659 166277 89660
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 96618
rect 168238 90813 168298 139435
rect 171234 136894 171854 172338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 173019 145076 173085 145077
rect 173019 145012 173020 145076
rect 173084 145012 173085 145076
rect 173019 145011 173085 145012
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 170259 135284 170325 135285
rect 170259 135220 170260 135284
rect 170324 135220 170325 135284
rect 170259 135219 170325 135220
rect 168971 128484 169037 128485
rect 168971 128420 168972 128484
rect 169036 128420 169037 128484
rect 168971 128419 169037 128420
rect 168235 90812 168301 90813
rect 168235 90748 168236 90812
rect 168300 90748 168301 90812
rect 168235 90747 168301 90748
rect 168974 81429 169034 128419
rect 169155 127124 169221 127125
rect 169155 127060 169156 127124
rect 169220 127060 169221 127124
rect 169155 127059 169221 127060
rect 169158 82789 169218 127059
rect 169155 82788 169221 82789
rect 169155 82724 169156 82788
rect 169220 82724 169221 82788
rect 169155 82723 169221 82724
rect 168971 81428 169037 81429
rect 168971 81364 168972 81428
rect 169036 81364 169037 81428
rect 168971 81363 169037 81364
rect 170262 81293 170322 135219
rect 170443 108356 170509 108357
rect 170443 108292 170444 108356
rect 170508 108292 170509 108356
rect 170443 108291 170509 108292
rect 170446 92309 170506 108291
rect 171234 100894 171854 136338
rect 172099 102372 172165 102373
rect 172099 102308 172100 102372
rect 172164 102308 172165 102372
rect 172099 102307 172165 102308
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 170443 92308 170509 92309
rect 170443 92244 170444 92308
rect 170508 92244 170509 92308
rect 170443 92243 170509 92244
rect 170259 81292 170325 81293
rect 170259 81228 170260 81292
rect 170324 81228 170325 81292
rect 170259 81227 170325 81228
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 100338
rect 172102 90949 172162 102307
rect 172099 90948 172165 90949
rect 172099 90884 172100 90948
rect 172164 90884 172165 90948
rect 172099 90883 172165 90884
rect 173022 85509 173082 145011
rect 173203 142220 173269 142221
rect 173203 142156 173204 142220
rect 173268 142156 173269 142220
rect 173203 142155 173269 142156
rect 173206 86869 173266 142155
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 173203 86868 173269 86869
rect 173203 86804 173204 86868
rect 173268 86804 173269 86868
rect 173203 86803 173269 86804
rect 173019 85508 173085 85509
rect 173019 85444 173020 85508
rect 173084 85444 173085 85508
rect 173019 85443 173085 85444
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 189234 694894 189854 708122
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 191603 697508 191669 697509
rect 191603 697444 191604 697508
rect 191668 697444 191669 697508
rect 191603 697443 191669 697444
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 187555 456924 187621 456925
rect 187555 456860 187556 456924
rect 187620 456860 187621 456924
rect 187555 456859 187621 456860
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 187558 241637 187618 456859
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 190499 397492 190565 397493
rect 190499 397428 190500 397492
rect 190564 397428 190565 397492
rect 190499 397427 190565 397428
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 187555 241636 187621 241637
rect 187555 241572 187556 241636
rect 187620 241572 187621 241636
rect 187555 241571 187621 241572
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 226894 189854 262338
rect 190502 240141 190562 397427
rect 191606 242997 191666 697443
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 294182 200414 308898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 294182 204134 312618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 294182 207854 316338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 294182 211574 320058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 294182 218414 326898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 294182 222134 294618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 294182 225854 298338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 294182 229574 302058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 294182 236414 308898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 294182 240134 312618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 294182 243854 316338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 294182 247574 320058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 255819 576876 255885 576877
rect 255819 576812 255820 576876
rect 255884 576812 255885 576876
rect 255819 576811 255885 576812
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 249011 294268 249077 294269
rect 249011 294204 249012 294268
rect 249076 294204 249077 294268
rect 249011 294203 249077 294204
rect 200251 293996 200317 293997
rect 200251 293932 200252 293996
rect 200316 293932 200317 293996
rect 200251 293931 200317 293932
rect 200067 291548 200133 291549
rect 200067 291484 200068 291548
rect 200132 291484 200133 291548
rect 200067 291483 200133 291484
rect 200070 291410 200130 291483
rect 199886 291350 200130 291410
rect 195835 289916 195901 289917
rect 195835 289852 195836 289916
rect 195900 289852 195901 289916
rect 195835 289851 195901 289852
rect 195651 283796 195717 283797
rect 195651 283732 195652 283796
rect 195716 283732 195717 283796
rect 195651 283731 195717 283732
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 191603 242996 191669 242997
rect 191603 242932 191604 242996
rect 191668 242932 191669 242996
rect 191603 242931 191669 242932
rect 192339 242180 192405 242181
rect 192339 242116 192340 242180
rect 192404 242116 192405 242180
rect 192339 242115 192405 242116
rect 190499 240140 190565 240141
rect 190499 240076 190500 240140
rect 190564 240076 190565 240140
rect 190499 240075 190565 240076
rect 192342 238509 192402 242115
rect 192339 238508 192405 238509
rect 192339 238444 192340 238508
rect 192404 238444 192405 238508
rect 192339 238443 192405 238444
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 195654 93669 195714 283731
rect 195838 95165 195898 289851
rect 199886 273869 199946 291350
rect 200067 290732 200133 290733
rect 200067 290668 200068 290732
rect 200132 290730 200133 290732
rect 200254 290730 200314 293931
rect 200132 290670 200314 290730
rect 200132 290668 200133 290670
rect 200067 290667 200133 290668
rect 249014 287070 249074 294203
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 249014 287010 249626 287070
rect 199883 273868 199949 273869
rect 199883 273804 199884 273868
rect 199948 273804 199949 273868
rect 199883 273803 199949 273804
rect 219768 273454 220088 273486
rect 219768 273218 219810 273454
rect 220046 273218 220088 273454
rect 219768 273134 220088 273218
rect 219768 272898 219810 273134
rect 220046 272898 220088 273134
rect 219768 272866 220088 272898
rect 249566 268429 249626 287010
rect 253059 285156 253125 285157
rect 253059 285092 253060 285156
rect 253124 285092 253125 285156
rect 253059 285091 253125 285092
rect 250299 281756 250365 281757
rect 250299 281692 250300 281756
rect 250364 281692 250365 281756
rect 250299 281691 250365 281692
rect 249747 269244 249813 269245
rect 249747 269180 249748 269244
rect 249812 269180 249813 269244
rect 249747 269179 249813 269180
rect 249563 268428 249629 268429
rect 249563 268364 249564 268428
rect 249628 268364 249629 268428
rect 249563 268363 249629 268364
rect 204408 255454 204728 255486
rect 204408 255218 204450 255454
rect 204686 255218 204728 255454
rect 204408 255134 204728 255218
rect 204408 254898 204450 255134
rect 204686 254898 204728 255134
rect 204408 254866 204728 254898
rect 235128 255454 235448 255486
rect 235128 255218 235170 255454
rect 235406 255218 235448 255454
rect 235128 255134 235448 255218
rect 235128 254898 235170 255134
rect 235406 254898 235448 255134
rect 235128 254866 235448 254898
rect 197123 252380 197189 252381
rect 197123 252316 197124 252380
rect 197188 252316 197189 252380
rect 197123 252315 197189 252316
rect 195835 95164 195901 95165
rect 195835 95100 195836 95164
rect 195900 95100 195901 95164
rect 195835 95099 195901 95100
rect 195651 93668 195717 93669
rect 195651 93604 195652 93668
rect 195716 93604 195717 93668
rect 195651 93603 195717 93604
rect 197126 93533 197186 252315
rect 200619 245988 200685 245989
rect 200619 245924 200620 245988
rect 200684 245924 200685 245988
rect 200619 245923 200685 245924
rect 199794 237454 200414 238182
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 200622 236605 200682 245923
rect 236499 239732 236565 239733
rect 236499 239668 236500 239732
rect 236564 239668 236565 239732
rect 236499 239667 236565 239668
rect 238523 239732 238589 239733
rect 238523 239668 238524 239732
rect 238588 239668 238589 239732
rect 238523 239667 238589 239668
rect 200619 236604 200685 236605
rect 200619 236540 200620 236604
rect 200684 236540 200685 236604
rect 200619 236539 200685 236540
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 197123 93532 197189 93533
rect 197123 93468 197124 93532
rect 197188 93468 197189 93532
rect 197123 93467 197189 93468
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 205174 204134 238182
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 208894 207854 238182
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 212614 211574 238182
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 217794 219454 218414 238182
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 223174 222134 238182
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 225234 226894 225854 238182
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 228954 230614 229574 238182
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228771 181524 228837 181525
rect 228771 181460 228772 181524
rect 228836 181460 228837 181524
rect 228771 181459 228837 181460
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 228774 174450 228834 181459
rect 228954 178000 229574 194058
rect 235794 237454 236414 238182
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 233371 186964 233437 186965
rect 233371 186900 233372 186964
rect 233436 186900 233437 186964
rect 233371 186899 233437 186900
rect 233187 177444 233253 177445
rect 233187 177380 233188 177444
rect 233252 177380 233253 177444
rect 233187 177379 233253 177380
rect 228774 174390 229202 174450
rect 229142 174317 229202 174390
rect 229139 174316 229205 174317
rect 229139 174252 229140 174316
rect 229204 174252 229205 174316
rect 229139 174251 229205 174252
rect 214419 173228 214485 173229
rect 214419 173164 214420 173228
rect 214484 173164 214485 173228
rect 214419 173163 214485 173164
rect 214422 160853 214482 173163
rect 221207 165454 221527 165486
rect 221207 165218 221249 165454
rect 221485 165218 221527 165454
rect 221207 165134 221527 165218
rect 221207 164898 221249 165134
rect 221485 164898 221527 165134
rect 221207 164866 221527 164898
rect 224471 165454 224791 165486
rect 224471 165218 224513 165454
rect 224749 165218 224791 165454
rect 224471 165134 224791 165218
rect 224471 164898 224513 165134
rect 224749 164898 224791 165134
rect 224471 164866 224791 164898
rect 214419 160852 214485 160853
rect 214419 160788 214420 160852
rect 214484 160788 214485 160852
rect 214419 160787 214485 160788
rect 232451 153236 232517 153237
rect 232451 153172 232452 153236
rect 232516 153172 232517 153236
rect 232451 153171 232517 153172
rect 219575 147454 219895 147486
rect 219575 147218 219617 147454
rect 219853 147218 219895 147454
rect 219575 147134 219895 147218
rect 219575 146898 219617 147134
rect 219853 146898 219895 147134
rect 219575 146866 219895 146898
rect 222839 147454 223159 147486
rect 222839 147218 222881 147454
rect 223117 147218 223159 147454
rect 222839 147134 223159 147218
rect 222839 146898 222881 147134
rect 223117 146898 223159 147134
rect 222839 146866 223159 146898
rect 226103 147454 226423 147486
rect 226103 147218 226145 147454
rect 226381 147218 226423 147454
rect 226103 147134 226423 147218
rect 226103 146898 226145 147134
rect 226381 146898 226423 147134
rect 226103 146866 226423 146898
rect 230979 144124 231045 144125
rect 230979 144060 230980 144124
rect 231044 144060 231045 144124
rect 230979 144059 231045 144060
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 221207 129454 221527 129486
rect 221207 129218 221249 129454
rect 221485 129218 221527 129454
rect 221207 129134 221527 129218
rect 221207 128898 221249 129134
rect 221485 128898 221527 129134
rect 221207 128866 221527 128898
rect 224471 129454 224791 129486
rect 224471 129218 224513 129454
rect 224749 129218 224791 129454
rect 224471 129134 224791 129218
rect 224471 128898 224513 129134
rect 224749 128898 224791 129134
rect 224471 128866 224791 128898
rect 230982 125493 231042 144059
rect 232454 139229 232514 153171
rect 232451 139228 232517 139229
rect 232451 139164 232452 139228
rect 232516 139164 232517 139228
rect 232451 139163 232517 139164
rect 233190 138821 233250 177379
rect 233374 148749 233434 186899
rect 234659 178804 234725 178805
rect 234659 178740 234660 178804
rect 234724 178740 234725 178804
rect 234659 178739 234725 178740
rect 234662 163437 234722 178739
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 234659 163436 234725 163437
rect 234659 163372 234660 163436
rect 234724 163372 234725 163436
rect 234659 163371 234725 163372
rect 233371 148748 233437 148749
rect 233371 148684 233372 148748
rect 233436 148684 233437 148748
rect 233371 148683 233437 148684
rect 233739 141132 233805 141133
rect 233739 141068 233740 141132
rect 233804 141068 233805 141132
rect 233739 141067 233805 141068
rect 233187 138820 233253 138821
rect 233187 138756 233188 138820
rect 233252 138756 233253 138820
rect 233187 138755 233253 138756
rect 232451 137188 232517 137189
rect 232451 137124 232452 137188
rect 232516 137124 232517 137188
rect 232451 137123 232517 137124
rect 230979 125492 231045 125493
rect 230979 125428 230980 125492
rect 231044 125428 231045 125492
rect 230979 125427 231045 125428
rect 219575 111454 219895 111486
rect 219575 111218 219617 111454
rect 219853 111218 219895 111454
rect 219575 111134 219895 111218
rect 219575 110898 219617 111134
rect 219853 110898 219895 111134
rect 219575 110866 219895 110898
rect 222839 111454 223159 111486
rect 222839 111218 222881 111454
rect 223117 111218 223159 111454
rect 222839 111134 223159 111218
rect 222839 110898 222881 111134
rect 223117 110898 223159 111134
rect 222839 110866 223159 110898
rect 226103 111454 226423 111486
rect 226103 111218 226145 111454
rect 226381 111218 226423 111454
rect 226103 111134 226423 111218
rect 226103 110898 226145 111134
rect 226381 110898 226423 111134
rect 226103 110866 226423 110898
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 214419 103596 214485 103597
rect 214419 103532 214420 103596
rect 214484 103532 214485 103596
rect 214419 103531 214485 103532
rect 214422 91085 214482 103531
rect 229139 97068 229205 97069
rect 229139 97004 229140 97068
rect 229204 97004 229205 97068
rect 229139 97003 229205 97004
rect 229142 96630 229202 97003
rect 228958 96570 229202 96630
rect 228958 95301 229018 96570
rect 227667 95300 227733 95301
rect 227667 95236 227668 95300
rect 227732 95236 227733 95300
rect 227667 95235 227733 95236
rect 228955 95300 229021 95301
rect 228955 95236 228956 95300
rect 229020 95236 229021 95300
rect 228955 95235 229021 95236
rect 214419 91084 214485 91085
rect 214419 91020 214420 91084
rect 214484 91020 214485 91084
rect 214419 91019 214485 91020
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 227670 44845 227730 95235
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 227667 44844 227733 44845
rect 227667 44780 227668 44844
rect 227732 44780 227733 44844
rect 227667 44779 227733 44780
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 232454 10437 232514 137123
rect 233742 98021 233802 141067
rect 235794 129454 236414 164898
rect 236502 163845 236562 239667
rect 237419 239596 237485 239597
rect 237419 239532 237420 239596
rect 237484 239532 237485 239596
rect 237419 239531 237485 239532
rect 236499 163844 236565 163845
rect 236499 163780 236500 163844
rect 236564 163780 236565 163844
rect 236499 163779 236565 163780
rect 237422 153917 237482 239531
rect 237603 177308 237669 177309
rect 237603 177244 237604 177308
rect 237668 177244 237669 177308
rect 237603 177243 237669 177244
rect 237419 153916 237485 153917
rect 237419 153852 237420 153916
rect 237484 153852 237485 153916
rect 237419 153851 237485 153852
rect 237606 141677 237666 177243
rect 237603 141676 237669 141677
rect 237603 141612 237604 141676
rect 237668 141612 237669 141676
rect 237603 141611 237669 141612
rect 236499 139908 236565 139909
rect 236499 139844 236500 139908
rect 236564 139844 236565 139908
rect 236499 139843 236565 139844
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 233739 98020 233805 98021
rect 233739 97956 233740 98020
rect 233804 97956 233805 98020
rect 233739 97955 233805 97956
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 236502 62797 236562 139843
rect 238526 137869 238586 239667
rect 241651 239460 241717 239461
rect 241651 239396 241652 239460
rect 241716 239396 241717 239460
rect 241651 239395 241717 239396
rect 239514 205174 240134 238182
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 241654 180810 241714 239395
rect 241470 180750 241714 180810
rect 243234 208894 243854 238182
rect 244779 235244 244845 235245
rect 244779 235180 244780 235244
rect 244844 235180 244845 235244
rect 244779 235179 244845 235180
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 240363 175948 240429 175949
rect 240363 175884 240364 175948
rect 240428 175884 240429 175948
rect 240363 175883 240429 175884
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 238523 137868 238589 137869
rect 238523 137804 238524 137868
rect 238588 137804 238589 137868
rect 238523 137803 238589 137804
rect 239514 133174 240134 168618
rect 240366 136373 240426 175883
rect 241470 151830 241530 180750
rect 241651 180164 241717 180165
rect 241651 180100 241652 180164
rect 241716 180100 241717 180164
rect 241651 180099 241717 180100
rect 241654 171150 241714 180099
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 241654 171090 241898 171150
rect 241470 151770 241714 151830
rect 241654 138277 241714 151770
rect 241838 144941 241898 171090
rect 241835 144940 241901 144941
rect 241835 144876 241836 144940
rect 241900 144876 241901 144940
rect 241835 144875 241901 144876
rect 241651 138276 241717 138277
rect 241651 138212 241652 138276
rect 241716 138212 241717 138276
rect 241651 138211 241717 138212
rect 243234 136894 243854 172338
rect 244782 139773 244842 235179
rect 246954 212614 247574 238182
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 249750 145621 249810 269179
rect 250302 160037 250362 281691
rect 251219 274956 251285 274957
rect 251219 274892 251220 274956
rect 251284 274892 251285 274956
rect 251219 274891 251285 274892
rect 250299 160036 250365 160037
rect 250299 159972 250300 160036
rect 250364 159972 250365 160036
rect 250299 159971 250365 159972
rect 251222 155277 251282 274891
rect 252507 246396 252573 246397
rect 252507 246332 252508 246396
rect 252572 246332 252573 246396
rect 252507 246331 252573 246332
rect 251219 155276 251285 155277
rect 251219 155212 251220 155276
rect 251284 155212 251285 155276
rect 251219 155211 251285 155212
rect 252510 151061 252570 246331
rect 253062 177309 253122 285091
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 255822 238645 255882 576811
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 258395 296988 258461 296989
rect 258395 296924 258396 296988
rect 258460 296924 258461 296988
rect 258395 296923 258461 296924
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 258398 277410 258458 296923
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 255819 238644 255885 238645
rect 255819 238580 255820 238644
rect 255884 238580 255885 238644
rect 255819 238579 255885 238580
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253059 177308 253125 177309
rect 253059 177244 253060 177308
rect 253124 177244 253125 177308
rect 253059 177243 253125 177244
rect 252507 151060 252573 151061
rect 252507 150996 252508 151060
rect 252572 150996 252573 151060
rect 252507 150995 252573 150996
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 249747 145620 249813 145621
rect 249747 145556 249748 145620
rect 249812 145556 249813 145620
rect 249747 145555 249813 145556
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 244779 139772 244845 139773
rect 244779 139708 244780 139772
rect 244844 139708 244845 139772
rect 244779 139707 244845 139708
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 240363 136372 240429 136373
rect 240363 136308 240364 136372
rect 240428 136308 240429 136372
rect 240363 136307 240429 136308
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 236499 62796 236565 62797
rect 236499 62732 236500 62796
rect 236564 62732 236565 62796
rect 236499 62731 236565 62732
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 232451 10436 232517 10437
rect 232451 10372 232452 10436
rect 232516 10372 232517 10436
rect 232451 10371 232517 10372
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 104614 247574 140058
rect 251771 139772 251837 139773
rect 251771 139708 251772 139772
rect 251836 139708 251837 139772
rect 251771 139707 251837 139708
rect 250299 130252 250365 130253
rect 250299 130188 250300 130252
rect 250364 130188 250365 130252
rect 250299 130187 250365 130188
rect 249011 114884 249077 114885
rect 249011 114820 249012 114884
rect 249076 114820 249077 114884
rect 249011 114819 249077 114820
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 249014 7581 249074 114819
rect 250302 17237 250362 130187
rect 250299 17236 250365 17237
rect 250299 17172 250300 17236
rect 250364 17172 250365 17236
rect 250299 17171 250365 17172
rect 251774 10301 251834 139707
rect 253794 111454 254414 146898
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 258214 277350 258458 277410
rect 258214 151830 258274 277350
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 258214 151770 258458 151830
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 255819 128484 255885 128485
rect 255819 128420 255820 128484
rect 255884 128420 255885 128484
rect 255819 128419 255885 128420
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253059 102508 253125 102509
rect 253059 102444 253060 102508
rect 253124 102444 253125 102508
rect 253059 102443 253125 102444
rect 253062 57221 253122 102443
rect 253243 96660 253309 96661
rect 253243 96596 253244 96660
rect 253308 96596 253309 96660
rect 253243 96595 253309 96596
rect 253059 57220 253125 57221
rect 253059 57156 253060 57220
rect 253124 57156 253125 57220
rect 253059 57155 253125 57156
rect 253246 55861 253306 96595
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253243 55860 253309 55861
rect 253243 55796 253244 55860
rect 253308 55796 253309 55860
rect 253243 55795 253309 55796
rect 253794 39454 254414 74898
rect 255822 40629 255882 128419
rect 257514 115174 258134 150618
rect 258398 142085 258458 151770
rect 258395 142084 258461 142085
rect 258395 142020 258396 142084
rect 258460 142020 258461 142084
rect 258395 142019 258461 142020
rect 258763 133244 258829 133245
rect 258763 133180 258764 133244
rect 258828 133180 258829 133244
rect 258763 133179 258829 133180
rect 258579 118828 258645 118829
rect 258579 118764 258580 118828
rect 258644 118764 258645 118828
rect 258579 118763 258645 118764
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 258582 51781 258642 118763
rect 258766 72453 258826 133179
rect 260051 129844 260117 129845
rect 260051 129780 260052 129844
rect 260116 129780 260117 129844
rect 260051 129779 260117 129780
rect 258763 72452 258829 72453
rect 258763 72388 258764 72452
rect 258828 72388 258829 72452
rect 258763 72387 258829 72388
rect 258579 51780 258645 51781
rect 258579 51716 258580 51780
rect 258644 51716 258645 51780
rect 258579 51715 258645 51716
rect 260054 46205 260114 129779
rect 261234 118894 261854 154338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 178000 272414 200898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 278819 279036 278885 279037
rect 278819 278972 278820 279036
rect 278884 278972 278885 279036
rect 278819 278971 278885 278972
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 178000 276134 204618
rect 276611 185604 276677 185605
rect 276611 185540 276612 185604
rect 276676 185540 276677 185604
rect 276611 185539 276677 185540
rect 276614 177581 276674 185539
rect 276611 177580 276677 177581
rect 276611 177516 276612 177580
rect 276676 177516 276677 177580
rect 276611 177515 276677 177516
rect 278822 175130 278882 278971
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 178000 279854 208338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 288387 294132 288453 294133
rect 288387 294068 288388 294132
rect 288452 294068 288453 294132
rect 288387 294067 288453 294068
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 287099 197980 287165 197981
rect 287099 197916 287100 197980
rect 287164 197916 287165 197980
rect 287099 197915 287165 197916
rect 285627 193900 285693 193901
rect 285627 193836 285628 193900
rect 285692 193836 285693 193900
rect 285627 193835 285693 193836
rect 284339 181524 284405 181525
rect 284339 181460 284340 181524
rect 284404 181460 284405 181524
rect 284339 181459 284405 181460
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 281579 175948 281645 175949
rect 281579 175884 281580 175948
rect 281644 175884 281645 175948
rect 281579 175883 281645 175884
rect 279371 175132 279437 175133
rect 279371 175130 279372 175132
rect 278822 175070 279372 175130
rect 279371 175068 279372 175070
rect 279436 175068 279437 175132
rect 279371 175067 279437 175068
rect 268515 168604 268581 168605
rect 268515 168540 268516 168604
rect 268580 168540 268581 168604
rect 268515 168539 268581 168540
rect 268518 168197 268578 168539
rect 268515 168196 268581 168197
rect 268515 168132 268516 168196
rect 268580 168132 268581 168196
rect 268515 168131 268581 168132
rect 268515 167244 268581 167245
rect 268515 167180 268516 167244
rect 268580 167180 268581 167244
rect 268515 167179 268581 167180
rect 268518 166837 268578 167179
rect 268515 166836 268581 166837
rect 268515 166772 268516 166836
rect 268580 166772 268581 166836
rect 268515 166771 268581 166772
rect 272207 165454 272527 165486
rect 272207 165218 272249 165454
rect 272485 165218 272527 165454
rect 272207 165134 272527 165218
rect 272207 164898 272249 165134
rect 272485 164898 272527 165134
rect 272207 164866 272527 164898
rect 275471 165454 275791 165486
rect 275471 165218 275513 165454
rect 275749 165218 275791 165454
rect 275471 165134 275791 165218
rect 275471 164898 275513 165134
rect 275749 164898 275791 165134
rect 275471 164866 275791 164898
rect 268515 161668 268581 161669
rect 268515 161604 268516 161668
rect 268580 161604 268581 161668
rect 268515 161603 268581 161604
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 262811 128212 262877 128213
rect 262811 128148 262812 128212
rect 262876 128148 262877 128212
rect 262811 128147 262877 128148
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 260235 116108 260301 116109
rect 260235 116044 260236 116108
rect 260300 116044 260301 116108
rect 260235 116043 260301 116044
rect 260051 46204 260117 46205
rect 260051 46140 260052 46204
rect 260116 46140 260117 46204
rect 260051 46139 260117 46140
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 255819 40628 255885 40629
rect 255819 40564 255820 40628
rect 255884 40564 255885 40628
rect 255819 40563 255885 40564
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 251771 10300 251837 10301
rect 251771 10236 251772 10300
rect 251836 10236 251837 10300
rect 251771 10235 251837 10236
rect 249011 7580 249077 7581
rect 249011 7516 249012 7580
rect 249076 7516 249077 7580
rect 249011 7515 249077 7516
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 42618
rect 260238 33829 260298 116043
rect 261234 82894 261854 118338
rect 262075 102780 262141 102781
rect 262075 102716 262076 102780
rect 262140 102716 262141 102780
rect 262075 102715 262141 102716
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 260235 33828 260301 33829
rect 260235 33764 260236 33828
rect 260300 33764 260301 33828
rect 260235 33763 260301 33764
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 46338
rect 262078 22677 262138 102715
rect 262814 43485 262874 128147
rect 264099 126852 264165 126853
rect 264099 126788 264100 126852
rect 264164 126788 264165 126852
rect 264099 126787 264165 126788
rect 262995 114748 263061 114749
rect 262995 114684 262996 114748
rect 263060 114684 263061 114748
rect 262995 114683 263061 114684
rect 262998 71093 263058 114683
rect 262995 71092 263061 71093
rect 262995 71028 262996 71092
rect 263060 71028 263061 71092
rect 262995 71027 263061 71028
rect 262811 43484 262877 43485
rect 262811 43420 262812 43484
rect 262876 43420 262877 43484
rect 262811 43419 262877 43420
rect 264102 36549 264162 126787
rect 264954 122614 265574 158058
rect 268518 157317 268578 161603
rect 268515 157316 268581 157317
rect 268515 157252 268516 157316
rect 268580 157252 268581 157316
rect 268515 157251 268581 157252
rect 281582 157045 281642 175883
rect 281579 157044 281645 157045
rect 281579 156980 281580 157044
rect 281644 156980 281645 157044
rect 281579 156979 281645 156980
rect 268515 147932 268581 147933
rect 268515 147868 268516 147932
rect 268580 147868 268581 147932
rect 268515 147867 268581 147868
rect 268518 146165 268578 147867
rect 270575 147454 270895 147486
rect 270575 147218 270617 147454
rect 270853 147218 270895 147454
rect 270575 147134 270895 147218
rect 270575 146898 270617 147134
rect 270853 146898 270895 147134
rect 270575 146866 270895 146898
rect 273839 147454 274159 147486
rect 273839 147218 273881 147454
rect 274117 147218 274159 147454
rect 273839 147134 274159 147218
rect 273839 146898 273881 147134
rect 274117 146898 274159 147134
rect 273839 146866 274159 146898
rect 277103 147454 277423 147486
rect 277103 147218 277145 147454
rect 277381 147218 277423 147454
rect 277103 147134 277423 147218
rect 277103 146898 277145 147134
rect 277381 146898 277423 147134
rect 277103 146866 277423 146898
rect 268515 146164 268581 146165
rect 268515 146100 268516 146164
rect 268580 146100 268581 146164
rect 268515 146099 268581 146100
rect 268515 142356 268581 142357
rect 268515 142292 268516 142356
rect 268580 142292 268581 142356
rect 268515 142291 268581 142292
rect 268518 141949 268578 142291
rect 268515 141948 268581 141949
rect 268515 141884 268516 141948
rect 268580 141884 268581 141948
rect 268515 141883 268581 141884
rect 267779 141132 267845 141133
rect 267779 141068 267780 141132
rect 267844 141130 267845 141132
rect 267844 141070 268394 141130
rect 267844 141068 267845 141070
rect 267779 141067 267845 141068
rect 268334 140997 268394 141070
rect 268331 140996 268397 140997
rect 268331 140932 268332 140996
rect 268396 140932 268397 140996
rect 268331 140931 268397 140932
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 272207 129454 272527 129486
rect 272207 129218 272249 129454
rect 272485 129218 272527 129454
rect 272207 129134 272527 129218
rect 272207 128898 272249 129134
rect 272485 128898 272527 129134
rect 272207 128866 272527 128898
rect 275471 129454 275791 129486
rect 275471 129218 275513 129454
rect 275749 129218 275791 129454
rect 275471 129134 275791 129218
rect 275471 128898 275513 129134
rect 275749 128898 275791 129134
rect 275471 128866 275791 128898
rect 268515 128620 268581 128621
rect 268515 128556 268516 128620
rect 268580 128556 268581 128620
rect 268515 128555 268581 128556
rect 268518 128213 268578 128555
rect 268515 128212 268581 128213
rect 268515 128148 268516 128212
rect 268580 128148 268581 128212
rect 268515 128147 268581 128148
rect 268515 127260 268581 127261
rect 268515 127196 268516 127260
rect 268580 127196 268581 127260
rect 268515 127195 268581 127196
rect 268518 126853 268578 127195
rect 268515 126852 268581 126853
rect 268515 126788 268516 126852
rect 268580 126788 268581 126852
rect 268515 126787 268581 126788
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264283 120460 264349 120461
rect 264283 120396 264284 120460
rect 264348 120396 264349 120460
rect 264283 120395 264349 120396
rect 264286 47565 264346 120395
rect 264954 86614 265574 122058
rect 268515 121684 268581 121685
rect 268515 121620 268516 121684
rect 268580 121620 268581 121684
rect 268515 121619 268581 121620
rect 268518 119917 268578 121619
rect 268515 119916 268581 119917
rect 268515 119852 268516 119916
rect 268580 119852 268581 119916
rect 268515 119851 268581 119852
rect 268331 116108 268397 116109
rect 268331 116044 268332 116108
rect 268396 116044 268397 116108
rect 268331 116043 268397 116044
rect 267779 115972 267845 115973
rect 267779 115908 267780 115972
rect 267844 115970 267845 115972
rect 268334 115970 268394 116043
rect 267844 115910 268394 115970
rect 267844 115908 267845 115910
rect 267779 115907 267845 115908
rect 270575 111454 270895 111486
rect 270575 111218 270617 111454
rect 270853 111218 270895 111454
rect 270575 111134 270895 111218
rect 270575 110898 270617 111134
rect 270853 110898 270895 111134
rect 270575 110866 270895 110898
rect 273839 111454 274159 111486
rect 273839 111218 273881 111454
rect 274117 111218 274159 111454
rect 273839 111134 274159 111218
rect 273839 110898 273881 111134
rect 274117 110898 274159 111134
rect 273839 110866 274159 110898
rect 277103 111454 277423 111486
rect 277103 111218 277145 111454
rect 277381 111218 277423 111454
rect 277103 111134 277423 111218
rect 277103 110898 277145 111134
rect 277381 110898 277423 111134
rect 277103 110866 277423 110898
rect 268331 107948 268397 107949
rect 268331 107884 268332 107948
rect 268396 107884 268397 107948
rect 268331 107883 268397 107884
rect 268334 107541 268394 107883
rect 268331 107540 268397 107541
rect 268331 107476 268332 107540
rect 268396 107476 268397 107540
rect 268331 107475 268397 107476
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 268331 102780 268397 102781
rect 268331 102778 268332 102780
rect 267782 102718 268332 102778
rect 267782 102509 267842 102718
rect 268331 102716 268332 102718
rect 268396 102716 268397 102780
rect 268331 102715 268397 102716
rect 267779 102508 267845 102509
rect 267779 102444 267780 102508
rect 267844 102444 267845 102508
rect 267779 102443 267845 102444
rect 266859 98836 266925 98837
rect 266859 98772 266860 98836
rect 266924 98772 266925 98836
rect 266859 98771 266925 98772
rect 265755 96660 265821 96661
rect 265755 96596 265756 96660
rect 265820 96596 265821 96660
rect 265755 96595 265821 96596
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264283 47564 264349 47565
rect 264283 47500 264284 47564
rect 264348 47500 264349 47564
rect 264283 47499 264349 47500
rect 264099 36548 264165 36549
rect 264099 36484 264100 36548
rect 264164 36484 264165 36548
rect 264099 36483 264165 36484
rect 262075 22676 262141 22677
rect 262075 22612 262076 22676
rect 262140 22612 262141 22676
rect 262075 22611 262141 22612
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 265758 4861 265818 96595
rect 266862 11661 266922 98771
rect 268331 96796 268397 96797
rect 268331 96732 268332 96796
rect 268396 96732 268397 96796
rect 268331 96731 268397 96732
rect 267779 96660 267845 96661
rect 267779 96596 267780 96660
rect 267844 96630 267845 96660
rect 268334 96630 268394 96731
rect 267844 96596 268394 96630
rect 267779 96595 268394 96596
rect 267782 96570 268394 96595
rect 271794 93454 272414 94000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 266859 11660 266925 11661
rect 266859 11596 266860 11660
rect 266924 11596 266925 11660
rect 266859 11595 266925 11596
rect 265755 4860 265821 4861
rect 265755 4796 265756 4860
rect 265820 4796 265821 4860
rect 265755 4795 265821 4796
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 94000
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 94000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 104058
rect 284342 104005 284402 181459
rect 285630 143173 285690 193835
rect 285627 143172 285693 143173
rect 285627 143108 285628 143172
rect 285692 143108 285693 143172
rect 285627 143107 285693 143108
rect 287102 127125 287162 197915
rect 287283 184244 287349 184245
rect 287283 184180 287284 184244
rect 287348 184180 287349 184244
rect 287283 184179 287349 184180
rect 287286 128757 287346 184179
rect 287283 128756 287349 128757
rect 287283 128692 287284 128756
rect 287348 128692 287349 128756
rect 287283 128691 287349 128692
rect 287099 127124 287165 127125
rect 287099 127060 287100 127124
rect 287164 127060 287165 127124
rect 287099 127059 287165 127060
rect 288390 104957 288450 294067
rect 288571 292636 288637 292637
rect 288571 292572 288572 292636
rect 288636 292572 288637 292636
rect 288571 292571 288637 292572
rect 288574 131205 288634 292571
rect 289794 291454 290414 326898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 291147 299572 291213 299573
rect 291147 299508 291148 299572
rect 291212 299508 291213 299572
rect 291147 299507 291213 299508
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 290595 191180 290661 191181
rect 290595 191116 290596 191180
rect 290660 191116 290661 191180
rect 290595 191115 290661 191116
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 288571 131204 288637 131205
rect 288571 131140 288572 131204
rect 288636 131140 288637 131204
rect 288571 131139 288637 131140
rect 289794 111454 290414 146898
rect 290598 134197 290658 191115
rect 290595 134196 290661 134197
rect 290595 134132 290596 134196
rect 290660 134132 290661 134196
rect 290595 134131 290661 134132
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 288387 104956 288453 104957
rect 288387 104892 288388 104956
rect 288452 104892 288453 104956
rect 288387 104891 288453 104892
rect 284339 104004 284405 104005
rect 284339 103940 284340 104004
rect 284404 103940 284405 104004
rect 284339 103939 284405 103940
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 75454 290414 110898
rect 291150 109581 291210 299507
rect 293514 295174 294134 330618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 295563 298212 295629 298213
rect 295563 298148 295564 298212
rect 295628 298148 295629 298212
rect 295563 298147 295629 298148
rect 295379 296852 295445 296853
rect 295379 296788 295380 296852
rect 295444 296788 295445 296852
rect 295379 296787 295445 296788
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 294275 191044 294341 191045
rect 294275 190980 294276 191044
rect 294340 190980 294341 191044
rect 294275 190979 294341 190980
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 292619 181388 292685 181389
rect 292619 181324 292620 181388
rect 292684 181324 292685 181388
rect 292619 181323 292685 181324
rect 291331 177444 291397 177445
rect 291331 177380 291332 177444
rect 291396 177380 291397 177444
rect 291331 177379 291397 177380
rect 291334 140861 291394 177379
rect 291331 140860 291397 140861
rect 291331 140796 291332 140860
rect 291396 140796 291397 140860
rect 291331 140795 291397 140796
rect 292622 113253 292682 181323
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 294278 121549 294338 190979
rect 294275 121548 294341 121549
rect 294275 121484 294276 121548
rect 294340 121484 294341 121548
rect 294275 121483 294341 121484
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 292619 113252 292685 113253
rect 292619 113188 292620 113252
rect 292684 113188 292685 113252
rect 292619 113187 292685 113188
rect 291147 109580 291213 109581
rect 291147 109516 291148 109580
rect 291212 109516 291213 109580
rect 291147 109515 291213 109516
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 79174 294134 114618
rect 295382 109173 295442 296787
rect 295566 171189 295626 298147
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 298691 228308 298757 228309
rect 298691 228244 298692 228308
rect 298756 228244 298757 228308
rect 298691 228243 298757 228244
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 295563 171188 295629 171189
rect 295563 171124 295564 171188
rect 295628 171124 295629 171188
rect 296667 171188 296733 171189
rect 296667 171150 296668 171188
rect 295563 171123 295629 171124
rect 296486 171124 296668 171150
rect 296732 171124 296733 171188
rect 296486 171123 296733 171124
rect 296486 171090 296730 171123
rect 296486 135285 296546 171090
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 296483 135284 296549 135285
rect 296483 135220 296484 135284
rect 296548 135220 296549 135284
rect 296483 135219 296549 135220
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 295379 109172 295445 109173
rect 295379 109108 295380 109172
rect 295444 109108 295445 109172
rect 295379 109107 295445 109108
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 298694 59397 298754 228243
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 298691 59396 298757 59397
rect 298691 59332 298692 59396
rect 298756 59332 298757 59396
rect 298691 59331 298757 59332
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 219810 273218 220046 273454
rect 219810 272898 220046 273134
rect 204450 255218 204686 255454
rect 204450 254898 204686 255134
rect 235170 255218 235406 255454
rect 235170 254898 235406 255134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 221249 165218 221485 165454
rect 221249 164898 221485 165134
rect 224513 165218 224749 165454
rect 224513 164898 224749 165134
rect 219617 147218 219853 147454
rect 219617 146898 219853 147134
rect 222881 147218 223117 147454
rect 222881 146898 223117 147134
rect 226145 147218 226381 147454
rect 226145 146898 226381 147134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 221249 129218 221485 129454
rect 221249 128898 221485 129134
rect 224513 129218 224749 129454
rect 224513 128898 224749 129134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 219617 111218 219853 111454
rect 219617 110898 219853 111134
rect 222881 111218 223117 111454
rect 222881 110898 223117 111134
rect 226145 111218 226381 111454
rect 226145 110898 226381 111134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 272249 165218 272485 165454
rect 272249 164898 272485 165134
rect 275513 165218 275749 165454
rect 275513 164898 275749 165134
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 270617 147218 270853 147454
rect 270617 146898 270853 147134
rect 273881 147218 274117 147454
rect 273881 146898 274117 147134
rect 277145 147218 277381 147454
rect 277145 146898 277381 147134
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 272249 129218 272485 129454
rect 272249 128898 272485 129134
rect 275513 129218 275749 129454
rect 275513 128898 275749 129134
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 270617 111218 270853 111454
rect 270617 110898 270853 111134
rect 273881 111218 274117 111454
rect 273881 110898 274117 111134
rect 277145 111218 277381 111454
rect 277145 110898 277381 111134
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219810 273454
rect 220046 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219810 273134
rect 220046 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204450 255454
rect 204686 255218 235170 255454
rect 235406 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204450 255134
rect 204686 254898 235170 255134
rect 235406 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 221249 165454
rect 221485 165218 224513 165454
rect 224749 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 272249 165454
rect 272485 165218 275513 165454
rect 275749 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 221249 165134
rect 221485 164898 224513 165134
rect 224749 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 272249 165134
rect 272485 164898 275513 165134
rect 275749 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 219617 147454
rect 219853 147218 222881 147454
rect 223117 147218 226145 147454
rect 226381 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 270617 147454
rect 270853 147218 273881 147454
rect 274117 147218 277145 147454
rect 277381 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 219617 147134
rect 219853 146898 222881 147134
rect 223117 146898 226145 147134
rect 226381 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 270617 147134
rect 270853 146898 273881 147134
rect 274117 146898 277145 147134
rect 277381 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 221249 129454
rect 221485 129218 224513 129454
rect 224749 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 272249 129454
rect 272485 129218 275513 129454
rect 275749 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 221249 129134
rect 221485 128898 224513 129134
rect 224749 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 272249 129134
rect 272485 128898 275513 129134
rect 275749 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 219617 111454
rect 219853 111218 222881 111454
rect 223117 111218 226145 111454
rect 226381 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 270617 111454
rect 270853 111218 273881 111454
rect 274117 111218 277145 111454
rect 277381 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 219617 111134
rect 219853 110898 222881 111134
rect 223117 110898 226145 111134
rect 226381 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 270617 111134
rect 270853 110898 273881 111134
rect 274117 110898 277145 111134
rect 277381 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 268000 0 1 96000
box 0 0 12000 79688
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 12000 79688
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 200200 0 1 240182
box 0 0 50000 52000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 238182 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 294182 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 238182 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 294182 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 238182 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 294182 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 238182 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 294182 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 294182 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 294182 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 178000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 238182 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 238182 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 294182 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 294182 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 294182 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 294182 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 178000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 294182 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 294182 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 178000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
