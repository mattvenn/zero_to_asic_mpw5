VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_hack_soc_dffram
  CLASS BLOCK ;
  FOREIGN wrapped_hack_soc_dffram ;
  ORIGIN 0.000 0.000 ;
  SIZE 372.350 BY 398.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 338.680 372.350 339.280 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 394.000 63.850 398.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 394.000 52.350 398.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 394.000 40.390 398.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 394.000 28.890 398.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 282.240 372.350 282.840 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 276.800 372.350 277.400 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 394.000 17.390 398.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 394.000 5.890 398.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 58.520 372.350 59.120 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 53.080 372.350 53.680 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 333.240 372.350 333.840 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 271.360 372.350 271.960 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 265.920 372.350 266.520 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 46.960 372.350 47.560 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 41.520 372.350 42.120 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 36.080 372.350 36.680 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 30.640 372.350 31.240 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 24.520 372.350 25.120 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 260.480 372.350 261.080 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 254.360 372.350 254.960 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 248.920 372.350 249.520 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 327.120 372.350 327.720 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 19.080 372.350 19.680 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 13.640 372.350 14.240 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 8.200 372.350 8.800 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 2.760 372.350 3.360 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 243.480 372.350 244.080 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 238.040 372.350 238.640 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 231.920 372.350 232.520 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 226.480 372.350 227.080 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 321.680 372.350 322.280 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 316.240 372.350 316.840 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 310.800 372.350 311.400 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 304.680 372.350 305.280 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 299.240 372.350 299.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 293.800 372.350 294.400 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 288.360 372.350 288.960 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 394.000 366.070 398.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 394.000 354.570 398.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 394.000 343.070 398.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 394.000 331.110 398.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 394.000 319.610 398.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 394.000 308.110 398.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 394.000 296.610 398.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 394.000 284.650 398.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 394.000 273.150 398.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 394.000 261.650 398.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 394.000 249.690 398.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 394.000 238.190 398.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 394.000 226.690 398.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 394.000 215.190 398.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 394.000 203.230 398.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 394.000 191.730 398.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 394.000 180.230 398.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 221.040 372.350 221.640 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 164.600 372.350 165.200 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 159.160 372.350 159.760 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 153.720 372.350 154.320 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 148.280 372.350 148.880 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 142.160 372.350 142.760 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 136.720 372.350 137.320 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 131.280 372.350 131.880 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 125.840 372.350 126.440 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 120.400 372.350 121.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 114.280 372.350 114.880 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 215.600 372.350 216.200 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 108.840 372.350 109.440 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 103.400 372.350 104.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 97.960 372.350 98.560 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 91.840 372.350 92.440 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 86.400 372.350 87.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 80.960 372.350 81.560 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 75.520 372.350 76.120 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 69.400 372.350 70.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 63.960 372.350 64.560 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 394.000 168.270 398.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 209.480 372.350 210.080 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 394.000 156.770 398.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 394.000 145.270 398.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 394.000 133.770 398.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 394.000 121.810 398.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 394.000 110.310 398.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 394.000 98.810 398.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 394.000 86.850 398.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 394.000 75.350 398.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 204.040 372.350 204.640 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 198.600 372.350 199.200 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 193.160 372.350 193.760 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 187.040 372.350 187.640 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 181.600 372.350 182.200 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 176.160 372.350 176.760 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 170.720 372.350 171.320 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 361.120 372.350 361.720 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 355.680 372.350 356.280 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 349.560 372.350 350.160 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 344.120 372.350 344.720 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 394.440 372.350 395.040 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 389.000 372.350 389.600 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 383.560 372.350 384.160 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 378.120 372.350 378.720 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.080 4.000 376.680 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 372.000 372.350 372.600 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 368.350 366.560 372.350 367.160 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 386.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 386.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 386.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 386.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 386.480 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 366.620 386.325 ;
      LAYER met1 ;
        RECT 2.830 7.860 368.850 386.480 ;
      LAYER met2 ;
        RECT 2.860 393.720 5.330 394.810 ;
        RECT 6.170 393.720 16.830 394.810 ;
        RECT 17.670 393.720 28.330 394.810 ;
        RECT 29.170 393.720 39.830 394.810 ;
        RECT 40.670 393.720 51.790 394.810 ;
        RECT 52.630 393.720 63.290 394.810 ;
        RECT 64.130 393.720 74.790 394.810 ;
        RECT 75.630 393.720 86.290 394.810 ;
        RECT 87.130 393.720 98.250 394.810 ;
        RECT 99.090 393.720 109.750 394.810 ;
        RECT 110.590 393.720 121.250 394.810 ;
        RECT 122.090 393.720 133.210 394.810 ;
        RECT 134.050 393.720 144.710 394.810 ;
        RECT 145.550 393.720 156.210 394.810 ;
        RECT 157.050 393.720 167.710 394.810 ;
        RECT 168.550 393.720 179.670 394.810 ;
        RECT 180.510 393.720 191.170 394.810 ;
        RECT 192.010 393.720 202.670 394.810 ;
        RECT 203.510 393.720 214.630 394.810 ;
        RECT 215.470 393.720 226.130 394.810 ;
        RECT 226.970 393.720 237.630 394.810 ;
        RECT 238.470 393.720 249.130 394.810 ;
        RECT 249.970 393.720 261.090 394.810 ;
        RECT 261.930 393.720 272.590 394.810 ;
        RECT 273.430 393.720 284.090 394.810 ;
        RECT 284.930 393.720 296.050 394.810 ;
        RECT 296.890 393.720 307.550 394.810 ;
        RECT 308.390 393.720 319.050 394.810 ;
        RECT 319.890 393.720 330.550 394.810 ;
        RECT 331.390 393.720 342.510 394.810 ;
        RECT 343.350 393.720 354.010 394.810 ;
        RECT 354.850 393.720 365.510 394.810 ;
        RECT 366.350 393.720 368.820 394.810 ;
        RECT 2.860 4.280 368.820 393.720 ;
        RECT 3.410 2.875 8.550 4.280 ;
        RECT 9.390 2.875 14.530 4.280 ;
        RECT 15.370 2.875 20.510 4.280 ;
        RECT 21.350 2.875 26.490 4.280 ;
        RECT 27.330 2.875 32.470 4.280 ;
        RECT 33.310 2.875 38.450 4.280 ;
        RECT 39.290 2.875 44.430 4.280 ;
        RECT 45.270 2.875 50.410 4.280 ;
        RECT 51.250 2.875 56.390 4.280 ;
        RECT 57.230 2.875 62.370 4.280 ;
        RECT 63.210 2.875 68.350 4.280 ;
        RECT 69.190 2.875 74.330 4.280 ;
        RECT 75.170 2.875 80.310 4.280 ;
        RECT 81.150 2.875 86.290 4.280 ;
        RECT 87.130 2.875 92.270 4.280 ;
        RECT 93.110 2.875 98.250 4.280 ;
        RECT 99.090 2.875 104.230 4.280 ;
        RECT 105.070 2.875 110.210 4.280 ;
        RECT 111.050 2.875 116.190 4.280 ;
        RECT 117.030 2.875 122.170 4.280 ;
        RECT 123.010 2.875 128.610 4.280 ;
        RECT 129.450 2.875 134.590 4.280 ;
        RECT 135.430 2.875 140.570 4.280 ;
        RECT 141.410 2.875 146.550 4.280 ;
        RECT 147.390 2.875 152.530 4.280 ;
        RECT 153.370 2.875 158.510 4.280 ;
        RECT 159.350 2.875 164.490 4.280 ;
        RECT 165.330 2.875 170.470 4.280 ;
        RECT 171.310 2.875 176.450 4.280 ;
        RECT 177.290 2.875 182.430 4.280 ;
        RECT 183.270 2.875 188.410 4.280 ;
        RECT 189.250 2.875 194.390 4.280 ;
        RECT 195.230 2.875 200.370 4.280 ;
        RECT 201.210 2.875 206.350 4.280 ;
        RECT 207.190 2.875 212.330 4.280 ;
        RECT 213.170 2.875 218.310 4.280 ;
        RECT 219.150 2.875 224.290 4.280 ;
        RECT 225.130 2.875 230.270 4.280 ;
        RECT 231.110 2.875 236.250 4.280 ;
        RECT 237.090 2.875 242.230 4.280 ;
        RECT 243.070 2.875 248.210 4.280 ;
        RECT 249.050 2.875 254.650 4.280 ;
        RECT 255.490 2.875 260.630 4.280 ;
        RECT 261.470 2.875 266.610 4.280 ;
        RECT 267.450 2.875 272.590 4.280 ;
        RECT 273.430 2.875 278.570 4.280 ;
        RECT 279.410 2.875 284.550 4.280 ;
        RECT 285.390 2.875 290.530 4.280 ;
        RECT 291.370 2.875 296.510 4.280 ;
        RECT 297.350 2.875 302.490 4.280 ;
        RECT 303.330 2.875 308.470 4.280 ;
        RECT 309.310 2.875 314.450 4.280 ;
        RECT 315.290 2.875 320.430 4.280 ;
        RECT 321.270 2.875 326.410 4.280 ;
        RECT 327.250 2.875 332.390 4.280 ;
        RECT 333.230 2.875 338.370 4.280 ;
        RECT 339.210 2.875 344.350 4.280 ;
        RECT 345.190 2.875 350.330 4.280 ;
        RECT 351.170 2.875 356.310 4.280 ;
        RECT 357.150 2.875 362.290 4.280 ;
        RECT 363.130 2.875 368.270 4.280 ;
      LAYER met3 ;
        RECT 4.000 385.920 368.350 386.405 ;
        RECT 4.400 384.560 368.350 385.920 ;
        RECT 4.400 384.520 367.950 384.560 ;
        RECT 4.000 383.160 367.950 384.520 ;
        RECT 4.000 379.120 368.350 383.160 ;
        RECT 4.000 377.720 367.950 379.120 ;
        RECT 4.000 377.080 368.350 377.720 ;
        RECT 4.400 375.680 368.350 377.080 ;
        RECT 4.000 373.000 368.350 375.680 ;
        RECT 4.000 371.600 367.950 373.000 ;
        RECT 4.000 368.920 368.350 371.600 ;
        RECT 4.400 367.560 368.350 368.920 ;
        RECT 4.400 367.520 367.950 367.560 ;
        RECT 4.000 366.160 367.950 367.520 ;
        RECT 4.000 362.120 368.350 366.160 ;
        RECT 4.000 360.720 367.950 362.120 ;
        RECT 4.000 360.080 368.350 360.720 ;
        RECT 4.400 358.680 368.350 360.080 ;
        RECT 4.000 356.680 368.350 358.680 ;
        RECT 4.000 355.280 367.950 356.680 ;
        RECT 4.000 351.920 368.350 355.280 ;
        RECT 4.400 350.560 368.350 351.920 ;
        RECT 4.400 350.520 367.950 350.560 ;
        RECT 4.000 349.160 367.950 350.520 ;
        RECT 4.000 345.120 368.350 349.160 ;
        RECT 4.000 343.720 367.950 345.120 ;
        RECT 4.000 343.080 368.350 343.720 ;
        RECT 4.400 341.680 368.350 343.080 ;
        RECT 4.000 339.680 368.350 341.680 ;
        RECT 4.000 338.280 367.950 339.680 ;
        RECT 4.000 334.920 368.350 338.280 ;
        RECT 4.400 334.240 368.350 334.920 ;
        RECT 4.400 333.520 367.950 334.240 ;
        RECT 4.000 332.840 367.950 333.520 ;
        RECT 4.000 328.120 368.350 332.840 ;
        RECT 4.000 326.720 367.950 328.120 ;
        RECT 4.000 326.080 368.350 326.720 ;
        RECT 4.400 324.680 368.350 326.080 ;
        RECT 4.000 322.680 368.350 324.680 ;
        RECT 4.000 321.280 367.950 322.680 ;
        RECT 4.000 317.920 368.350 321.280 ;
        RECT 4.400 317.240 368.350 317.920 ;
        RECT 4.400 316.520 367.950 317.240 ;
        RECT 4.000 315.840 367.950 316.520 ;
        RECT 4.000 311.800 368.350 315.840 ;
        RECT 4.000 310.400 367.950 311.800 ;
        RECT 4.000 309.760 368.350 310.400 ;
        RECT 4.400 308.360 368.350 309.760 ;
        RECT 4.000 305.680 368.350 308.360 ;
        RECT 4.000 304.280 367.950 305.680 ;
        RECT 4.000 300.920 368.350 304.280 ;
        RECT 4.400 300.240 368.350 300.920 ;
        RECT 4.400 299.520 367.950 300.240 ;
        RECT 4.000 298.840 367.950 299.520 ;
        RECT 4.000 294.800 368.350 298.840 ;
        RECT 4.000 293.400 367.950 294.800 ;
        RECT 4.000 292.760 368.350 293.400 ;
        RECT 4.400 291.360 368.350 292.760 ;
        RECT 4.000 289.360 368.350 291.360 ;
        RECT 4.000 287.960 367.950 289.360 ;
        RECT 4.000 283.920 368.350 287.960 ;
        RECT 4.400 283.240 368.350 283.920 ;
        RECT 4.400 282.520 367.950 283.240 ;
        RECT 4.000 281.840 367.950 282.520 ;
        RECT 4.000 277.800 368.350 281.840 ;
        RECT 4.000 276.400 367.950 277.800 ;
        RECT 4.000 275.760 368.350 276.400 ;
        RECT 4.400 274.360 368.350 275.760 ;
        RECT 4.000 272.360 368.350 274.360 ;
        RECT 4.000 270.960 367.950 272.360 ;
        RECT 4.000 266.920 368.350 270.960 ;
        RECT 4.400 265.520 367.950 266.920 ;
        RECT 4.000 261.480 368.350 265.520 ;
        RECT 4.000 260.080 367.950 261.480 ;
        RECT 4.000 258.760 368.350 260.080 ;
        RECT 4.400 257.360 368.350 258.760 ;
        RECT 4.000 255.360 368.350 257.360 ;
        RECT 4.000 253.960 367.950 255.360 ;
        RECT 4.000 249.920 368.350 253.960 ;
        RECT 4.400 248.520 367.950 249.920 ;
        RECT 4.000 244.480 368.350 248.520 ;
        RECT 4.000 243.080 367.950 244.480 ;
        RECT 4.000 241.760 368.350 243.080 ;
        RECT 4.400 240.360 368.350 241.760 ;
        RECT 4.000 239.040 368.350 240.360 ;
        RECT 4.000 237.640 367.950 239.040 ;
        RECT 4.000 233.600 368.350 237.640 ;
        RECT 4.400 232.920 368.350 233.600 ;
        RECT 4.400 232.200 367.950 232.920 ;
        RECT 4.000 231.520 367.950 232.200 ;
        RECT 4.000 227.480 368.350 231.520 ;
        RECT 4.000 226.080 367.950 227.480 ;
        RECT 4.000 224.760 368.350 226.080 ;
        RECT 4.400 223.360 368.350 224.760 ;
        RECT 4.000 222.040 368.350 223.360 ;
        RECT 4.000 220.640 367.950 222.040 ;
        RECT 4.000 216.600 368.350 220.640 ;
        RECT 4.400 215.200 367.950 216.600 ;
        RECT 4.000 210.480 368.350 215.200 ;
        RECT 4.000 209.080 367.950 210.480 ;
        RECT 4.000 207.760 368.350 209.080 ;
        RECT 4.400 206.360 368.350 207.760 ;
        RECT 4.000 205.040 368.350 206.360 ;
        RECT 4.000 203.640 367.950 205.040 ;
        RECT 4.000 199.600 368.350 203.640 ;
        RECT 4.400 198.200 367.950 199.600 ;
        RECT 4.000 194.160 368.350 198.200 ;
        RECT 4.000 192.760 367.950 194.160 ;
        RECT 4.000 190.760 368.350 192.760 ;
        RECT 4.400 189.360 368.350 190.760 ;
        RECT 4.000 188.040 368.350 189.360 ;
        RECT 4.000 186.640 367.950 188.040 ;
        RECT 4.000 182.600 368.350 186.640 ;
        RECT 4.400 181.200 367.950 182.600 ;
        RECT 4.000 177.160 368.350 181.200 ;
        RECT 4.000 175.760 367.950 177.160 ;
        RECT 4.000 173.760 368.350 175.760 ;
        RECT 4.400 172.360 368.350 173.760 ;
        RECT 4.000 171.720 368.350 172.360 ;
        RECT 4.000 170.320 367.950 171.720 ;
        RECT 4.000 165.600 368.350 170.320 ;
        RECT 4.400 164.200 367.950 165.600 ;
        RECT 4.000 160.160 368.350 164.200 ;
        RECT 4.000 158.760 367.950 160.160 ;
        RECT 4.000 157.440 368.350 158.760 ;
        RECT 4.400 156.040 368.350 157.440 ;
        RECT 4.000 154.720 368.350 156.040 ;
        RECT 4.000 153.320 367.950 154.720 ;
        RECT 4.000 149.280 368.350 153.320 ;
        RECT 4.000 148.600 367.950 149.280 ;
        RECT 4.400 147.880 367.950 148.600 ;
        RECT 4.400 147.200 368.350 147.880 ;
        RECT 4.000 143.160 368.350 147.200 ;
        RECT 4.000 141.760 367.950 143.160 ;
        RECT 4.000 140.440 368.350 141.760 ;
        RECT 4.400 139.040 368.350 140.440 ;
        RECT 4.000 137.720 368.350 139.040 ;
        RECT 4.000 136.320 367.950 137.720 ;
        RECT 4.000 132.280 368.350 136.320 ;
        RECT 4.000 131.600 367.950 132.280 ;
        RECT 4.400 130.880 367.950 131.600 ;
        RECT 4.400 130.200 368.350 130.880 ;
        RECT 4.000 126.840 368.350 130.200 ;
        RECT 4.000 125.440 367.950 126.840 ;
        RECT 4.000 123.440 368.350 125.440 ;
        RECT 4.400 122.040 368.350 123.440 ;
        RECT 4.000 121.400 368.350 122.040 ;
        RECT 4.000 120.000 367.950 121.400 ;
        RECT 4.000 115.280 368.350 120.000 ;
        RECT 4.000 114.600 367.950 115.280 ;
        RECT 4.400 113.880 367.950 114.600 ;
        RECT 4.400 113.200 368.350 113.880 ;
        RECT 4.000 109.840 368.350 113.200 ;
        RECT 4.000 108.440 367.950 109.840 ;
        RECT 4.000 106.440 368.350 108.440 ;
        RECT 4.400 105.040 368.350 106.440 ;
        RECT 4.000 104.400 368.350 105.040 ;
        RECT 4.000 103.000 367.950 104.400 ;
        RECT 4.000 98.960 368.350 103.000 ;
        RECT 4.000 97.600 367.950 98.960 ;
        RECT 4.400 97.560 367.950 97.600 ;
        RECT 4.400 96.200 368.350 97.560 ;
        RECT 4.000 92.840 368.350 96.200 ;
        RECT 4.000 91.440 367.950 92.840 ;
        RECT 4.000 89.440 368.350 91.440 ;
        RECT 4.400 88.040 368.350 89.440 ;
        RECT 4.000 87.400 368.350 88.040 ;
        RECT 4.000 86.000 367.950 87.400 ;
        RECT 4.000 81.960 368.350 86.000 ;
        RECT 4.000 81.280 367.950 81.960 ;
        RECT 4.400 80.560 367.950 81.280 ;
        RECT 4.400 79.880 368.350 80.560 ;
        RECT 4.000 76.520 368.350 79.880 ;
        RECT 4.000 75.120 367.950 76.520 ;
        RECT 4.000 72.440 368.350 75.120 ;
        RECT 4.400 71.040 368.350 72.440 ;
        RECT 4.000 70.400 368.350 71.040 ;
        RECT 4.000 69.000 367.950 70.400 ;
        RECT 4.000 64.960 368.350 69.000 ;
        RECT 4.000 64.280 367.950 64.960 ;
        RECT 4.400 63.560 367.950 64.280 ;
        RECT 4.400 62.880 368.350 63.560 ;
        RECT 4.000 59.520 368.350 62.880 ;
        RECT 4.000 58.120 367.950 59.520 ;
        RECT 4.000 55.440 368.350 58.120 ;
        RECT 4.400 54.080 368.350 55.440 ;
        RECT 4.400 54.040 367.950 54.080 ;
        RECT 4.000 52.680 367.950 54.040 ;
        RECT 4.000 47.960 368.350 52.680 ;
        RECT 4.000 47.280 367.950 47.960 ;
        RECT 4.400 46.560 367.950 47.280 ;
        RECT 4.400 45.880 368.350 46.560 ;
        RECT 4.000 42.520 368.350 45.880 ;
        RECT 4.000 41.120 367.950 42.520 ;
        RECT 4.000 38.440 368.350 41.120 ;
        RECT 4.400 37.080 368.350 38.440 ;
        RECT 4.400 37.040 367.950 37.080 ;
        RECT 4.000 35.680 367.950 37.040 ;
        RECT 4.000 31.640 368.350 35.680 ;
        RECT 4.000 30.280 367.950 31.640 ;
        RECT 4.400 30.240 367.950 30.280 ;
        RECT 4.400 28.880 368.350 30.240 ;
        RECT 4.000 25.520 368.350 28.880 ;
        RECT 4.000 24.120 367.950 25.520 ;
        RECT 4.000 21.440 368.350 24.120 ;
        RECT 4.400 20.080 368.350 21.440 ;
        RECT 4.400 20.040 367.950 20.080 ;
        RECT 4.000 18.680 367.950 20.040 ;
        RECT 4.000 14.640 368.350 18.680 ;
        RECT 4.000 13.280 367.950 14.640 ;
        RECT 4.400 13.240 367.950 13.280 ;
        RECT 4.400 11.880 368.350 13.240 ;
        RECT 4.000 9.200 368.350 11.880 ;
        RECT 4.000 7.800 367.950 9.200 ;
        RECT 4.000 5.120 368.350 7.800 ;
        RECT 4.400 3.760 368.350 5.120 ;
        RECT 4.400 3.720 367.950 3.760 ;
        RECT 4.000 2.895 367.950 3.720 ;
      LAYER met4 ;
        RECT 10.415 15.135 20.640 384.705 ;
        RECT 23.040 15.135 97.440 384.705 ;
        RECT 99.840 15.135 174.240 384.705 ;
        RECT 176.640 15.135 251.040 384.705 ;
        RECT 253.440 15.135 327.840 384.705 ;
        RECT 330.240 15.135 357.585 384.705 ;
  END
END wrapped_hack_soc_dffram
END LIBRARY

