magic
tech sky130A
magscale 1 2
timestamp 1646327704
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 251818 700680 251824 700732
rect 251876 700720 251882 700732
rect 267642 700720 267648 700732
rect 251876 700692 267648 700720
rect 251876 700680 251882 700692
rect 267642 700680 267648 700692
rect 267700 700680 267706 700732
rect 195790 700612 195796 700664
rect 195848 700652 195854 700664
rect 300118 700652 300124 700664
rect 195848 700624 300124 700652
rect 195848 700612 195854 700624
rect 300118 700612 300124 700624
rect 300176 700612 300182 700664
rect 198642 700544 198648 700596
rect 198700 700584 198706 700596
rect 332502 700584 332508 700596
rect 198700 700556 332508 700584
rect 198700 700544 198706 700556
rect 332502 700544 332508 700556
rect 332560 700544 332566 700596
rect 235534 700476 235540 700528
rect 235592 700516 235598 700528
rect 413646 700516 413652 700528
rect 235592 700488 413652 700516
rect 235592 700476 235598 700488
rect 413646 700476 413652 700488
rect 413704 700476 413710 700528
rect 197262 700408 197268 700460
rect 197320 700448 197326 700460
rect 397454 700448 397460 700460
rect 197320 700420 397460 700448
rect 197320 700408 197326 700420
rect 397454 700408 397460 700420
rect 397512 700408 397518 700460
rect 234614 700340 234620 700392
rect 234672 700380 234678 700392
rect 478506 700380 478512 700392
rect 234672 700352 478512 700380
rect 234672 700340 234678 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 529198 700340 529204 700392
rect 529256 700380 529262 700392
rect 559650 700380 559656 700392
rect 529256 700352 559656 700380
rect 529256 700340 529262 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 40494 700272 40500 700324
rect 40552 700312 40558 700324
rect 50338 700312 50344 700324
rect 40552 700284 50344 700312
rect 40552 700272 40558 700284
rect 50338 700272 50344 700284
rect 50396 700272 50402 700324
rect 195882 700272 195888 700324
rect 195940 700312 195946 700324
rect 218974 700312 218980 700324
rect 195940 700284 218980 700312
rect 195940 700272 195946 700284
rect 218974 700272 218980 700284
rect 219032 700272 219038 700324
rect 247678 700272 247684 700324
rect 247736 700312 247742 700324
rect 543458 700312 543464 700324
rect 247736 700284 543464 700312
rect 247736 700272 247742 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 154114 700068 154120 700120
rect 154172 700108 154178 700120
rect 155218 700108 155224 700120
rect 154172 700080 155224 700108
rect 154172 700068 154178 700080
rect 155218 700068 155224 700080
rect 155276 700068 155282 700120
rect 105446 699728 105452 699780
rect 105504 699768 105510 699780
rect 108298 699768 108304 699780
rect 105504 699740 108304 699768
rect 105504 699728 105510 699740
rect 108298 699728 108304 699740
rect 108356 699728 108362 699780
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 26878 699700 26884 699712
rect 24360 699672 26884 699700
rect 24360 699660 24366 699672
rect 26878 699660 26884 699672
rect 26936 699660 26942 699712
rect 347038 699660 347044 699712
rect 347096 699700 347102 699712
rect 348786 699700 348792 699712
rect 347096 699672 348792 699700
rect 347096 699660 347102 699672
rect 348786 699660 348792 699672
rect 348844 699660 348850 699712
rect 422938 699660 422944 699712
rect 422996 699700 423002 699712
rect 429838 699700 429844 699712
rect 422996 699672 429844 699700
rect 422996 699660 423002 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 526438 699660 526444 699712
rect 526496 699700 526502 699712
rect 527174 699700 527180 699712
rect 526496 699672 527180 699700
rect 526496 699660 526502 699672
rect 527174 699660 527180 699672
rect 527232 699660 527238 699712
rect 212902 696940 212908 696992
rect 212960 696980 212966 696992
rect 580166 696980 580172 696992
rect 212960 696952 580172 696980
rect 212960 696940 212966 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 253198 696192 253204 696244
rect 253256 696232 253262 696244
rect 283834 696232 283840 696244
rect 253256 696204 283840 696232
rect 253256 696192 253262 696204
rect 283834 696192 283840 696204
rect 283892 696192 283898 696244
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 246206 683176 246212 683188
rect 3476 683148 246212 683176
rect 3476 683136 3482 683148
rect 246206 683136 246212 683148
rect 246264 683136 246270 683188
rect 295978 683136 295984 683188
rect 296036 683176 296042 683188
rect 580166 683176 580172 683188
rect 296036 683148 580172 683176
rect 296036 683136 296042 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 156598 670732 156604 670744
rect 3568 670704 156604 670732
rect 3568 670692 3574 670704
rect 156598 670692 156604 670704
rect 156656 670692 156662 670744
rect 223022 670692 223028 670744
rect 223080 670732 223086 670744
rect 580166 670732 580172 670744
rect 223080 670704 580172 670732
rect 223080 670692 223086 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 233878 656928 233884 656940
rect 3476 656900 233884 656928
rect 3476 656888 3482 656900
rect 233878 656888 233884 656900
rect 233936 656888 233942 656940
rect 249058 643084 249064 643136
rect 249116 643124 249122 643136
rect 580166 643124 580172 643136
rect 249116 643096 580172 643124
rect 249116 643084 249122 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 28258 632108 28264 632120
rect 3476 632080 28264 632108
rect 3476 632068 3482 632080
rect 28258 632068 28264 632080
rect 28316 632068 28322 632120
rect 260098 630640 260104 630692
rect 260156 630680 260162 630692
rect 580166 630680 580172 630692
rect 260156 630652 580172 630680
rect 260156 630640 260162 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 29638 618304 29644 618316
rect 3200 618276 29644 618304
rect 3200 618264 3206 618276
rect 29638 618264 29644 618276
rect 29696 618264 29702 618316
rect 255958 616836 255964 616888
rect 256016 616876 256022 616888
rect 580166 616876 580172 616888
rect 256016 616848 580172 616876
rect 256016 616836 256022 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 224218 605860 224224 605872
rect 3292 605832 224224 605860
rect 3292 605820 3298 605832
rect 224218 605820 224224 605832
rect 224276 605820 224282 605872
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 240778 579680 240784 579692
rect 3384 579652 240784 579680
rect 3384 579640 3390 579652
rect 240778 579640 240784 579652
rect 240836 579640 240842 579692
rect 225966 563048 225972 563100
rect 226024 563088 226030 563100
rect 579890 563088 579896 563100
rect 226024 563060 579896 563088
rect 226024 563048 226030 563060
rect 579890 563048 579896 563060
rect 579948 563048 579954 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 25498 553432 25504 553444
rect 3384 553404 25504 553432
rect 3384 553392 3390 553404
rect 25498 553392 25504 553404
rect 25556 553392 25562 553444
rect 250438 536800 250444 536852
rect 250496 536840 250502 536852
rect 580166 536840 580172 536852
rect 250496 536812 580172 536840
rect 250496 536800 250502 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 10318 527184 10324 527196
rect 3016 527156 10324 527184
rect 3016 527144 3022 527156
rect 10318 527144 10324 527156
rect 10376 527144 10382 527196
rect 294598 524424 294604 524476
rect 294656 524464 294662 524476
rect 580166 524464 580172 524476
rect 294656 524436 580172 524464
rect 294656 524424 294662 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 198550 510620 198556 510672
rect 198608 510660 198614 510672
rect 580166 510660 580172 510672
rect 198608 510632 580172 510660
rect 198608 510620 198614 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3326 500964 3332 501016
rect 3384 501004 3390 501016
rect 244918 501004 244924 501016
rect 3384 500976 244924 501004
rect 3384 500964 3390 500976
rect 244918 500964 244924 500976
rect 244976 500964 244982 501016
rect 286318 484372 286324 484424
rect 286376 484412 286382 484424
rect 580166 484412 580172 484424
rect 286376 484384 580172 484412
rect 286376 484372 286382 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3050 474716 3056 474768
rect 3108 474756 3114 474768
rect 86218 474756 86224 474768
rect 3108 474728 86224 474756
rect 3108 474716 3114 474728
rect 86218 474716 86224 474728
rect 86276 474716 86282 474768
rect 258718 470568 258724 470620
rect 258776 470608 258782 470620
rect 580166 470608 580172 470620
rect 258776 470580 580172 470608
rect 258776 470568 258782 470580
rect 580166 470568 580172 470580
rect 580224 470568 580230 470620
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 175918 462380 175924 462392
rect 3384 462352 175924 462380
rect 3384 462340 3390 462352
rect 175918 462340 175924 462352
rect 175976 462340 175982 462392
rect 197170 456764 197176 456816
rect 197228 456804 197234 456816
rect 580166 456804 580172 456816
rect 197228 456776 580172 456804
rect 197228 456764 197234 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3326 448536 3332 448588
rect 3384 448576 3390 448588
rect 204898 448576 204904 448588
rect 3384 448548 204904 448576
rect 3384 448536 3390 448548
rect 204898 448536 204904 448548
rect 204956 448536 204962 448588
rect 251910 430584 251916 430636
rect 251968 430624 251974 430636
rect 580166 430624 580172 430636
rect 251968 430596 580172 430624
rect 251968 430584 251974 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3142 422288 3148 422340
rect 3200 422328 3206 422340
rect 15838 422328 15844 422340
rect 3200 422300 15844 422328
rect 3200 422288 3206 422300
rect 15838 422288 15844 422300
rect 15896 422288 15902 422340
rect 213454 418140 213460 418192
rect 213512 418180 213518 418192
rect 580166 418180 580172 418192
rect 213512 418152 580172 418180
rect 213512 418140 213518 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 200114 404336 200120 404388
rect 200172 404376 200178 404388
rect 579982 404376 579988 404388
rect 200172 404348 579988 404376
rect 200172 404336 200178 404348
rect 579982 404336 579988 404348
rect 580040 404336 580046 404388
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 195330 397508 195336 397520
rect 3384 397480 195336 397508
rect 3384 397468 3390 397480
rect 195330 397468 195336 397480
rect 195388 397468 195394 397520
rect 305638 378156 305644 378208
rect 305696 378196 305702 378208
rect 580166 378196 580172 378208
rect 305696 378168 580172 378196
rect 305696 378156 305702 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 196710 371260 196716 371272
rect 3384 371232 196716 371260
rect 3384 371220 3390 371232
rect 196710 371220 196716 371232
rect 196768 371220 196774 371272
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 226978 357456 226984 357468
rect 3384 357428 226984 357456
rect 3384 357416 3390 357428
rect 226978 357416 226984 357428
rect 227036 357416 227042 357468
rect 209958 351908 209964 351960
rect 210016 351948 210022 351960
rect 580166 351948 580172 351960
rect 210016 351920 580172 351948
rect 210016 351908 210022 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 232498 345080 232504 345092
rect 3384 345052 232504 345080
rect 3384 345040 3390 345052
rect 232498 345040 232504 345052
rect 232556 345040 232562 345092
rect 250622 324300 250628 324352
rect 250680 324340 250686 324352
rect 579614 324340 579620 324352
rect 250680 324312 579620 324340
rect 250680 324300 250686 324312
rect 579614 324300 579620 324312
rect 579672 324300 579678 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 214558 318832 214564 318844
rect 3384 318804 214564 318832
rect 3384 318792 3390 318804
rect 214558 318792 214564 318804
rect 214616 318792 214622 318844
rect 234706 312536 234712 312588
rect 234764 312576 234770 312588
rect 246850 312576 246856 312588
rect 234764 312548 246856 312576
rect 234764 312536 234770 312548
rect 246850 312536 246856 312548
rect 246908 312536 246914 312588
rect 316678 311856 316684 311908
rect 316736 311896 316742 311908
rect 580166 311896 580172 311908
rect 316736 311868 580172 311896
rect 316736 311856 316742 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 3050 298732 3056 298784
rect 3108 298772 3114 298784
rect 244366 298772 244372 298784
rect 3108 298744 244372 298772
rect 3108 298732 3114 298744
rect 244366 298732 244372 298744
rect 244424 298732 244430 298784
rect 250714 298120 250720 298172
rect 250772 298160 250778 298172
rect 580166 298160 580172 298172
rect 250772 298132 580172 298160
rect 250772 298120 250778 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 88334 297372 88340 297424
rect 88392 297412 88398 297424
rect 232774 297412 232780 297424
rect 88392 297384 232780 297412
rect 88392 297372 88398 297384
rect 232774 297372 232780 297384
rect 232832 297372 232838 297424
rect 218606 295944 218612 295996
rect 218664 295984 218670 295996
rect 347038 295984 347044 295996
rect 218664 295956 347044 295984
rect 218664 295944 218670 295956
rect 347038 295944 347044 295956
rect 347096 295944 347102 295996
rect 71774 294584 71780 294636
rect 71832 294624 71838 294636
rect 240502 294624 240508 294636
rect 71832 294596 240508 294624
rect 71832 294584 71838 294596
rect 240502 294584 240508 294596
rect 240560 294584 240566 294636
rect 201494 293224 201500 293276
rect 201552 293264 201558 293276
rect 244274 293264 244280 293276
rect 201552 293236 244280 293264
rect 201552 293224 201558 293236
rect 244274 293224 244280 293236
rect 244332 293224 244338 293276
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 11698 292584 11704 292596
rect 3384 292556 11704 292584
rect 3384 292544 3390 292556
rect 11698 292544 11704 292556
rect 11756 292544 11762 292596
rect 15838 291796 15844 291848
rect 15896 291836 15902 291848
rect 209038 291836 209044 291848
rect 15896 291808 209044 291836
rect 15896 291796 15902 291808
rect 209038 291796 209044 291808
rect 209096 291796 209102 291848
rect 214558 291796 214564 291848
rect 214616 291836 214622 291848
rect 241422 291836 241428 291848
rect 214616 291808 241428 291836
rect 214616 291796 214622 291808
rect 241422 291796 241428 291808
rect 241480 291796 241486 291848
rect 233878 289144 233884 289196
rect 233936 289184 233942 289196
rect 245654 289184 245660 289196
rect 233936 289156 245660 289184
rect 233936 289144 233942 289156
rect 245654 289144 245660 289156
rect 245712 289144 245718 289196
rect 198366 289076 198372 289128
rect 198424 289116 198430 289128
rect 422938 289116 422944 289128
rect 198424 289088 422944 289116
rect 198424 289076 198430 289088
rect 422938 289076 422944 289088
rect 422996 289076 423002 289128
rect 224494 288736 224500 288788
rect 224552 288776 224558 288788
rect 251358 288776 251364 288788
rect 224552 288748 251364 288776
rect 224552 288736 224558 288748
rect 251358 288736 251364 288748
rect 251416 288736 251422 288788
rect 222470 288668 222476 288720
rect 222528 288708 222534 288720
rect 250070 288708 250076 288720
rect 222528 288680 250076 288708
rect 222528 288668 222534 288680
rect 250070 288668 250076 288680
rect 250128 288668 250134 288720
rect 216214 288600 216220 288652
rect 216272 288640 216278 288652
rect 247126 288640 247132 288652
rect 216272 288612 247132 288640
rect 216272 288600 216278 288612
rect 247126 288600 247132 288612
rect 247184 288600 247190 288652
rect 220078 288532 220084 288584
rect 220136 288572 220142 288584
rect 251266 288572 251272 288584
rect 220136 288544 251272 288572
rect 220136 288532 220142 288544
rect 251266 288532 251272 288544
rect 251324 288532 251330 288584
rect 214374 288464 214380 288516
rect 214432 288504 214438 288516
rect 249886 288504 249892 288516
rect 214432 288476 249892 288504
rect 214432 288464 214438 288476
rect 249886 288464 249892 288476
rect 249944 288464 249950 288516
rect 235166 288396 235172 288448
rect 235224 288436 235230 288448
rect 287054 288436 287060 288448
rect 235224 288408 287060 288436
rect 235224 288396 235230 288408
rect 287054 288396 287060 288408
rect 287112 288396 287118 288448
rect 204898 288328 204904 288380
rect 204956 288368 204962 288380
rect 208118 288368 208124 288380
rect 204956 288340 208124 288368
rect 204956 288328 204962 288340
rect 208118 288328 208124 288340
rect 208176 288328 208182 288380
rect 224218 288328 224224 288380
rect 224276 288368 224282 288380
rect 225414 288368 225420 288380
rect 224276 288340 225420 288368
rect 224276 288328 224282 288340
rect 225414 288328 225420 288340
rect 225472 288328 225478 288380
rect 226978 288328 226984 288380
rect 227036 288368 227042 288380
rect 228358 288368 228364 288380
rect 227036 288340 228364 288368
rect 227036 288328 227042 288340
rect 228358 288328 228364 288340
rect 228416 288328 228422 288380
rect 201310 287920 201316 287972
rect 201368 287960 201374 287972
rect 287330 287960 287336 287972
rect 201368 287932 287336 287960
rect 201368 287920 201374 287932
rect 287330 287920 287336 287932
rect 287388 287920 287394 287972
rect 202230 287852 202236 287904
rect 202288 287892 202294 287904
rect 289814 287892 289820 287904
rect 202288 287864 289820 287892
rect 202288 287852 202294 287864
rect 289814 287852 289820 287864
rect 289872 287852 289878 287904
rect 220630 287784 220636 287836
rect 220688 287824 220694 287836
rect 247218 287824 247224 287836
rect 220688 287796 247224 287824
rect 220688 287784 220694 287796
rect 247218 287784 247224 287796
rect 247276 287784 247282 287836
rect 86218 287716 86224 287768
rect 86276 287756 86282 287768
rect 246114 287756 246120 287768
rect 86276 287728 246120 287756
rect 86276 287716 86282 287728
rect 246114 287716 246120 287728
rect 246172 287716 246178 287768
rect 26878 287648 26884 287700
rect 26936 287688 26942 287700
rect 218238 287688 218244 287700
rect 26936 287660 218244 287688
rect 26936 287648 26942 287660
rect 218238 287648 218244 287660
rect 218296 287648 218302 287700
rect 232498 287648 232504 287700
rect 232556 287688 232562 287700
rect 243630 287688 243636 287700
rect 232556 287660 243636 287688
rect 232556 287648 232562 287660
rect 243630 287648 243636 287660
rect 243688 287648 243694 287700
rect 231302 287580 231308 287632
rect 231360 287620 231366 287632
rect 251174 287620 251180 287632
rect 231360 287592 251180 287620
rect 231360 287580 231366 287592
rect 251174 287580 251180 287592
rect 251232 287580 251238 287632
rect 217318 287512 217324 287564
rect 217376 287552 217382 287564
rect 248598 287552 248604 287564
rect 217376 287524 248604 287552
rect 217376 287512 217382 287524
rect 248598 287512 248604 287524
rect 248656 287512 248662 287564
rect 216766 287444 216772 287496
rect 216824 287484 216830 287496
rect 248690 287484 248696 287496
rect 216824 287456 248696 287484
rect 216824 287444 216830 287456
rect 248690 287444 248696 287456
rect 248748 287444 248754 287496
rect 239582 287376 239588 287428
rect 239640 287416 239646 287428
rect 291194 287416 291200 287428
rect 239640 287388 291200 287416
rect 239640 287376 239646 287388
rect 291194 287376 291200 287388
rect 291252 287376 291258 287428
rect 232222 287308 232228 287360
rect 232280 287348 232286 287360
rect 292574 287348 292580 287360
rect 232280 287320 292580 287348
rect 232280 287308 232286 287320
rect 292574 287308 292580 287320
rect 292632 287308 292638 287360
rect 222102 287240 222108 287292
rect 222160 287280 222166 287292
rect 287146 287280 287152 287292
rect 222160 287252 287152 287280
rect 222160 287240 222166 287252
rect 287146 287240 287152 287252
rect 287204 287240 287210 287292
rect 211982 287172 211988 287224
rect 212040 287212 212046 287224
rect 287238 287212 287244 287224
rect 212040 287184 287244 287212
rect 212040 287172 212046 287184
rect 287238 287172 287244 287184
rect 287296 287172 287302 287224
rect 230750 287104 230756 287156
rect 230808 287144 230814 287156
rect 249978 287144 249984 287156
rect 230808 287116 249984 287144
rect 230808 287104 230814 287116
rect 249978 287104 249984 287116
rect 250036 287104 250042 287156
rect 229278 287036 229284 287088
rect 229336 287076 229342 287088
rect 249794 287076 249800 287088
rect 229336 287048 249800 287076
rect 229336 287036 229342 287048
rect 249794 287036 249800 287048
rect 249852 287036 249858 287088
rect 209406 286560 209412 286612
rect 209464 286600 209470 286612
rect 280890 286600 280896 286612
rect 209464 286572 280896 286600
rect 209464 286560 209470 286572
rect 280890 286560 280896 286572
rect 280948 286560 280954 286612
rect 219158 286492 219164 286544
rect 219216 286532 219222 286544
rect 248782 286532 248788 286544
rect 219216 286504 248788 286532
rect 219216 286492 219222 286504
rect 248782 286492 248788 286504
rect 248840 286492 248846 286544
rect 208486 286424 208492 286476
rect 208544 286464 208550 286476
rect 283190 286464 283196 286476
rect 208544 286436 283196 286464
rect 208544 286424 208550 286436
rect 283190 286424 283196 286436
rect 283248 286424 283254 286476
rect 156598 286356 156604 286408
rect 156656 286396 156662 286408
rect 202782 286396 202788 286408
rect 156656 286368 202788 286396
rect 156656 286356 156662 286368
rect 202782 286356 202788 286368
rect 202840 286356 202846 286408
rect 207566 286356 207572 286408
rect 207624 286396 207630 286408
rect 283650 286396 283656 286408
rect 207624 286368 283656 286396
rect 207624 286356 207630 286368
rect 283650 286356 283656 286368
rect 283708 286356 283714 286408
rect 155218 286288 155224 286340
rect 155276 286328 155282 286340
rect 204254 286328 204260 286340
rect 155276 286300 204260 286328
rect 155276 286288 155282 286300
rect 204254 286288 204260 286300
rect 204312 286288 204318 286340
rect 215294 286288 215300 286340
rect 215352 286328 215358 286340
rect 248506 286328 248512 286340
rect 215352 286300 248512 286328
rect 215352 286288 215358 286300
rect 248506 286288 248512 286300
rect 248564 286288 248570 286340
rect 210878 286220 210884 286272
rect 210936 286260 210942 286272
rect 247034 286260 247040 286272
rect 210936 286232 247040 286260
rect 210936 286220 210942 286232
rect 247034 286220 247040 286232
rect 247092 286220 247098 286272
rect 195422 286152 195428 286204
rect 195480 286192 195486 286204
rect 207014 286192 207020 286204
rect 195480 286164 207020 286192
rect 195480 286152 195486 286164
rect 207014 286152 207020 286164
rect 207072 286152 207078 286204
rect 236086 286152 236092 286204
rect 236144 286192 236150 286204
rect 278038 286192 278044 286204
rect 236144 286164 278044 286192
rect 236144 286152 236150 286164
rect 278038 286152 278044 286164
rect 278096 286152 278102 286204
rect 195606 286084 195612 286136
rect 195664 286124 195670 286136
rect 203702 286124 203708 286136
rect 195664 286096 203708 286124
rect 195664 286084 195670 286096
rect 203702 286084 203708 286096
rect 203760 286084 203766 286136
rect 205174 286084 205180 286136
rect 205232 286124 205238 286136
rect 247770 286124 247776 286136
rect 205232 286096 247776 286124
rect 205232 286084 205238 286096
rect 247770 286084 247776 286096
rect 247828 286084 247834 286136
rect 3694 286016 3700 286068
rect 3752 286056 3758 286068
rect 206094 286056 206100 286068
rect 3752 286028 206100 286056
rect 3752 286016 3758 286028
rect 206094 286016 206100 286028
rect 206152 286016 206158 286068
rect 237558 286016 237564 286068
rect 237616 286056 237622 286068
rect 285858 286056 285864 286068
rect 237616 286028 285864 286056
rect 237616 286016 237622 286028
rect 285858 286016 285864 286028
rect 285916 286016 285922 286068
rect 197078 285948 197084 286000
rect 197136 285988 197142 286000
rect 217686 285988 217692 286000
rect 197136 285960 217692 285988
rect 197136 285948 197142 285960
rect 217686 285948 217692 285960
rect 217744 285948 217750 286000
rect 228910 285948 228916 286000
rect 228968 285988 228974 286000
rect 280798 285988 280804 286000
rect 228968 285960 280804 285988
rect 228968 285948 228974 285960
rect 280798 285948 280804 285960
rect 280856 285948 280862 286000
rect 194410 285880 194416 285932
rect 194468 285920 194474 285932
rect 204622 285920 204628 285932
rect 194468 285892 204628 285920
rect 194468 285880 194474 285892
rect 204622 285880 204628 285892
rect 204680 285880 204686 285932
rect 211430 285880 211436 285932
rect 211488 285920 211494 285932
rect 265618 285920 265624 285932
rect 211488 285892 265624 285920
rect 211488 285880 211494 285892
rect 265618 285880 265624 285892
rect 265676 285880 265682 285932
rect 196986 285812 196992 285864
rect 197044 285852 197050 285864
rect 203150 285852 203156 285864
rect 197044 285824 203156 285852
rect 197044 285812 197050 285824
rect 203150 285812 203156 285824
rect 203208 285812 203214 285864
rect 234246 285812 234252 285864
rect 234304 285852 234310 285864
rect 244090 285852 244096 285864
rect 234304 285824 244096 285852
rect 234304 285812 234310 285824
rect 244090 285812 244096 285824
rect 244148 285812 244154 285864
rect 196894 285744 196900 285796
rect 196952 285784 196958 285796
rect 210510 285784 210516 285796
rect 196952 285756 210516 285784
rect 196952 285744 196958 285756
rect 210510 285744 210516 285756
rect 210568 285744 210574 285796
rect 227806 285744 227812 285796
rect 227864 285784 227870 285796
rect 243906 285784 243912 285796
rect 227864 285756 243912 285784
rect 227864 285744 227870 285756
rect 243906 285744 243912 285756
rect 243964 285744 243970 285796
rect 195514 285676 195520 285728
rect 195572 285716 195578 285728
rect 205542 285716 205548 285728
rect 195572 285688 205548 285716
rect 195572 285676 195578 285688
rect 205542 285676 205548 285688
rect 205600 285676 205606 285728
rect 226518 285676 226524 285728
rect 226576 285716 226582 285728
rect 250530 285716 250536 285728
rect 226576 285688 250536 285716
rect 226576 285676 226582 285688
rect 250530 285676 250536 285688
rect 250588 285676 250594 285728
rect 196618 285200 196624 285252
rect 196676 285240 196682 285252
rect 242894 285240 242900 285252
rect 196676 285212 242900 285240
rect 196676 285200 196682 285212
rect 242894 285200 242900 285212
rect 242952 285200 242958 285252
rect 229830 285132 229836 285184
rect 229888 285172 229894 285184
rect 250162 285172 250168 285184
rect 229888 285144 250168 285172
rect 229888 285132 229894 285144
rect 250162 285132 250168 285144
rect 250220 285132 250226 285184
rect 201678 285064 201684 285116
rect 201736 285104 201742 285116
rect 249150 285104 249156 285116
rect 201736 285076 249156 285104
rect 201736 285064 201742 285076
rect 249150 285064 249156 285076
rect 249208 285064 249214 285116
rect 214742 284996 214748 285048
rect 214800 285036 214806 285048
rect 256050 285036 256056 285048
rect 214800 285008 256056 285036
rect 214800 284996 214806 285008
rect 256050 284996 256056 285008
rect 256108 284996 256114 285048
rect 231670 284928 231676 284980
rect 231728 284968 231734 284980
rect 284294 284968 284300 284980
rect 231728 284940 284300 284968
rect 231728 284928 231734 284940
rect 284294 284928 284300 284940
rect 284352 284928 284358 284980
rect 223574 284860 223580 284912
rect 223632 284900 223638 284912
rect 247310 284900 247316 284912
rect 223632 284872 247316 284900
rect 223632 284860 223638 284872
rect 247310 284860 247316 284872
rect 247368 284860 247374 284912
rect 225046 284792 225052 284844
rect 225104 284832 225110 284844
rect 251542 284832 251548 284844
rect 225104 284804 251548 284832
rect 225104 284792 225110 284804
rect 251542 284792 251548 284804
rect 251600 284792 251606 284844
rect 212350 284724 212356 284776
rect 212408 284764 212414 284776
rect 243998 284764 244004 284776
rect 212408 284736 244004 284764
rect 212408 284724 212414 284736
rect 243998 284724 244004 284736
rect 244056 284724 244062 284776
rect 192478 284656 192484 284708
rect 192536 284696 192542 284708
rect 223942 284696 223948 284708
rect 192536 284668 223948 284696
rect 192536 284656 192542 284668
rect 223942 284656 223948 284668
rect 224000 284656 224006 284708
rect 238110 284656 238116 284708
rect 238168 284696 238174 284708
rect 283098 284696 283104 284708
rect 238168 284668 283104 284696
rect 238168 284656 238174 284668
rect 283098 284656 283104 284668
rect 283156 284656 283162 284708
rect 195238 284588 195244 284640
rect 195296 284628 195302 284640
rect 230382 284628 230388 284640
rect 195296 284600 230388 284628
rect 195296 284588 195302 284600
rect 230382 284588 230388 284600
rect 230440 284588 230446 284640
rect 241974 284588 241980 284640
rect 242032 284628 242038 284640
rect 288710 284628 288716 284640
rect 242032 284600 288716 284628
rect 242032 284588 242038 284600
rect 288710 284588 288716 284600
rect 288768 284588 288774 284640
rect 236638 284520 236644 284572
rect 236696 284560 236702 284572
rect 252002 284560 252008 284572
rect 236696 284532 252008 284560
rect 236696 284520 236702 284532
rect 252002 284520 252008 284532
rect 252060 284520 252066 284572
rect 239950 284452 239956 284504
rect 240008 284492 240014 284504
rect 289262 284492 289268 284504
rect 240008 284464 289268 284492
rect 240008 284452 240014 284464
rect 289262 284452 289268 284464
rect 289320 284452 289326 284504
rect 188338 284384 188344 284436
rect 188396 284424 188402 284436
rect 227438 284424 227444 284436
rect 188396 284396 227444 284424
rect 188396 284384 188402 284396
rect 227438 284384 227444 284396
rect 227496 284384 227502 284436
rect 233142 284384 233148 284436
rect 233200 284424 233206 284436
rect 249242 284424 249248 284436
rect 233200 284396 249248 284424
rect 233200 284384 233206 284396
rect 249242 284384 249248 284396
rect 249300 284384 249306 284436
rect 18598 284316 18604 284368
rect 18656 284356 18662 284368
rect 213822 284356 213828 284368
rect 18656 284328 213828 284356
rect 18656 284316 18662 284328
rect 213822 284316 213828 284328
rect 213880 284316 213886 284368
rect 240870 284316 240876 284368
rect 240928 284356 240934 284368
rect 298738 284356 298744 284368
rect 240928 284328 298744 284356
rect 240928 284316 240934 284328
rect 298738 284316 298744 284328
rect 298796 284316 298802 284368
rect 242618 284044 242624 284096
rect 242676 284084 242682 284096
rect 283742 284084 283748 284096
rect 242676 284056 283748 284084
rect 242676 284044 242682 284056
rect 283742 284044 283748 284056
rect 283800 284044 283806 284096
rect 238570 283976 238576 284028
rect 238628 284016 238634 284028
rect 251450 284016 251456 284028
rect 238628 283988 251456 284016
rect 238628 283976 238634 283988
rect 251450 283976 251456 283988
rect 251508 283976 251514 284028
rect 237282 283908 237288 283960
rect 237340 283948 237346 283960
rect 244458 283948 244464 283960
rect 237340 283920 244464 283948
rect 237340 283908 237346 283920
rect 244458 283908 244464 283920
rect 244516 283908 244522 283960
rect 243906 283840 243912 283892
rect 243964 283880 243970 283892
rect 282178 283880 282184 283892
rect 243964 283852 282184 283880
rect 243964 283840 243970 283852
rect 282178 283840 282184 283852
rect 282236 283840 282242 283892
rect 244090 283568 244096 283620
rect 244148 283608 244154 283620
rect 282362 283608 282368 283620
rect 244148 283580 282368 283608
rect 244148 283568 244154 283580
rect 282362 283568 282368 283580
rect 282420 283568 282426 283620
rect 245930 282820 245936 282872
rect 245988 282860 245994 282872
rect 305638 282860 305644 282872
rect 245988 282832 305644 282860
rect 245988 282820 245994 282832
rect 305638 282820 305644 282832
rect 305696 282820 305702 282872
rect 58618 281528 58624 281580
rect 58676 281568 58682 281580
rect 197354 281568 197360 281580
rect 58676 281540 197360 281568
rect 58676 281528 58682 281540
rect 197354 281528 197360 281540
rect 197412 281528 197418 281580
rect 245654 280236 245660 280288
rect 245712 280276 245718 280288
rect 287422 280276 287428 280288
rect 245712 280248 287428 280276
rect 245712 280236 245718 280248
rect 287422 280236 287428 280248
rect 287480 280236 287486 280288
rect 193122 280168 193128 280220
rect 193180 280208 193186 280220
rect 197354 280208 197360 280220
rect 193180 280180 197360 280208
rect 193180 280168 193186 280180
rect 197354 280168 197360 280180
rect 197412 280168 197418 280220
rect 245930 280168 245936 280220
rect 245988 280208 245994 280220
rect 289906 280208 289912 280220
rect 245988 280180 289912 280208
rect 245988 280168 245994 280180
rect 289906 280168 289912 280180
rect 289964 280168 289970 280220
rect 193030 278740 193036 278792
rect 193088 278780 193094 278792
rect 197354 278780 197360 278792
rect 193088 278752 197360 278780
rect 193088 278740 193094 278752
rect 197354 278740 197360 278752
rect 197412 278740 197418 278792
rect 245654 278740 245660 278792
rect 245712 278780 245718 278792
rect 454678 278780 454684 278792
rect 245712 278752 454684 278780
rect 245712 278740 245718 278752
rect 454678 278740 454684 278752
rect 454736 278740 454742 278792
rect 194318 276020 194324 276072
rect 194376 276060 194382 276072
rect 197446 276060 197452 276072
rect 194376 276032 197452 276060
rect 194376 276020 194382 276032
rect 197446 276020 197452 276032
rect 197504 276020 197510 276072
rect 29638 275952 29644 276004
rect 29696 275992 29702 276004
rect 197354 275992 197360 276004
rect 29696 275964 197360 275992
rect 29696 275952 29702 275964
rect 197354 275952 197360 275964
rect 197412 275952 197418 276004
rect 246114 275952 246120 276004
rect 246172 275992 246178 276004
rect 526438 275992 526444 276004
rect 246172 275964 526444 275992
rect 246172 275952 246178 275964
rect 526438 275952 526444 275964
rect 526496 275952 526502 276004
rect 245746 275884 245752 275936
rect 245804 275924 245810 275936
rect 258718 275924 258724 275936
rect 245804 275896 258724 275924
rect 245804 275884 245810 275896
rect 258718 275884 258724 275896
rect 258776 275884 258782 275936
rect 245746 273232 245752 273284
rect 245804 273272 245810 273284
rect 285766 273272 285772 273284
rect 245804 273244 285772 273272
rect 245804 273232 245810 273244
rect 285766 273232 285772 273244
rect 285824 273232 285830 273284
rect 169754 273164 169760 273216
rect 169812 273204 169818 273216
rect 197354 273204 197360 273216
rect 169812 273176 197360 273204
rect 169812 273164 169818 273176
rect 197354 273164 197360 273176
rect 197412 273164 197418 273216
rect 245746 271940 245752 271992
rect 245804 271980 245810 271992
rect 288526 271980 288532 271992
rect 245804 271952 288532 271980
rect 245804 271940 245810 271952
rect 288526 271940 288532 271952
rect 288584 271940 288590 271992
rect 194502 271872 194508 271924
rect 194560 271912 194566 271924
rect 197446 271912 197452 271924
rect 194560 271884 197452 271912
rect 194560 271872 194566 271884
rect 197446 271872 197452 271884
rect 197504 271872 197510 271924
rect 258718 271872 258724 271924
rect 258776 271912 258782 271924
rect 580166 271912 580172 271924
rect 258776 271884 580172 271912
rect 258776 271872 258782 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 15838 269084 15844 269136
rect 15896 269124 15902 269136
rect 197354 269124 197360 269136
rect 15896 269096 197360 269124
rect 15896 269084 15902 269096
rect 197354 269084 197360 269096
rect 197412 269084 197418 269136
rect 245746 269084 245752 269136
rect 245804 269124 245810 269136
rect 288618 269124 288624 269136
rect 245804 269096 288624 269124
rect 245804 269084 245810 269096
rect 288618 269084 288624 269096
rect 288676 269084 288682 269136
rect 3418 269016 3424 269068
rect 3476 269056 3482 269068
rect 197446 269056 197452 269068
rect 3476 269028 197452 269056
rect 3476 269016 3482 269028
rect 197446 269016 197452 269028
rect 197504 269016 197510 269068
rect 6914 268948 6920 269000
rect 6972 268988 6978 269000
rect 197354 268988 197360 269000
rect 6972 268960 197360 268988
rect 6972 268948 6978 268960
rect 197354 268948 197360 268960
rect 197412 268948 197418 269000
rect 245654 267792 245660 267844
rect 245712 267832 245718 267844
rect 291286 267832 291292 267844
rect 245712 267804 291292 267832
rect 245712 267792 245718 267804
rect 291286 267792 291292 267804
rect 291344 267792 291350 267844
rect 245746 267724 245752 267776
rect 245804 267764 245810 267776
rect 291930 267764 291936 267776
rect 245804 267736 291936 267764
rect 245804 267724 245810 267736
rect 291930 267724 291936 267736
rect 291988 267724 291994 267776
rect 28258 267656 28264 267708
rect 28316 267696 28322 267708
rect 197354 267696 197360 267708
rect 28316 267668 197360 267696
rect 28316 267656 28322 267668
rect 197354 267656 197360 267668
rect 197412 267656 197418 267708
rect 245654 266704 245660 266756
rect 245712 266744 245718 266756
rect 245930 266744 245936 266756
rect 245712 266716 245936 266744
rect 245712 266704 245718 266716
rect 245930 266704 245936 266716
rect 245988 266704 245994 266756
rect 3326 266568 3332 266620
rect 3384 266608 3390 266620
rect 7558 266608 7564 266620
rect 3384 266580 7564 266608
rect 3384 266568 3390 266580
rect 7558 266568 7564 266580
rect 7616 266568 7622 266620
rect 245746 266432 245752 266484
rect 245804 266472 245810 266484
rect 284386 266472 284392 266484
rect 245804 266444 284392 266472
rect 245804 266432 245810 266444
rect 284386 266432 284392 266444
rect 284444 266432 284450 266484
rect 192938 266364 192944 266416
rect 192996 266404 193002 266416
rect 197446 266404 197452 266416
rect 192996 266376 197452 266404
rect 192996 266364 193002 266376
rect 197446 266364 197452 266376
rect 197504 266364 197510 266416
rect 245930 266364 245936 266416
rect 245988 266404 245994 266416
rect 565078 266404 565084 266416
rect 245988 266376 565084 266404
rect 245988 266364 245994 266376
rect 565078 266364 565084 266376
rect 565136 266364 565142 266416
rect 246114 266296 246120 266348
rect 246172 266336 246178 266348
rect 316678 266336 316684 266348
rect 246172 266308 316684 266336
rect 246172 266296 246178 266308
rect 316678 266296 316684 266308
rect 316736 266296 316742 266348
rect 192846 265004 192852 265056
rect 192904 265044 192910 265056
rect 197354 265044 197360 265056
rect 192904 265016 197360 265044
rect 192904 265004 192910 265016
rect 197354 265004 197360 265016
rect 197412 265004 197418 265056
rect 17218 264936 17224 264988
rect 17276 264976 17282 264988
rect 197446 264976 197452 264988
rect 17276 264948 197452 264976
rect 17276 264936 17282 264948
rect 197446 264936 197452 264948
rect 197504 264936 197510 264988
rect 25498 264868 25504 264920
rect 25556 264908 25562 264920
rect 197354 264908 197360 264920
rect 25556 264880 197360 264908
rect 25556 264868 25562 264880
rect 197354 264868 197360 264880
rect 197412 264868 197418 264920
rect 196434 263576 196440 263628
rect 196492 263616 196498 263628
rect 197354 263616 197360 263628
rect 196492 263588 197360 263616
rect 196492 263576 196498 263588
rect 197354 263576 197360 263588
rect 197412 263576 197418 263628
rect 10318 262148 10324 262200
rect 10376 262188 10382 262200
rect 197354 262188 197360 262200
rect 10376 262160 197360 262188
rect 10376 262148 10382 262160
rect 197354 262148 197360 262160
rect 197412 262148 197418 262200
rect 245930 259428 245936 259480
rect 245988 259468 245994 259480
rect 286502 259468 286508 259480
rect 245988 259440 286508 259468
rect 245988 259428 245994 259440
rect 286502 259428 286508 259440
rect 286560 259428 286566 259480
rect 244090 259360 244096 259412
rect 244148 259400 244154 259412
rect 580166 259400 580172 259412
rect 244148 259372 580172 259400
rect 244148 259360 244154 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 245838 259292 245844 259344
rect 245896 259292 245902 259344
rect 245856 259072 245884 259292
rect 245838 259020 245844 259072
rect 245896 259020 245902 259072
rect 195146 258612 195152 258664
rect 195204 258652 195210 258664
rect 197446 258652 197452 258664
rect 195204 258624 197452 258652
rect 195204 258612 195210 258624
rect 197446 258612 197452 258624
rect 197504 258612 197510 258664
rect 246482 258136 246488 258188
rect 246540 258176 246546 258188
rect 288802 258176 288808 258188
rect 246540 258148 288808 258176
rect 246540 258136 246546 258148
rect 288802 258136 288808 258148
rect 288860 258136 288866 258188
rect 26878 258068 26884 258120
rect 26936 258108 26942 258120
rect 197354 258108 197360 258120
rect 26936 258080 197360 258108
rect 26936 258068 26942 258080
rect 197354 258068 197360 258080
rect 197412 258068 197418 258120
rect 245746 258068 245752 258120
rect 245804 258108 245810 258120
rect 292666 258108 292672 258120
rect 245804 258080 292672 258108
rect 245804 258068 245810 258080
rect 292666 258068 292672 258080
rect 292724 258068 292730 258120
rect 246206 256912 246212 256964
rect 246264 256952 246270 256964
rect 246482 256952 246488 256964
rect 246264 256924 246488 256952
rect 246264 256912 246270 256924
rect 246482 256912 246488 256924
rect 246540 256912 246546 256964
rect 246022 256776 246028 256828
rect 246080 256816 246086 256828
rect 246206 256816 246212 256828
rect 246080 256788 246212 256816
rect 246080 256776 246086 256788
rect 246206 256776 246212 256788
rect 246264 256776 246270 256828
rect 194226 256708 194232 256760
rect 194284 256748 194290 256760
rect 197354 256748 197360 256760
rect 194284 256720 197360 256748
rect 194284 256708 194290 256720
rect 197354 256708 197360 256720
rect 197412 256708 197418 256760
rect 246022 256640 246028 256692
rect 246080 256680 246086 256692
rect 286318 256680 286324 256692
rect 246080 256652 286324 256680
rect 246080 256640 246086 256652
rect 286318 256640 286324 256652
rect 286376 256640 286382 256692
rect 245746 255280 245752 255332
rect 245804 255320 245810 255332
rect 267090 255320 267096 255332
rect 245804 255292 267096 255320
rect 245804 255280 245810 255292
rect 267090 255280 267096 255292
rect 267148 255280 267154 255332
rect 195698 253988 195704 254040
rect 195756 254028 195762 254040
rect 197446 254028 197452 254040
rect 195756 254000 197452 254028
rect 195756 253988 195762 254000
rect 197446 253988 197452 254000
rect 197504 253988 197510 254040
rect 47578 253920 47584 253972
rect 47636 253960 47642 253972
rect 197354 253960 197360 253972
rect 47636 253932 197360 253960
rect 47636 253920 47642 253932
rect 197354 253920 197360 253932
rect 197412 253920 197418 253972
rect 3418 253172 3424 253224
rect 3476 253212 3482 253224
rect 191098 253212 191104 253224
rect 3476 253184 191104 253212
rect 3476 253172 3482 253184
rect 191098 253172 191104 253184
rect 191156 253172 191162 253224
rect 194134 252560 194140 252612
rect 194192 252600 194198 252612
rect 197354 252600 197360 252612
rect 194192 252572 197360 252600
rect 194192 252560 194198 252572
rect 197354 252560 197360 252572
rect 197412 252560 197418 252612
rect 246022 252560 246028 252612
rect 246080 252600 246086 252612
rect 280982 252600 280988 252612
rect 246080 252572 280988 252600
rect 246080 252560 246086 252572
rect 280982 252560 280988 252572
rect 281040 252560 281046 252612
rect 246482 252084 246488 252136
rect 246540 252124 246546 252136
rect 246666 252124 246672 252136
rect 246540 252096 246672 252124
rect 246540 252084 246546 252096
rect 246666 252084 246672 252096
rect 246724 252084 246730 252136
rect 246022 251200 246028 251252
rect 246080 251240 246086 251252
rect 291838 251240 291844 251252
rect 246080 251212 291844 251240
rect 246080 251200 246086 251212
rect 291838 251200 291844 251212
rect 291896 251200 291902 251252
rect 136634 251132 136640 251184
rect 136692 251172 136698 251184
rect 197354 251172 197360 251184
rect 136692 251144 197360 251172
rect 136692 251132 136698 251144
rect 197354 251132 197360 251144
rect 197412 251132 197418 251184
rect 246022 249772 246028 249824
rect 246080 249812 246086 249824
rect 284478 249812 284484 249824
rect 246080 249784 284484 249812
rect 246080 249772 246086 249784
rect 284478 249772 284484 249784
rect 284536 249772 284542 249824
rect 196342 248480 196348 248532
rect 196400 248520 196406 248532
rect 197538 248520 197544 248532
rect 196400 248492 197544 248520
rect 196400 248480 196406 248492
rect 197538 248480 197544 248492
rect 197596 248480 197602 248532
rect 245654 248344 245660 248396
rect 245712 248384 245718 248396
rect 251910 248384 251916 248396
rect 245712 248356 251916 248384
rect 245712 248344 245718 248356
rect 251910 248344 251916 248356
rect 251968 248344 251974 248396
rect 246022 248140 246028 248192
rect 246080 248180 246086 248192
rect 250622 248180 250628 248192
rect 246080 248152 250628 248180
rect 246080 248140 246086 248152
rect 250622 248140 250628 248152
rect 250680 248140 250686 248192
rect 196526 247052 196532 247104
rect 196584 247092 196590 247104
rect 197998 247092 198004 247104
rect 196584 247064 198004 247092
rect 196584 247052 196590 247064
rect 197998 247052 198004 247064
rect 198056 247052 198062 247104
rect 3602 246984 3608 247036
rect 3660 247024 3666 247036
rect 197354 247024 197360 247036
rect 3660 246996 197360 247024
rect 3660 246984 3666 246996
rect 197354 246984 197360 246996
rect 197412 246984 197418 247036
rect 246022 246984 246028 247036
rect 246080 247024 246086 247036
rect 255958 247024 255964 247036
rect 246080 246996 255964 247024
rect 246080 246984 246086 246996
rect 255958 246984 255964 246996
rect 256016 246984 256022 247036
rect 246022 245624 246028 245676
rect 246080 245664 246086 245676
rect 280154 245664 280160 245676
rect 246080 245636 280160 245664
rect 246080 245624 246086 245636
rect 280154 245624 280160 245636
rect 280212 245624 280218 245676
rect 248966 244264 248972 244316
rect 249024 244304 249030 244316
rect 579798 244304 579804 244316
rect 249024 244276 579804 244304
rect 249024 244264 249030 244276
rect 579798 244264 579804 244276
rect 579856 244264 579862 244316
rect 11698 244196 11704 244248
rect 11756 244236 11762 244248
rect 197354 244236 197360 244248
rect 11756 244208 197360 244236
rect 11756 244196 11762 244208
rect 197354 244196 197360 244208
rect 197412 244196 197418 244248
rect 245654 244196 245660 244248
rect 245712 244236 245718 244248
rect 295978 244236 295984 244248
rect 245712 244208 295984 244236
rect 245712 244196 245718 244208
rect 295978 244196 295984 244208
rect 296036 244196 296042 244248
rect 195790 244128 195796 244180
rect 195848 244168 195854 244180
rect 197446 244168 197452 244180
rect 195848 244140 197452 244168
rect 195848 244128 195854 244140
rect 197446 244128 197452 244140
rect 197504 244128 197510 244180
rect 246022 242904 246028 242956
rect 246080 242944 246086 242956
rect 292758 242944 292764 242956
rect 246080 242916 292764 242944
rect 246080 242904 246086 242916
rect 292758 242904 292764 242916
rect 292816 242904 292822 242956
rect 249426 242156 249432 242208
rect 249484 242196 249490 242208
rect 580350 242196 580356 242208
rect 249484 242168 580356 242196
rect 249484 242156 249490 242168
rect 580350 242156 580356 242168
rect 580408 242156 580414 242208
rect 195790 241476 195796 241528
rect 195848 241516 195854 241528
rect 197998 241516 198004 241528
rect 195848 241488 198004 241516
rect 195848 241476 195854 241488
rect 197998 241476 198004 241488
rect 198056 241476 198062 241528
rect 246022 241408 246028 241460
rect 246080 241448 246086 241460
rect 294598 241448 294604 241460
rect 246080 241420 294604 241448
rect 246080 241408 246086 241420
rect 294598 241408 294604 241420
rect 294656 241408 294662 241460
rect 245286 240864 245292 240916
rect 245344 240904 245350 240916
rect 462314 240904 462320 240916
rect 245344 240876 462320 240904
rect 245344 240864 245350 240876
rect 462314 240864 462320 240876
rect 462372 240864 462378 240916
rect 580258 240836 580264 240848
rect 244200 240808 580264 240836
rect 243906 240292 243912 240304
rect 242912 240264 243912 240292
rect 242912 240168 242940 240264
rect 243906 240252 243912 240264
rect 243964 240252 243970 240304
rect 3050 240116 3056 240168
rect 3108 240156 3114 240168
rect 201402 240156 201408 240168
rect 3108 240128 201408 240156
rect 3108 240116 3114 240128
rect 201402 240116 201408 240128
rect 201460 240116 201466 240168
rect 242894 240116 242900 240168
rect 242952 240116 242958 240168
rect 243814 240116 243820 240168
rect 243872 240156 243878 240168
rect 244200 240156 244228 240808
rect 580258 240796 580264 240808
rect 580316 240796 580322 240848
rect 244274 240728 244280 240780
rect 244332 240768 244338 240780
rect 580442 240768 580448 240780
rect 244332 240740 580448 240768
rect 244332 240728 244338 240740
rect 580442 240728 580448 240740
rect 580500 240728 580506 240780
rect 243872 240128 244228 240156
rect 243872 240116 243878 240128
rect 7558 240048 7564 240100
rect 7616 240088 7622 240100
rect 212718 240088 212724 240100
rect 7616 240060 212724 240088
rect 7616 240048 7622 240060
rect 212718 240048 212724 240060
rect 212776 240048 212782 240100
rect 238854 240048 238860 240100
rect 238912 240088 238918 240100
rect 529198 240088 529204 240100
rect 238912 240060 529204 240088
rect 238912 240048 238918 240060
rect 529198 240048 529204 240060
rect 529256 240048 529262 240100
rect 175918 239980 175924 240032
rect 175976 240020 175982 240032
rect 232958 240020 232964 240032
rect 175976 239992 232964 240020
rect 175976 239980 175982 239992
rect 232958 239980 232964 239992
rect 233016 239980 233022 240032
rect 235910 239980 235916 240032
rect 235968 240020 235974 240032
rect 235968 239992 248414 240020
rect 235968 239980 235974 239992
rect 201402 239912 201408 239964
rect 201460 239952 201466 239964
rect 225230 239952 225236 239964
rect 201460 239924 225236 239952
rect 201460 239912 201466 239924
rect 225230 239912 225236 239924
rect 225288 239912 225294 239964
rect 248386 239952 248414 239992
rect 249058 239952 249064 239964
rect 248386 239924 249064 239952
rect 249058 239912 249064 239924
rect 249116 239912 249122 239964
rect 216582 239844 216588 239896
rect 216640 239884 216646 239896
rect 243538 239884 243544 239896
rect 216640 239856 243544 239884
rect 216640 239844 216646 239856
rect 243538 239844 243544 239856
rect 243596 239844 243602 239896
rect 243814 239844 243820 239896
rect 243872 239884 243878 239896
rect 244274 239884 244280 239896
rect 243872 239856 244280 239884
rect 243872 239844 243878 239856
rect 244274 239844 244280 239856
rect 244332 239844 244338 239896
rect 245286 239844 245292 239896
rect 245344 239884 245350 239896
rect 248966 239884 248972 239896
rect 245344 239856 248972 239884
rect 245344 239844 245350 239856
rect 248966 239844 248972 239856
rect 249024 239844 249030 239896
rect 196710 239776 196716 239828
rect 196768 239816 196774 239828
rect 221918 239816 221924 239828
rect 196768 239788 221924 239816
rect 196768 239776 196774 239788
rect 221918 239776 221924 239788
rect 221976 239776 221982 239828
rect 227622 239776 227628 239828
rect 227680 239816 227686 239828
rect 251818 239816 251824 239828
rect 227680 239788 251824 239816
rect 227680 239776 227686 239788
rect 251818 239776 251824 239788
rect 251876 239776 251882 239828
rect 233510 239708 233516 239760
rect 233568 239748 233574 239760
rect 243446 239748 243452 239760
rect 233568 239720 243452 239748
rect 233568 239708 233574 239720
rect 243446 239708 243452 239720
rect 243504 239708 243510 239760
rect 243538 239708 243544 239760
rect 243596 239748 243602 239760
rect 250714 239748 250720 239760
rect 243596 239720 250720 239748
rect 243596 239708 243602 239720
rect 250714 239708 250720 239720
rect 250772 239708 250778 239760
rect 221366 239640 221372 239692
rect 221424 239680 221430 239692
rect 364334 239680 364340 239692
rect 221424 239652 364340 239680
rect 221424 239640 221430 239652
rect 364334 239640 364340 239652
rect 364392 239640 364398 239692
rect 232590 239572 232596 239624
rect 232648 239612 232654 239624
rect 494054 239612 494060 239624
rect 232648 239584 494060 239612
rect 232648 239572 232654 239584
rect 494054 239572 494060 239584
rect 494112 239572 494118 239624
rect 198182 239504 198188 239556
rect 198240 239544 198246 239556
rect 231946 239544 231952 239556
rect 198240 239516 231952 239544
rect 198240 239504 198246 239516
rect 231946 239504 231952 239516
rect 232004 239504 232010 239556
rect 243446 239504 243452 239556
rect 243504 239544 243510 239556
rect 250438 239544 250444 239556
rect 243504 239516 250444 239544
rect 243504 239504 243510 239516
rect 250438 239504 250444 239516
rect 250496 239504 250502 239556
rect 199286 239436 199292 239488
rect 199344 239476 199350 239488
rect 281718 239476 281724 239488
rect 199344 239448 281724 239476
rect 199344 239436 199350 239448
rect 281718 239436 281724 239448
rect 281776 239436 281782 239488
rect 3510 239368 3516 239420
rect 3568 239408 3574 239420
rect 233142 239408 233148 239420
rect 3568 239380 233148 239408
rect 3568 239368 3574 239380
rect 233142 239368 233148 239380
rect 233200 239368 233206 239420
rect 239214 239368 239220 239420
rect 239272 239408 239278 239420
rect 245286 239408 245292 239420
rect 239272 239380 245292 239408
rect 239272 239368 239278 239380
rect 245286 239368 245292 239380
rect 245344 239368 245350 239420
rect 228174 239300 228180 239352
rect 228232 239340 228238 239352
rect 247678 239340 247684 239352
rect 228232 239312 247684 239340
rect 228232 239300 228238 239312
rect 247678 239300 247684 239312
rect 247736 239300 247742 239352
rect 50338 238688 50344 238740
rect 50396 238728 50402 238740
rect 219526 238728 219532 238740
rect 50396 238700 219532 238728
rect 50396 238688 50402 238700
rect 219526 238688 219532 238700
rect 219584 238688 219590 238740
rect 240686 238688 240692 238740
rect 240744 238728 240750 238740
rect 243906 238728 243912 238740
rect 240744 238700 243912 238728
rect 240744 238688 240750 238700
rect 243906 238688 243912 238700
rect 243964 238688 243970 238740
rect 108298 238620 108304 238672
rect 108356 238660 108362 238672
rect 214558 238660 214564 238672
rect 108356 238632 214564 238660
rect 108356 238620 108362 238632
rect 214558 238620 214564 238632
rect 214616 238620 214622 238672
rect 239766 238620 239772 238672
rect 239824 238660 239830 238672
rect 253198 238660 253204 238672
rect 239824 238632 253204 238660
rect 239824 238620 239830 238632
rect 253198 238620 253204 238632
rect 253256 238620 253262 238672
rect 202046 238552 202052 238604
rect 202104 238592 202110 238604
rect 243814 238592 243820 238604
rect 202104 238564 243820 238592
rect 202104 238552 202110 238564
rect 243814 238552 243820 238564
rect 243872 238552 243878 238604
rect 204438 238484 204444 238536
rect 204496 238524 204502 238536
rect 243722 238524 243728 238536
rect 204496 238496 243728 238524
rect 204496 238484 204502 238496
rect 243722 238484 243728 238496
rect 243780 238484 243786 238536
rect 191098 238416 191104 238468
rect 191156 238456 191162 238468
rect 231486 238456 231492 238468
rect 191156 238428 231492 238456
rect 191156 238416 191162 238428
rect 231486 238416 231492 238428
rect 231544 238416 231550 238468
rect 236454 238416 236460 238468
rect 236512 238456 236518 238468
rect 249426 238456 249432 238468
rect 236512 238428 249432 238456
rect 236512 238416 236518 238428
rect 249426 238416 249432 238428
rect 249484 238416 249490 238468
rect 195330 238348 195336 238400
rect 195388 238388 195394 238400
rect 209222 238388 209228 238400
rect 195388 238360 209228 238388
rect 195388 238348 195394 238360
rect 209222 238348 209228 238360
rect 209280 238348 209286 238400
rect 215662 238348 215668 238400
rect 215720 238388 215726 238400
rect 229738 238388 229744 238400
rect 215720 238360 229744 238388
rect 215720 238348 215726 238360
rect 229738 238348 229744 238360
rect 229796 238348 229802 238400
rect 233142 238348 233148 238400
rect 233200 238388 233206 238400
rect 242710 238388 242716 238400
rect 233200 238360 242716 238388
rect 233200 238348 233206 238360
rect 242710 238348 242716 238360
rect 242768 238348 242774 238400
rect 195882 238280 195888 238332
rect 195940 238320 195946 238332
rect 208854 238320 208860 238332
rect 195940 238292 208860 238320
rect 195940 238280 195946 238292
rect 208854 238280 208860 238292
rect 208912 238280 208918 238332
rect 215110 238280 215116 238332
rect 215168 238320 215174 238332
rect 234614 238320 234620 238332
rect 215168 238292 234620 238320
rect 215168 238280 215174 238292
rect 234614 238280 234620 238292
rect 234672 238280 234678 238332
rect 218974 238212 218980 238264
rect 219032 238252 219038 238264
rect 290090 238252 290096 238264
rect 219032 238224 290096 238252
rect 219032 238212 219038 238224
rect 290090 238212 290096 238224
rect 290148 238212 290154 238264
rect 213086 238144 213092 238196
rect 213144 238184 213150 238196
rect 289998 238184 290004 238196
rect 213144 238156 290004 238184
rect 213144 238144 213150 238156
rect 289998 238144 290004 238156
rect 290056 238144 290062 238196
rect 207382 238076 207388 238128
rect 207440 238116 207446 238128
rect 290182 238116 290188 238128
rect 207440 238088 290188 238116
rect 207440 238076 207446 238088
rect 290182 238076 290188 238088
rect 290240 238076 290246 238128
rect 200574 238008 200580 238060
rect 200632 238048 200638 238060
rect 287514 238048 287520 238060
rect 200632 238020 287520 238048
rect 200632 238008 200638 238020
rect 287514 238008 287520 238020
rect 287572 238008 287578 238060
rect 234982 237940 234988 237992
rect 235040 237980 235046 237992
rect 260098 237980 260104 237992
rect 235040 237952 260104 237980
rect 235040 237940 235046 237952
rect 260098 237940 260104 237952
rect 260156 237940 260162 237992
rect 240870 237396 240876 237448
rect 240928 237436 240934 237448
rect 244458 237436 244464 237448
rect 240928 237408 244464 237436
rect 240928 237396 240934 237408
rect 244458 237396 244464 237408
rect 244516 237396 244522 237448
rect 216030 237328 216036 237380
rect 216088 237368 216094 237380
rect 258718 237368 258724 237380
rect 216088 237340 258724 237368
rect 216088 237328 216094 237340
rect 258718 237328 258724 237340
rect 258776 237328 258782 237380
rect 197630 237124 197636 237176
rect 197688 237164 197694 237176
rect 229554 237164 229560 237176
rect 197688 237136 229560 237164
rect 197688 237124 197694 237136
rect 229554 237124 229560 237136
rect 229612 237124 229618 237176
rect 230566 237124 230572 237176
rect 230624 237164 230630 237176
rect 231854 237164 231860 237176
rect 230624 237136 231860 237164
rect 230624 237124 230630 237136
rect 231854 237124 231860 237136
rect 231912 237124 231918 237176
rect 209038 236988 209044 237040
rect 209096 237028 209102 237040
rect 229646 237028 229652 237040
rect 209096 237000 229652 237028
rect 209096 236988 209102 237000
rect 229646 236988 229652 237000
rect 229704 236988 229710 237040
rect 199654 236852 199660 236904
rect 199712 236892 199718 236904
rect 230750 236892 230756 236904
rect 199712 236864 230756 236892
rect 199712 236852 199718 236864
rect 230750 236852 230756 236864
rect 230808 236852 230814 236904
rect 199562 236784 199568 236836
rect 199620 236824 199626 236836
rect 231210 236824 231216 236836
rect 199620 236796 231216 236824
rect 199620 236784 199626 236796
rect 231210 236784 231216 236796
rect 231268 236784 231274 236836
rect 212166 236716 212172 236768
rect 212224 236756 212230 236768
rect 266998 236756 267004 236768
rect 212224 236728 267004 236756
rect 212224 236716 212230 236728
rect 266998 236716 267004 236728
rect 267056 236716 267062 236768
rect 25498 236648 25504 236700
rect 25556 236688 25562 236700
rect 230198 236688 230204 236700
rect 25556 236660 230204 236688
rect 25556 236648 25562 236660
rect 230198 236648 230204 236660
rect 230256 236648 230262 236700
rect 238018 236648 238024 236700
rect 238076 236688 238082 236700
rect 245746 236688 245752 236700
rect 238076 236660 245752 236688
rect 238076 236648 238082 236660
rect 245746 236648 245752 236660
rect 245804 236648 245810 236700
rect 240778 236036 240784 236088
rect 240836 236076 240842 236088
rect 245838 236076 245844 236088
rect 240836 236048 245844 236076
rect 240836 236036 240842 236048
rect 245838 236036 245844 236048
rect 245896 236036 245902 236088
rect 204990 235968 204996 236020
rect 205048 236008 205054 236020
rect 206278 236008 206284 236020
rect 205048 235980 206284 236008
rect 205048 235968 205054 235980
rect 206278 235968 206284 235980
rect 206336 235968 206342 236020
rect 239398 235968 239404 236020
rect 239456 236008 239462 236020
rect 243262 236008 243268 236020
rect 239456 235980 243268 236008
rect 239456 235968 239462 235980
rect 243262 235968 243268 235980
rect 243320 235968 243326 236020
rect 238110 235424 238116 235476
rect 238168 235464 238174 235476
rect 245654 235464 245660 235476
rect 238168 235436 245660 235464
rect 238168 235424 238174 235436
rect 245654 235424 245660 235436
rect 245712 235424 245718 235476
rect 236638 235356 236644 235408
rect 236696 235396 236702 235408
rect 246114 235396 246120 235408
rect 236696 235368 246120 235396
rect 236696 235356 236702 235368
rect 246114 235356 246120 235368
rect 246172 235356 246178 235408
rect 199470 235288 199476 235340
rect 199528 235328 199534 235340
rect 230658 235328 230664 235340
rect 199528 235300 230664 235328
rect 199528 235288 199534 235300
rect 230658 235288 230664 235300
rect 230716 235288 230722 235340
rect 197722 235220 197728 235272
rect 197780 235260 197786 235272
rect 281810 235260 281816 235272
rect 197780 235232 281816 235260
rect 197780 235220 197786 235232
rect 281810 235220 281816 235232
rect 281868 235220 281874 235272
rect 237282 234608 237288 234660
rect 237340 234648 237346 234660
rect 238294 234648 238300 234660
rect 237340 234620 238300 234648
rect 237340 234608 237346 234620
rect 238294 234608 238300 234620
rect 238352 234608 238358 234660
rect 199378 233928 199384 233980
rect 199436 233968 199442 233980
rect 230566 233968 230572 233980
rect 199436 233940 230572 233968
rect 199436 233928 199442 233940
rect 230566 233928 230572 233940
rect 230624 233928 230630 233980
rect 7558 233860 7564 233912
rect 7616 233900 7622 233912
rect 210326 233900 210332 233912
rect 7616 233872 210332 233900
rect 7616 233860 7622 233872
rect 210326 233860 210332 233872
rect 210384 233860 210390 233912
rect 235258 233656 235264 233708
rect 235316 233696 235322 233708
rect 237926 233696 237932 233708
rect 235316 233668 237932 233696
rect 235316 233656 235322 233668
rect 237926 233656 237932 233668
rect 237984 233656 237990 233708
rect 291930 233180 291936 233232
rect 291988 233220 291994 233232
rect 579982 233220 579988 233232
rect 291988 233192 579988 233220
rect 291988 233180 291994 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 180058 229712 180064 229764
rect 180116 229752 180122 229764
rect 245930 229752 245936 229764
rect 180116 229724 245936 229752
rect 180116 229712 180122 229724
rect 245930 229712 245936 229724
rect 245988 229712 245994 229764
rect 256050 219376 256056 219428
rect 256108 219416 256114 219428
rect 580166 219416 580172 219428
rect 256108 219388 580172 219416
rect 256108 219376 256114 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 17218 215268 17224 215280
rect 3384 215240 17224 215268
rect 3384 215228 3390 215240
rect 17218 215228 17224 215240
rect 17276 215228 17282 215280
rect 249242 206932 249248 206984
rect 249300 206972 249306 206984
rect 579798 206972 579804 206984
rect 249300 206944 579804 206972
rect 249300 206932 249306 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 238110 202824 238116 202836
rect 3108 202796 238116 202824
rect 3108 202784 3114 202796
rect 238110 202784 238116 202796
rect 238168 202784 238174 202836
rect 235350 199384 235356 199436
rect 235408 199424 235414 199436
rect 580258 199424 580264 199436
rect 235408 199396 580264 199424
rect 235408 199384 235414 199396
rect 580258 199384 580264 199396
rect 580316 199384 580322 199436
rect 208302 197956 208308 198008
rect 208360 197996 208366 198008
rect 286318 197996 286324 198008
rect 208360 197968 286324 197996
rect 208360 197956 208366 197968
rect 286318 197956 286324 197968
rect 286376 197956 286382 198008
rect 249150 193128 249156 193180
rect 249208 193168 249214 193180
rect 580166 193168 580172 193180
rect 249208 193140 580172 193168
rect 249208 193128 249214 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 214190 191088 214196 191140
rect 214248 191128 214254 191140
rect 286410 191128 286416 191140
rect 214248 191100 286416 191128
rect 214248 191088 214254 191100
rect 286410 191088 286416 191100
rect 286468 191088 286474 191140
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 192478 189020 192484 189032
rect 3476 188992 192484 189020
rect 3476 188980 3482 188992
rect 192478 188980 192484 188992
rect 192536 188980 192542 189032
rect 206462 188368 206468 188420
rect 206520 188408 206526 188420
rect 229462 188408 229468 188420
rect 206520 188380 229468 188408
rect 206520 188368 206526 188380
rect 229462 188368 229468 188380
rect 229520 188368 229526 188420
rect 229094 188300 229100 188352
rect 229152 188340 229158 188352
rect 284570 188340 284576 188352
rect 229152 188312 284576 188340
rect 229152 188300 229158 188312
rect 284570 188300 284576 188312
rect 284628 188300 284634 188352
rect 204070 187076 204076 187128
rect 204128 187116 204134 187128
rect 233418 187116 233424 187128
rect 204128 187088 233424 187116
rect 204128 187076 204134 187088
rect 233418 187076 233424 187088
rect 233476 187076 233482 187128
rect 222286 187008 222292 187060
rect 222344 187048 222350 187060
rect 285674 187048 285680 187060
rect 222344 187020 285680 187048
rect 222344 187008 222350 187020
rect 285674 187008 285680 187020
rect 285732 187008 285738 187060
rect 205910 186940 205916 186992
rect 205968 186980 205974 186992
rect 284662 186980 284668 186992
rect 205968 186952 284668 186980
rect 205968 186940 205974 186952
rect 284662 186940 284668 186952
rect 284720 186940 284726 186992
rect 218054 184356 218060 184408
rect 218112 184396 218118 184408
rect 233510 184396 233516 184408
rect 218112 184368 233516 184396
rect 218112 184356 218118 184368
rect 233510 184356 233516 184368
rect 233568 184356 233574 184408
rect 237374 184356 237380 184408
rect 237432 184396 237438 184408
rect 286226 184396 286232 184408
rect 237432 184368 286232 184396
rect 237432 184356 237438 184368
rect 286226 184356 286232 184368
rect 286284 184356 286290 184408
rect 224310 184288 224316 184340
rect 224368 184328 224374 184340
rect 281994 184328 282000 184340
rect 224368 184300 282000 184328
rect 224368 184288 224374 184300
rect 281994 184288 282000 184300
rect 282052 184288 282058 184340
rect 226702 184220 226708 184272
rect 226760 184260 226766 184272
rect 285950 184260 285956 184272
rect 226760 184232 285956 184260
rect 226760 184220 226766 184232
rect 285950 184220 285956 184232
rect 286008 184220 286014 184272
rect 211246 184152 211252 184204
rect 211304 184192 211310 184204
rect 284938 184192 284944 184204
rect 211304 184164 284944 184192
rect 211304 184152 211310 184164
rect 284938 184152 284944 184164
rect 284996 184152 285002 184204
rect 213638 182996 213644 183048
rect 213696 183036 213702 183048
rect 229278 183036 229284 183048
rect 213696 183008 229284 183036
rect 213696 182996 213702 183008
rect 229278 182996 229284 183008
rect 229336 182996 229342 183048
rect 203518 182928 203524 182980
rect 203576 182968 203582 182980
rect 281074 182968 281080 182980
rect 203576 182940 281080 182968
rect 203576 182928 203582 182940
rect 281074 182928 281080 182940
rect 281132 182928 281138 182980
rect 201494 182860 201500 182912
rect 201552 182900 201558 182912
rect 290274 182900 290280 182912
rect 201552 182872 290280 182900
rect 201552 182860 201558 182872
rect 290274 182860 290280 182872
rect 290332 182860 290338 182912
rect 194134 182792 194140 182844
rect 194192 182832 194198 182844
rect 289170 182832 289176 182844
rect 194192 182804 289176 182832
rect 194192 182792 194198 182804
rect 289170 182792 289176 182804
rect 289228 182792 289234 182844
rect 211798 181636 211804 181688
rect 211856 181676 211862 181688
rect 232130 181676 232136 181688
rect 211856 181648 232136 181676
rect 211856 181636 211862 181648
rect 232130 181636 232136 181648
rect 232188 181636 232194 181688
rect 236822 181636 236828 181688
rect 236880 181676 236886 181688
rect 284846 181676 284852 181688
rect 236880 181648 284852 181676
rect 236880 181636 236886 181648
rect 284846 181636 284852 181648
rect 284904 181636 284910 181688
rect 226150 181568 226156 181620
rect 226208 181608 226214 181620
rect 283282 181608 283288 181620
rect 226208 181580 283288 181608
rect 226208 181568 226214 181580
rect 283282 181568 283288 181580
rect 283340 181568 283346 181620
rect 218422 181500 218428 181552
rect 218480 181540 218486 181552
rect 280338 181540 280344 181552
rect 218480 181512 280344 181540
rect 218480 181500 218486 181512
rect 280338 181500 280344 181512
rect 280396 181500 280402 181552
rect 217502 181432 217508 181484
rect 217560 181472 217566 181484
rect 285122 181472 285128 181484
rect 217560 181444 285128 181472
rect 217560 181432 217566 181444
rect 285122 181432 285128 181444
rect 285180 181432 285186 181484
rect 199194 180752 199200 180804
rect 199252 180792 199258 180804
rect 230934 180792 230940 180804
rect 199252 180764 230940 180792
rect 199252 180752 199258 180764
rect 230934 180752 230940 180764
rect 230992 180752 230998 180804
rect 196894 180684 196900 180736
rect 196952 180724 196958 180736
rect 233970 180724 233976 180736
rect 196952 180696 233976 180724
rect 196952 180684 196958 180696
rect 233970 180684 233976 180696
rect 234028 180684 234034 180736
rect 196802 180616 196808 180668
rect 196860 180656 196866 180668
rect 233694 180656 233700 180668
rect 196860 180628 233700 180656
rect 196860 180616 196866 180628
rect 233694 180616 233700 180628
rect 233752 180616 233758 180668
rect 194410 180548 194416 180600
rect 194468 180588 194474 180600
rect 232314 180588 232320 180600
rect 194468 180560 232320 180588
rect 194468 180548 194474 180560
rect 232314 180548 232320 180560
rect 232372 180548 232378 180600
rect 195422 180480 195428 180532
rect 195480 180520 195486 180532
rect 229370 180520 229376 180532
rect 195480 180492 229376 180520
rect 195480 180480 195486 180492
rect 229370 180480 229376 180492
rect 229428 180480 229434 180532
rect 195514 180412 195520 180464
rect 195572 180452 195578 180464
rect 234890 180452 234896 180464
rect 195572 180424 234896 180452
rect 195572 180412 195578 180424
rect 234890 180412 234896 180424
rect 234948 180412 234954 180464
rect 193030 180344 193036 180396
rect 193088 180384 193094 180396
rect 233786 180384 233792 180396
rect 193088 180356 233792 180384
rect 193088 180344 193094 180356
rect 233786 180344 233792 180356
rect 233844 180344 233850 180396
rect 246666 180344 246672 180396
rect 246724 180384 246730 180396
rect 279142 180384 279148 180396
rect 246724 180356 279148 180384
rect 246724 180344 246730 180356
rect 279142 180344 279148 180356
rect 279200 180344 279206 180396
rect 228726 180276 228732 180328
rect 228784 180316 228790 180328
rect 285030 180316 285036 180328
rect 228784 180288 285036 180316
rect 228784 180276 228790 180288
rect 285030 180276 285036 180288
rect 285088 180276 285094 180328
rect 220998 180208 221004 180260
rect 221056 180248 221062 180260
rect 286042 180248 286048 180260
rect 221056 180220 286048 180248
rect 221056 180208 221062 180220
rect 286042 180208 286048 180220
rect 286100 180208 286106 180260
rect 205358 180140 205364 180192
rect 205416 180180 205422 180192
rect 284754 180180 284760 180192
rect 205416 180152 284760 180180
rect 205416 180140 205422 180152
rect 284754 180140 284760 180152
rect 284812 180140 284818 180192
rect 200206 180072 200212 180124
rect 200264 180112 200270 180124
rect 282914 180112 282920 180124
rect 200264 180084 282920 180112
rect 200264 180072 200270 180084
rect 282914 180072 282920 180084
rect 282972 180072 282978 180124
rect 201126 180004 201132 180056
rect 201184 180044 201190 180056
rect 229830 180044 229836 180056
rect 201184 180016 229836 180044
rect 201184 180004 201190 180016
rect 229830 180004 229836 180016
rect 229888 180004 229894 180056
rect 223390 179936 223396 179988
rect 223448 179976 223454 179988
rect 232222 179976 232228 179988
rect 223448 179948 232228 179976
rect 223448 179936 223454 179948
rect 232222 179936 232228 179948
rect 232280 179936 232286 179988
rect 222838 179460 222844 179512
rect 222896 179500 222902 179512
rect 229094 179500 229100 179512
rect 222896 179472 229100 179500
rect 222896 179460 222902 179472
rect 229094 179460 229100 179472
rect 229152 179460 229158 179512
rect 252002 179324 252008 179376
rect 252060 179364 252066 179376
rect 579982 179364 579988 179376
rect 252060 179336 579988 179364
rect 252060 179324 252066 179336
rect 579982 179324 579988 179336
rect 580040 179324 580046 179376
rect 223758 178916 223764 178968
rect 223816 178956 223822 178968
rect 232406 178956 232412 178968
rect 223816 178928 232412 178956
rect 223816 178916 223822 178928
rect 232406 178916 232412 178928
rect 232464 178916 232470 178968
rect 220446 178848 220452 178900
rect 220504 178888 220510 178900
rect 229554 178888 229560 178900
rect 220504 178860 229560 178888
rect 220504 178848 220510 178860
rect 229554 178848 229560 178860
rect 229612 178848 229618 178900
rect 199930 178780 199936 178832
rect 199988 178820 199994 178832
rect 230842 178820 230848 178832
rect 199988 178792 230848 178820
rect 199988 178780 199994 178792
rect 230842 178780 230848 178792
rect 230900 178780 230906 178832
rect 241238 178780 241244 178832
rect 241296 178820 241302 178832
rect 280522 178820 280528 178832
rect 241296 178792 280528 178820
rect 241296 178780 241302 178792
rect 280522 178780 280528 178792
rect 280580 178780 280586 178832
rect 200022 178712 200028 178764
rect 200080 178752 200086 178764
rect 231026 178752 231032 178764
rect 200080 178724 231032 178752
rect 200080 178712 200086 178724
rect 231026 178712 231032 178724
rect 231084 178712 231090 178764
rect 243630 178712 243636 178764
rect 243688 178752 243694 178764
rect 283374 178752 283380 178764
rect 243688 178724 283380 178752
rect 243688 178712 243694 178724
rect 283374 178712 283380 178724
rect 283432 178712 283438 178764
rect 202966 178644 202972 178696
rect 203024 178684 203030 178696
rect 283558 178684 283564 178696
rect 203024 178656 283564 178684
rect 203024 178644 203030 178656
rect 283558 178644 283564 178656
rect 283616 178644 283622 178696
rect 114002 178440 114008 178492
rect 114060 178480 114066 178492
rect 169294 178480 169300 178492
rect 114060 178452 169300 178480
rect 114060 178440 114066 178452
rect 169294 178440 169300 178452
rect 169352 178440 169358 178492
rect 114370 178372 114376 178424
rect 114428 178412 114434 178424
rect 170582 178412 170588 178424
rect 114428 178384 170588 178412
rect 114428 178372 114434 178384
rect 170582 178372 170588 178384
rect 170640 178372 170646 178424
rect 110690 178304 110696 178356
rect 110748 178344 110754 178356
rect 169202 178344 169208 178356
rect 110748 178316 169208 178344
rect 110748 178304 110754 178316
rect 169202 178304 169208 178316
rect 169260 178304 169266 178356
rect 112622 178236 112628 178288
rect 112680 178276 112686 178288
rect 173250 178276 173256 178288
rect 112680 178248 173256 178276
rect 112680 178236 112686 178248
rect 173250 178236 173256 178248
rect 173308 178236 173314 178288
rect 148226 178168 148232 178220
rect 148284 178208 148290 178220
rect 213178 178208 213184 178220
rect 148284 178180 213184 178208
rect 148284 178168 148290 178180
rect 213178 178168 213184 178180
rect 213236 178168 213242 178220
rect 97810 178100 97816 178152
rect 97868 178140 97874 178152
rect 170398 178140 170404 178152
rect 97868 178112 170404 178140
rect 97868 178100 97874 178112
rect 170398 178100 170404 178112
rect 170456 178100 170462 178152
rect 110046 178032 110052 178084
rect 110104 178072 110110 178084
rect 192478 178072 192484 178084
rect 110104 178044 192484 178072
rect 110104 178032 110110 178044
rect 192478 178032 192484 178044
rect 192536 178032 192542 178084
rect 196434 177964 196440 178016
rect 196492 178004 196498 178016
rect 234706 178004 234712 178016
rect 196492 177976 234712 178004
rect 196492 177964 196498 177976
rect 234706 177964 234712 177976
rect 234764 177964 234770 178016
rect 196342 177896 196348 177948
rect 196400 177936 196406 177948
rect 234154 177936 234160 177948
rect 196400 177908 234160 177936
rect 196400 177896 196406 177908
rect 234154 177896 234160 177908
rect 234212 177896 234218 177948
rect 196986 177828 196992 177880
rect 197044 177868 197050 177880
rect 235166 177868 235172 177880
rect 197044 177840 235172 177868
rect 197044 177828 197050 177840
rect 235166 177828 235172 177840
rect 235224 177828 235230 177880
rect 246574 177828 246580 177880
rect 246632 177868 246638 177880
rect 283466 177868 283472 177880
rect 246632 177840 283472 177868
rect 246632 177828 246638 177840
rect 283466 177828 283472 177840
rect 283524 177828 283530 177880
rect 195790 177760 195796 177812
rect 195848 177800 195854 177812
rect 234798 177800 234804 177812
rect 195848 177772 234804 177800
rect 195848 177760 195854 177772
rect 234798 177760 234804 177772
rect 234856 177760 234862 177812
rect 240318 177760 240324 177812
rect 240376 177800 240382 177812
rect 283006 177800 283012 177812
rect 240376 177772 283012 177800
rect 240376 177760 240382 177772
rect 283006 177760 283012 177772
rect 283064 177760 283070 177812
rect 195606 177692 195612 177744
rect 195664 177732 195670 177744
rect 235074 177732 235080 177744
rect 195664 177704 235080 177732
rect 195664 177692 195670 177704
rect 235074 177692 235080 177704
rect 235132 177692 235138 177744
rect 244182 177692 244188 177744
rect 244240 177732 244246 177744
rect 287882 177732 287888 177744
rect 244240 177704 287888 177732
rect 244240 177692 244246 177704
rect 287882 177692 287888 177704
rect 287940 177692 287946 177744
rect 196526 177624 196532 177676
rect 196584 177664 196590 177676
rect 233234 177664 233240 177676
rect 196584 177636 233240 177664
rect 196584 177624 196590 177636
rect 233234 177624 233240 177636
rect 233292 177624 233298 177676
rect 234062 177624 234068 177676
rect 234120 177664 234126 177676
rect 288986 177664 288992 177676
rect 234120 177636 288992 177664
rect 234120 177624 234126 177636
rect 288986 177624 288992 177636
rect 289044 177624 289050 177676
rect 199838 177556 199844 177608
rect 199896 177596 199902 177608
rect 199896 177568 219434 177596
rect 199896 177556 199902 177568
rect 134518 177488 134524 177540
rect 134576 177528 134582 177540
rect 165154 177528 165160 177540
rect 134576 177500 165160 177528
rect 134576 177488 134582 177500
rect 165154 177488 165160 177500
rect 165212 177488 165218 177540
rect 219406 177528 219434 177568
rect 224862 177556 224868 177608
rect 224920 177596 224926 177608
rect 229186 177596 229192 177608
rect 224920 177568 229192 177596
rect 224920 177556 224926 177568
rect 229186 177556 229192 177568
rect 229244 177556 229250 177608
rect 232038 177556 232044 177608
rect 232096 177596 232102 177608
rect 287790 177596 287796 177608
rect 232096 177568 287796 177596
rect 232096 177556 232102 177568
rect 287790 177556 287796 177568
rect 287848 177556 287854 177608
rect 230474 177528 230480 177540
rect 219406 177500 230480 177528
rect 230474 177488 230480 177500
rect 230532 177488 230538 177540
rect 233878 177488 233884 177540
rect 233936 177528 233942 177540
rect 286134 177528 286140 177540
rect 233936 177500 286140 177528
rect 233936 177488 233942 177500
rect 286134 177488 286140 177500
rect 286192 177488 286198 177540
rect 133138 177420 133144 177472
rect 133196 177460 133202 177472
rect 165246 177460 165252 177472
rect 133196 177432 165252 177460
rect 133196 177420 133202 177432
rect 165246 177420 165252 177432
rect 165304 177420 165310 177472
rect 219894 177420 219900 177472
rect 219952 177460 219958 177472
rect 281534 177460 281540 177472
rect 219952 177432 281540 177460
rect 219952 177420 219958 177432
rect 281534 177420 281540 177432
rect 281592 177420 281598 177472
rect 103330 177352 103336 177404
rect 103388 177392 103394 177404
rect 129734 177392 129740 177404
rect 103388 177364 129740 177392
rect 103388 177352 103394 177364
rect 129734 177352 129740 177364
rect 129792 177352 129798 177404
rect 130930 177352 130936 177404
rect 130988 177392 130994 177404
rect 165706 177392 165712 177404
rect 130988 177364 165712 177392
rect 130988 177352 130994 177364
rect 165706 177352 165712 177364
rect 165764 177352 165770 177404
rect 202598 177352 202604 177404
rect 202656 177392 202662 177404
rect 281626 177392 281632 177404
rect 202656 177364 281632 177392
rect 202656 177352 202662 177364
rect 281626 177352 281632 177364
rect 281684 177352 281690 177404
rect 127986 177284 127992 177336
rect 128044 177324 128050 177336
rect 165338 177324 165344 177336
rect 128044 177296 165344 177324
rect 128044 177284 128050 177296
rect 165338 177284 165344 177296
rect 165396 177284 165402 177336
rect 192938 177284 192944 177336
rect 192996 177324 193002 177336
rect 287698 177324 287704 177336
rect 192996 177296 287704 177324
rect 192996 177284 193002 177296
rect 287698 177284 287704 177296
rect 287756 177284 287762 177336
rect 129458 177216 129464 177268
rect 129516 177256 129522 177268
rect 165798 177256 165804 177268
rect 129516 177228 165804 177256
rect 129516 177216 129522 177228
rect 165798 177216 165804 177228
rect 165856 177216 165862 177268
rect 206830 177216 206836 177268
rect 206888 177256 206894 177268
rect 233602 177256 233608 177268
rect 206888 177228 233608 177256
rect 206888 177216 206894 177228
rect 233602 177216 233608 177228
rect 233660 177216 233666 177268
rect 124490 177148 124496 177200
rect 124548 177188 124554 177200
rect 166350 177188 166356 177200
rect 124548 177160 166356 177188
rect 124548 177148 124554 177160
rect 166350 177148 166356 177160
rect 166408 177148 166414 177200
rect 217134 177148 217140 177200
rect 217192 177188 217198 177200
rect 234982 177188 234988 177200
rect 217192 177160 234988 177188
rect 217192 177148 217198 177160
rect 234982 177148 234988 177160
rect 235040 177148 235046 177200
rect 122282 177080 122288 177132
rect 122340 177120 122346 177132
rect 169386 177120 169392 177132
rect 122340 177092 169392 177120
rect 122340 177080 122346 177092
rect 169386 177080 169392 177092
rect 169444 177080 169450 177132
rect 227254 177080 227260 177132
rect 227312 177120 227318 177132
rect 233878 177120 233884 177132
rect 227312 177092 233884 177120
rect 227312 177080 227318 177092
rect 233878 177080 233884 177092
rect 233936 177080 233942 177132
rect 120810 177012 120816 177064
rect 120868 177052 120874 177064
rect 170674 177052 170680 177064
rect 120868 177024 170680 177052
rect 120868 177012 120874 177024
rect 170674 177012 170680 177024
rect 170732 177012 170738 177064
rect 118418 176944 118424 176996
rect 118476 176984 118482 176996
rect 174630 176984 174636 176996
rect 118476 176956 174636 176984
rect 118476 176944 118482 176956
rect 174630 176944 174636 176956
rect 174688 176944 174694 176996
rect 107010 176876 107016 176928
rect 107068 176916 107074 176928
rect 167822 176916 167828 176928
rect 107068 176888 167828 176916
rect 107068 176876 107074 176888
rect 167822 176876 167828 176888
rect 167880 176876 167886 176928
rect 108114 176808 108120 176860
rect 108172 176848 108178 176860
rect 174538 176848 174544 176860
rect 108172 176820 174544 176848
rect 108172 176808 108178 176820
rect 174538 176808 174544 176820
rect 174596 176808 174602 176860
rect 116946 176740 116952 176792
rect 117004 176780 117010 176792
rect 191098 176780 191104 176792
rect 117004 176752 191104 176780
rect 117004 176740 117010 176752
rect 191098 176740 191104 176752
rect 191156 176740 191162 176792
rect 115842 176672 115848 176724
rect 115900 176712 115906 176724
rect 202138 176712 202144 176724
rect 115900 176684 202144 176712
rect 115900 176672 115906 176684
rect 202138 176672 202144 176684
rect 202196 176672 202202 176724
rect 125686 176604 125692 176656
rect 125744 176644 125750 176656
rect 166534 176644 166540 176656
rect 125744 176616 166540 176644
rect 125744 176604 125750 176616
rect 166534 176604 166540 176616
rect 166592 176604 166598 176656
rect 193122 176604 193128 176656
rect 193180 176644 193186 176656
rect 278774 176644 278780 176656
rect 193180 176616 278780 176644
rect 193180 176604 193186 176616
rect 278774 176604 278780 176616
rect 278832 176604 278838 176656
rect 135714 176536 135720 176588
rect 135772 176576 135778 176588
rect 213914 176576 213920 176588
rect 135772 176548 213920 176576
rect 135772 176536 135778 176548
rect 213914 176536 213920 176548
rect 213972 176536 213978 176588
rect 123110 176468 123116 176520
rect 123168 176508 123174 176520
rect 166442 176508 166448 176520
rect 123168 176480 166448 176508
rect 123168 176468 123174 176480
rect 166442 176468 166448 176480
rect 166500 176468 166506 176520
rect 197078 176468 197084 176520
rect 197136 176508 197142 176520
rect 227714 176508 227720 176520
rect 197136 176480 227720 176508
rect 197136 176468 197142 176480
rect 227714 176468 227720 176480
rect 227772 176468 227778 176520
rect 119430 176400 119436 176452
rect 119488 176440 119494 176452
rect 167730 176440 167736 176452
rect 119488 176412 167736 176440
rect 119488 176400 119494 176412
rect 167730 176400 167736 176412
rect 167788 176400 167794 176452
rect 104618 176332 104624 176384
rect 104676 176372 104682 176384
rect 167638 176372 167644 176384
rect 104676 176344 167644 176372
rect 104676 176332 104682 176344
rect 167638 176332 167644 176344
rect 167696 176332 167702 176384
rect 98362 176264 98368 176316
rect 98420 176304 98426 176316
rect 166258 176304 166264 176316
rect 98420 176276 166264 176304
rect 98420 176264 98426 176276
rect 166258 176264 166264 176276
rect 166316 176264 166322 176316
rect 100754 176196 100760 176248
rect 100812 176236 100818 176248
rect 170490 176236 170496 176248
rect 100812 176208 170496 176236
rect 100812 176196 100818 176208
rect 170490 176196 170496 176208
rect 170548 176196 170554 176248
rect 99466 176128 99472 176180
rect 99524 176168 99530 176180
rect 169110 176168 169116 176180
rect 99524 176140 169116 176168
rect 99524 176128 99530 176140
rect 169110 176128 169116 176140
rect 169168 176128 169174 176180
rect 105722 176060 105728 176112
rect 105780 176100 105786 176112
rect 175918 176100 175924 176112
rect 105780 176072 175924 176100
rect 105780 176060 105786 176072
rect 175918 176060 175924 176072
rect 175976 176060 175982 176112
rect 246298 176060 246304 176112
rect 246356 176100 246362 176112
rect 280706 176100 280712 176112
rect 246356 176072 280712 176100
rect 246356 176060 246362 176072
rect 280706 176060 280712 176072
rect 280764 176060 280770 176112
rect 129734 175992 129740 176044
rect 129792 176032 129798 176044
rect 214558 176032 214564 176044
rect 129792 176004 214564 176032
rect 129792 175992 129798 176004
rect 214558 175992 214564 176004
rect 214616 175992 214622 176044
rect 230750 175992 230756 176044
rect 230808 176032 230814 176044
rect 231302 176032 231308 176044
rect 230808 176004 231308 176032
rect 230808 175992 230814 176004
rect 231302 175992 231308 176004
rect 231360 175992 231366 176044
rect 246482 175992 246488 176044
rect 246540 176032 246546 176044
rect 280614 176032 280620 176044
rect 246540 176004 280620 176032
rect 246540 175992 246546 176004
rect 280614 175992 280620 176004
rect 280672 175992 280678 176044
rect 102042 175924 102048 175976
rect 102100 175964 102106 175976
rect 173158 175964 173164 175976
rect 102100 175936 173164 175964
rect 102100 175924 102106 175936
rect 173158 175924 173164 175936
rect 173216 175924 173222 175976
rect 194318 175924 194324 175976
rect 194376 175964 194382 175976
rect 288434 175964 288440 175976
rect 194376 175936 288440 175964
rect 194376 175924 194382 175936
rect 288434 175924 288440 175936
rect 288492 175924 288498 175976
rect 128170 175856 128176 175908
rect 128228 175896 128234 175908
rect 165430 175896 165436 175908
rect 128228 175868 165436 175896
rect 128228 175856 128234 175868
rect 165430 175856 165436 175868
rect 165488 175856 165494 175908
rect 280430 175856 280436 175908
rect 280488 175896 280494 175908
rect 281074 175896 281080 175908
rect 280488 175868 281080 175896
rect 280488 175856 280494 175868
rect 281074 175856 281080 175868
rect 281132 175856 281138 175908
rect 132034 175788 132040 175840
rect 132092 175828 132098 175840
rect 165522 175828 165528 175840
rect 132092 175800 165528 175828
rect 132092 175788 132098 175800
rect 165522 175788 165528 175800
rect 165580 175788 165586 175840
rect 278038 175788 278044 175840
rect 278096 175828 278102 175840
rect 282086 175828 282092 175840
rect 278096 175800 282092 175828
rect 278096 175788 278102 175800
rect 282086 175788 282092 175800
rect 282144 175788 282150 175840
rect 158898 175720 158904 175772
rect 158956 175760 158962 175772
rect 166626 175760 166632 175772
rect 158956 175732 166632 175760
rect 158956 175720 158962 175732
rect 166626 175720 166632 175732
rect 166684 175720 166690 175772
rect 165154 175176 165160 175228
rect 165212 175216 165218 175228
rect 213914 175216 213920 175228
rect 165212 175188 213920 175216
rect 165212 175176 165218 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 165246 175108 165252 175160
rect 165304 175148 165310 175160
rect 214006 175148 214012 175160
rect 165304 175120 214012 175148
rect 165304 175108 165310 175120
rect 214006 175108 214012 175120
rect 214064 175108 214070 175160
rect 231762 175108 231768 175160
rect 231820 175148 231826 175160
rect 242894 175148 242900 175160
rect 231820 175120 242900 175148
rect 231820 175108 231826 175120
rect 242894 175108 242900 175120
rect 242952 175108 242958 175160
rect 230750 175040 230756 175092
rect 230808 175080 230814 175092
rect 244642 175080 244648 175092
rect 230808 175052 244648 175080
rect 230808 175040 230814 175052
rect 244642 175040 244648 175052
rect 244700 175040 244706 175092
rect 165338 174496 165344 174548
rect 165396 174536 165402 174548
rect 214650 174536 214656 174548
rect 165396 174508 214656 174536
rect 165396 174496 165402 174508
rect 214650 174496 214656 174508
rect 214708 174496 214714 174548
rect 249242 174496 249248 174548
rect 249300 174536 249306 174548
rect 265894 174536 265900 174548
rect 249300 174508 265900 174536
rect 249300 174496 249306 174508
rect 265894 174496 265900 174508
rect 265952 174496 265958 174548
rect 229370 174156 229376 174208
rect 229428 174196 229434 174208
rect 229830 174196 229836 174208
rect 229428 174168 229836 174196
rect 229428 174156 229434 174168
rect 229830 174156 229836 174168
rect 229888 174156 229894 174208
rect 258902 174020 258908 174072
rect 258960 174060 258966 174072
rect 265802 174060 265808 174072
rect 258960 174032 265808 174060
rect 258960 174020 258966 174032
rect 265802 174020 265808 174032
rect 265860 174020 265866 174072
rect 256142 173952 256148 174004
rect 256200 173992 256206 174004
rect 265986 173992 265992 174004
rect 256200 173964 265992 173992
rect 256200 173952 256206 173964
rect 265986 173952 265992 173964
rect 266044 173952 266050 174004
rect 241054 173884 241060 173936
rect 241112 173924 241118 173936
rect 264422 173924 264428 173936
rect 241112 173896 264428 173924
rect 241112 173884 241118 173896
rect 264422 173884 264428 173896
rect 264480 173884 264486 173936
rect 165522 173816 165528 173868
rect 165580 173856 165586 173868
rect 213914 173856 213920 173868
rect 165580 173828 213920 173856
rect 165580 173816 165586 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 231118 173816 231124 173868
rect 231176 173856 231182 173868
rect 251542 173856 251548 173868
rect 231176 173828 251548 173856
rect 231176 173816 231182 173828
rect 251542 173816 251548 173828
rect 251600 173816 251606 173868
rect 165706 173748 165712 173800
rect 165764 173788 165770 173800
rect 214006 173788 214012 173800
rect 165764 173760 214012 173788
rect 165764 173748 165770 173760
rect 214006 173748 214012 173760
rect 214064 173748 214070 173800
rect 231486 173748 231492 173800
rect 231544 173788 231550 173800
rect 244734 173788 244740 173800
rect 231544 173760 244740 173788
rect 231544 173748 231550 173760
rect 244734 173748 244740 173760
rect 244792 173748 244798 173800
rect 263318 172864 263324 172916
rect 263376 172904 263382 172916
rect 266078 172904 266084 172916
rect 263376 172876 266084 172904
rect 263376 172864 263382 172876
rect 266078 172864 266084 172876
rect 266136 172864 266142 172916
rect 253474 172660 253480 172712
rect 253532 172700 253538 172712
rect 265802 172700 265808 172712
rect 253532 172672 265808 172700
rect 253532 172660 253538 172672
rect 265802 172660 265808 172672
rect 265860 172660 265866 172712
rect 252094 172592 252100 172644
rect 252152 172632 252158 172644
rect 265986 172632 265992 172644
rect 252152 172604 265992 172632
rect 252152 172592 252158 172604
rect 265986 172592 265992 172604
rect 266044 172592 266050 172644
rect 250806 172524 250812 172576
rect 250864 172564 250870 172576
rect 265894 172564 265900 172576
rect 250864 172536 265900 172564
rect 250864 172524 250870 172536
rect 265894 172524 265900 172536
rect 265952 172524 265958 172576
rect 165430 172456 165436 172508
rect 165488 172496 165494 172508
rect 214006 172496 214012 172508
rect 165488 172468 214012 172496
rect 165488 172456 165494 172468
rect 214006 172456 214012 172468
rect 214064 172456 214070 172508
rect 231762 172456 231768 172508
rect 231820 172496 231826 172508
rect 244826 172496 244832 172508
rect 231820 172468 244832 172496
rect 231820 172456 231826 172468
rect 244826 172456 244832 172468
rect 244884 172456 244890 172508
rect 165798 172388 165804 172440
rect 165856 172428 165862 172440
rect 213914 172428 213920 172440
rect 165856 172400 213920 172428
rect 165856 172388 165862 172400
rect 213914 172388 213920 172400
rect 213972 172388 213978 172440
rect 231486 172388 231492 172440
rect 231544 172428 231550 172440
rect 245010 172428 245016 172440
rect 231544 172400 245016 172428
rect 231544 172388 231550 172400
rect 245010 172388 245016 172400
rect 245068 172388 245074 172440
rect 231670 172320 231676 172372
rect 231728 172360 231734 172372
rect 239398 172360 239404 172372
rect 231728 172332 239404 172360
rect 231728 172320 231734 172332
rect 239398 172320 239404 172332
rect 239456 172320 239462 172372
rect 231394 171300 231400 171352
rect 231452 171340 231458 171352
rect 231670 171340 231676 171352
rect 231452 171312 231676 171340
rect 231452 171300 231458 171312
rect 231670 171300 231676 171312
rect 231728 171300 231734 171352
rect 256234 171232 256240 171284
rect 256292 171272 256298 171284
rect 265250 171272 265256 171284
rect 256292 171244 265256 171272
rect 256292 171232 256298 171244
rect 265250 171232 265256 171244
rect 265308 171232 265314 171284
rect 251818 171164 251824 171216
rect 251876 171204 251882 171216
rect 265434 171204 265440 171216
rect 251876 171176 265440 171204
rect 251876 171164 251882 171176
rect 265434 171164 265440 171176
rect 265492 171164 265498 171216
rect 250714 171096 250720 171148
rect 250772 171136 250778 171148
rect 265526 171136 265532 171148
rect 250772 171108 265532 171136
rect 250772 171096 250778 171108
rect 265526 171096 265532 171108
rect 265584 171096 265590 171148
rect 166534 171028 166540 171080
rect 166592 171068 166598 171080
rect 213914 171068 213920 171080
rect 166592 171040 213920 171068
rect 166592 171028 166598 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 231762 171028 231768 171080
rect 231820 171068 231826 171080
rect 248782 171068 248788 171080
rect 231820 171040 248788 171068
rect 231820 171028 231826 171040
rect 248782 171028 248788 171040
rect 248840 171028 248846 171080
rect 231026 170688 231032 170740
rect 231084 170728 231090 170740
rect 231084 170700 231164 170728
rect 231084 170688 231090 170700
rect 231136 170536 231164 170700
rect 231118 170484 231124 170536
rect 231176 170484 231182 170536
rect 231210 170484 231216 170536
rect 231268 170524 231274 170536
rect 233234 170524 233240 170536
rect 231268 170496 233240 170524
rect 231268 170484 231274 170496
rect 233234 170484 233240 170496
rect 233292 170484 233298 170536
rect 167822 170348 167828 170400
rect 167880 170388 167886 170400
rect 214742 170388 214748 170400
rect 167880 170360 214748 170388
rect 167880 170348 167886 170360
rect 214742 170348 214748 170360
rect 214800 170348 214806 170400
rect 229738 170076 229744 170128
rect 229796 170116 229802 170128
rect 230750 170116 230756 170128
rect 229796 170088 230756 170116
rect 229796 170076 229802 170088
rect 230750 170076 230756 170088
rect 230808 170076 230814 170128
rect 253382 169872 253388 169924
rect 253440 169912 253446 169924
rect 265802 169912 265808 169924
rect 253440 169884 265808 169912
rect 253440 169872 253446 169884
rect 265802 169872 265808 169884
rect 265860 169872 265866 169924
rect 249426 169804 249432 169856
rect 249484 169844 249490 169856
rect 265526 169844 265532 169856
rect 249484 169816 265532 169844
rect 249484 169804 249490 169816
rect 265526 169804 265532 169816
rect 265584 169804 265590 169856
rect 235626 169736 235632 169788
rect 235684 169776 235690 169788
rect 265158 169776 265164 169788
rect 235684 169748 265164 169776
rect 235684 169736 235690 169748
rect 265158 169736 265164 169748
rect 265216 169736 265222 169788
rect 166442 169668 166448 169720
rect 166500 169708 166506 169720
rect 214006 169708 214012 169720
rect 166500 169680 214012 169708
rect 166500 169668 166506 169680
rect 214006 169668 214012 169680
rect 214064 169668 214070 169720
rect 231762 169668 231768 169720
rect 231820 169708 231826 169720
rect 247218 169708 247224 169720
rect 231820 169680 247224 169708
rect 231820 169668 231826 169680
rect 247218 169668 247224 169680
rect 247276 169668 247282 169720
rect 166350 169600 166356 169652
rect 166408 169640 166414 169652
rect 213914 169640 213920 169652
rect 166408 169612 213920 169640
rect 166408 169600 166414 169612
rect 213914 169600 213920 169612
rect 213972 169600 213978 169652
rect 259086 168512 259092 168564
rect 259144 168552 259150 168564
rect 265894 168552 265900 168564
rect 259144 168524 265900 168552
rect 259144 168512 259150 168524
rect 265894 168512 265900 168524
rect 265952 168512 265958 168564
rect 257522 168444 257528 168496
rect 257580 168484 257586 168496
rect 265802 168484 265808 168496
rect 257580 168456 265808 168484
rect 257580 168444 257586 168456
rect 265802 168444 265808 168456
rect 265860 168444 265866 168496
rect 238294 168376 238300 168428
rect 238352 168416 238358 168428
rect 265986 168416 265992 168428
rect 238352 168388 265992 168416
rect 238352 168376 238358 168388
rect 265986 168376 265992 168388
rect 266044 168376 266050 168428
rect 169386 168308 169392 168360
rect 169444 168348 169450 168360
rect 213914 168348 213920 168360
rect 169444 168320 213920 168348
rect 169444 168308 169450 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 231762 168308 231768 168360
rect 231820 168348 231826 168360
rect 248690 168348 248696 168360
rect 231820 168320 248696 168348
rect 231820 168308 231826 168320
rect 248690 168308 248696 168320
rect 248748 168308 248754 168360
rect 170674 168240 170680 168292
rect 170732 168280 170738 168292
rect 214006 168280 214012 168292
rect 170732 168252 214012 168280
rect 170732 168240 170738 168252
rect 214006 168240 214012 168252
rect 214064 168240 214070 168292
rect 231486 168240 231492 168292
rect 231544 168280 231550 168292
rect 247310 168280 247316 168292
rect 231544 168252 247316 168280
rect 231544 168240 231550 168252
rect 247310 168240 247316 168252
rect 247368 168240 247374 168292
rect 231394 168172 231400 168224
rect 231452 168212 231458 168224
rect 243998 168212 244004 168224
rect 231452 168184 244004 168212
rect 231452 168172 231458 168184
rect 243998 168172 244004 168184
rect 244056 168172 244062 168224
rect 280890 167560 280896 167612
rect 280948 167600 280954 167612
rect 282546 167600 282552 167612
rect 280948 167572 282552 167600
rect 280948 167560 280954 167572
rect 282546 167560 282552 167572
rect 282604 167560 282610 167612
rect 242434 167084 242440 167136
rect 242492 167124 242498 167136
rect 265802 167124 265808 167136
rect 242492 167096 265808 167124
rect 242492 167084 242498 167096
rect 265802 167084 265808 167096
rect 265860 167084 265866 167136
rect 238110 167016 238116 167068
rect 238168 167056 238174 167068
rect 265342 167056 265348 167068
rect 238168 167028 265348 167056
rect 238168 167016 238174 167028
rect 265342 167016 265348 167028
rect 265400 167016 265406 167068
rect 167730 166948 167736 167000
rect 167788 166988 167794 167000
rect 213914 166988 213920 167000
rect 167788 166960 213920 166988
rect 167788 166948 167794 166960
rect 213914 166948 213920 166960
rect 213972 166948 213978 167000
rect 291838 166948 291844 167000
rect 291896 166988 291902 167000
rect 580166 166988 580172 167000
rect 291896 166960 580172 166988
rect 291896 166948 291902 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 174630 166880 174636 166932
rect 174688 166920 174694 166932
rect 214006 166920 214012 166932
rect 174688 166892 214012 166920
rect 174688 166880 174694 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 191098 166812 191104 166864
rect 191156 166852 191162 166864
rect 214098 166852 214104 166864
rect 191156 166824 214104 166852
rect 191156 166812 191162 166824
rect 214098 166812 214104 166824
rect 214156 166812 214162 166864
rect 231302 166676 231308 166728
rect 231360 166716 231366 166728
rect 235258 166716 235264 166728
rect 231360 166688 235264 166716
rect 231360 166676 231366 166688
rect 235258 166676 235264 166688
rect 235316 166676 235322 166728
rect 231762 166608 231768 166660
rect 231820 166648 231826 166660
rect 234706 166648 234712 166660
rect 231820 166620 234712 166648
rect 231820 166608 231826 166620
rect 234706 166608 234712 166620
rect 234764 166608 234770 166660
rect 240962 166268 240968 166320
rect 241020 166308 241026 166320
rect 265158 166308 265164 166320
rect 241020 166280 265164 166308
rect 241020 166268 241026 166280
rect 265158 166268 265164 166280
rect 265216 166268 265222 166320
rect 231762 165724 231768 165776
rect 231820 165764 231826 165776
rect 234982 165764 234988 165776
rect 231820 165736 234988 165764
rect 231820 165724 231826 165736
rect 234982 165724 234988 165736
rect 235040 165724 235046 165776
rect 249150 165724 249156 165776
rect 249208 165764 249214 165776
rect 265802 165764 265808 165776
rect 249208 165736 265808 165764
rect 249208 165724 249214 165736
rect 265802 165724 265808 165736
rect 265860 165724 265866 165776
rect 254670 165656 254676 165708
rect 254728 165696 254734 165708
rect 265434 165696 265440 165708
rect 254728 165668 265440 165696
rect 254728 165656 254734 165668
rect 265434 165656 265440 165668
rect 265492 165656 265498 165708
rect 170582 165520 170588 165572
rect 170640 165560 170646 165572
rect 214006 165560 214012 165572
rect 170640 165532 214012 165560
rect 170640 165520 170646 165532
rect 214006 165520 214012 165532
rect 214064 165520 214070 165572
rect 231762 165520 231768 165572
rect 231820 165560 231826 165572
rect 240870 165560 240876 165572
rect 231820 165532 240876 165560
rect 231820 165520 231826 165532
rect 240870 165520 240876 165532
rect 240928 165520 240934 165572
rect 202138 165452 202144 165504
rect 202196 165492 202202 165504
rect 213914 165492 213920 165504
rect 202196 165464 213920 165492
rect 202196 165452 202202 165464
rect 213914 165452 213920 165464
rect 213972 165452 213978 165504
rect 231762 164908 231768 164960
rect 231820 164948 231826 164960
rect 234614 164948 234620 164960
rect 231820 164920 234620 164948
rect 231820 164908 231826 164920
rect 234614 164908 234620 164920
rect 234672 164908 234678 164960
rect 231394 164772 231400 164824
rect 231452 164812 231458 164824
rect 233786 164812 233792 164824
rect 231452 164784 233792 164812
rect 231452 164772 231458 164784
rect 233786 164772 233792 164784
rect 233844 164772 233850 164824
rect 263226 164364 263232 164416
rect 263284 164404 263290 164416
rect 265802 164404 265808 164416
rect 263284 164376 265808 164404
rect 263284 164364 263290 164376
rect 265802 164364 265808 164376
rect 265860 164364 265866 164416
rect 254578 164296 254584 164348
rect 254636 164336 254642 164348
rect 265894 164336 265900 164348
rect 254636 164308 265900 164336
rect 254636 164296 254642 164308
rect 265894 164296 265900 164308
rect 265952 164296 265958 164348
rect 249518 164228 249524 164280
rect 249576 164268 249582 164280
rect 265434 164268 265440 164280
rect 249576 164240 265440 164268
rect 249576 164228 249582 164240
rect 265434 164228 265440 164240
rect 265492 164228 265498 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 18598 164200 18604 164212
rect 3292 164172 18604 164200
rect 3292 164160 3298 164172
rect 18598 164160 18604 164172
rect 18656 164160 18662 164212
rect 169294 164160 169300 164212
rect 169352 164200 169358 164212
rect 213914 164200 213920 164212
rect 169352 164172 213920 164200
rect 169352 164160 169358 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 231486 164160 231492 164212
rect 231544 164200 231550 164212
rect 244918 164200 244924 164212
rect 231544 164172 244924 164200
rect 231544 164160 231550 164172
rect 244918 164160 244924 164172
rect 244976 164160 244982 164212
rect 173250 164092 173256 164144
rect 173308 164132 173314 164144
rect 214006 164132 214012 164144
rect 173308 164104 214012 164132
rect 173308 164092 173314 164104
rect 214006 164092 214012 164104
rect 214064 164092 214070 164144
rect 231394 163820 231400 163872
rect 231452 163860 231458 163872
rect 233970 163860 233976 163872
rect 231452 163832 233976 163860
rect 231452 163820 231458 163832
rect 233970 163820 233976 163832
rect 234028 163820 234034 163872
rect 231762 163412 231768 163464
rect 231820 163452 231826 163464
rect 235074 163452 235080 163464
rect 231820 163424 235080 163452
rect 231820 163412 231826 163424
rect 235074 163412 235080 163424
rect 235132 163412 235138 163464
rect 239490 163072 239496 163124
rect 239548 163112 239554 163124
rect 265158 163112 265164 163124
rect 239548 163084 265164 163112
rect 239548 163072 239554 163084
rect 265158 163072 265164 163084
rect 265216 163072 265222 163124
rect 260098 162936 260104 162988
rect 260156 162976 260162 162988
rect 265802 162976 265808 162988
rect 260156 162948 265808 162976
rect 260156 162936 260162 162948
rect 265802 162936 265808 162948
rect 265860 162936 265866 162988
rect 169202 162800 169208 162852
rect 169260 162840 169266 162852
rect 213914 162840 213920 162852
rect 169260 162812 213920 162840
rect 169260 162800 169266 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 280798 162800 280804 162852
rect 280856 162840 280862 162852
rect 281534 162840 281540 162852
rect 280856 162812 281540 162840
rect 280856 162800 280862 162812
rect 281534 162800 281540 162812
rect 281592 162800 281598 162852
rect 192478 162732 192484 162784
rect 192536 162772 192542 162784
rect 214006 162772 214012 162784
rect 192536 162744 214012 162772
rect 192536 162732 192542 162744
rect 214006 162732 214012 162744
rect 214064 162732 214070 162784
rect 260558 161712 260564 161764
rect 260616 161752 260622 161764
rect 265434 161752 265440 161764
rect 260616 161724 265440 161752
rect 260616 161712 260622 161724
rect 265434 161712 265440 161724
rect 265492 161712 265498 161764
rect 256418 161440 256424 161492
rect 256476 161480 256482 161492
rect 265802 161480 265808 161492
rect 256476 161452 265808 161480
rect 256476 161440 256482 161452
rect 265802 161440 265808 161452
rect 265860 161440 265866 161492
rect 174538 161372 174544 161424
rect 174596 161412 174602 161424
rect 213914 161412 213920 161424
rect 174596 161384 213920 161412
rect 174596 161372 174602 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 231762 161372 231768 161424
rect 231820 161412 231826 161424
rect 248598 161412 248604 161424
rect 231820 161384 248604 161412
rect 231820 161372 231826 161384
rect 248598 161372 248604 161384
rect 248656 161372 248662 161424
rect 282178 161168 282184 161220
rect 282236 161208 282242 161220
rect 285858 161208 285864 161220
rect 282236 161180 285864 161208
rect 282236 161168 282242 161180
rect 285858 161168 285864 161180
rect 285916 161168 285922 161220
rect 231762 160556 231768 160608
rect 231820 160596 231826 160608
rect 234430 160596 234436 160608
rect 231820 160568 234436 160596
rect 231820 160556 231826 160568
rect 234430 160556 234436 160568
rect 234488 160556 234494 160608
rect 257706 160216 257712 160268
rect 257764 160256 257770 160268
rect 265526 160256 265532 160268
rect 257764 160228 265532 160256
rect 257764 160216 257770 160228
rect 265526 160216 265532 160228
rect 265584 160216 265590 160268
rect 250622 160148 250628 160200
rect 250680 160188 250686 160200
rect 265986 160188 265992 160200
rect 250680 160160 265992 160188
rect 250680 160148 250686 160160
rect 265986 160148 265992 160160
rect 266044 160148 266050 160200
rect 241146 160080 241152 160132
rect 241204 160120 241210 160132
rect 242158 160120 242164 160132
rect 241204 160092 242164 160120
rect 241204 160080 241210 160092
rect 242158 160080 242164 160092
rect 242216 160080 242222 160132
rect 242250 160080 242256 160132
rect 242308 160120 242314 160132
rect 265894 160120 265900 160132
rect 242308 160092 265900 160120
rect 242308 160080 242314 160092
rect 265894 160080 265900 160092
rect 265952 160080 265958 160132
rect 167638 160012 167644 160064
rect 167696 160052 167702 160064
rect 214006 160052 214012 160064
rect 167696 160024 214012 160052
rect 167696 160012 167702 160024
rect 214006 160012 214012 160024
rect 214064 160012 214070 160064
rect 175918 159944 175924 159996
rect 175976 159984 175982 159996
rect 213914 159984 213920 159996
rect 175976 159956 213920 159984
rect 175976 159944 175982 159956
rect 213914 159944 213920 159956
rect 213972 159944 213978 159996
rect 231210 159944 231216 159996
rect 231268 159984 231274 159996
rect 240778 159984 240784 159996
rect 231268 159956 240784 159984
rect 231268 159944 231274 159956
rect 240778 159944 240784 159956
rect 240836 159944 240842 159996
rect 231762 159876 231768 159928
rect 231820 159916 231826 159928
rect 244550 159916 244556 159928
rect 231820 159888 244556 159916
rect 231820 159876 231826 159888
rect 244550 159876 244556 159888
rect 244608 159876 244614 159928
rect 230658 159740 230664 159792
rect 230716 159780 230722 159792
rect 232314 159780 232320 159792
rect 230716 159752 232320 159780
rect 230716 159740 230722 159752
rect 232314 159740 232320 159752
rect 232372 159740 232378 159792
rect 264606 159264 264612 159316
rect 264664 159304 264670 159316
rect 266262 159304 266268 159316
rect 264664 159276 266268 159304
rect 264664 159264 264670 159276
rect 266262 159264 266268 159276
rect 266320 159264 266326 159316
rect 282822 159128 282828 159180
rect 282880 159168 282886 159180
rect 287514 159168 287520 159180
rect 282880 159140 287520 159168
rect 282880 159128 282886 159140
rect 287514 159128 287520 159140
rect 287572 159128 287578 159180
rect 235350 158788 235356 158840
rect 235408 158828 235414 158840
rect 265434 158828 265440 158840
rect 235408 158800 265440 158828
rect 235408 158788 235414 158800
rect 265434 158788 265440 158800
rect 265492 158788 265498 158840
rect 235534 158720 235540 158772
rect 235592 158760 235598 158772
rect 265894 158760 265900 158772
rect 235592 158732 265900 158760
rect 235592 158720 235598 158732
rect 265894 158720 265900 158732
rect 265952 158720 265958 158772
rect 173158 158652 173164 158704
rect 173216 158692 173222 158704
rect 213914 158692 213920 158704
rect 173216 158664 213920 158692
rect 173216 158652 173222 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 231762 158652 231768 158704
rect 231820 158692 231826 158704
rect 251358 158692 251364 158704
rect 231820 158664 251364 158692
rect 231820 158652 231826 158664
rect 251358 158652 251364 158664
rect 251416 158652 251422 158704
rect 231026 158312 231032 158364
rect 231084 158352 231090 158364
rect 233694 158352 233700 158364
rect 231084 158324 233700 158352
rect 231084 158312 231090 158324
rect 233694 158312 233700 158324
rect 233752 158312 233758 158364
rect 238478 158040 238484 158092
rect 238536 158080 238542 158092
rect 266078 158080 266084 158092
rect 238536 158052 266084 158080
rect 238536 158040 238542 158052
rect 266078 158040 266084 158052
rect 266136 158040 266142 158092
rect 235442 157972 235448 158024
rect 235500 158012 235506 158024
rect 265342 158012 265348 158024
rect 235500 157984 265348 158012
rect 235500 157972 235506 157984
rect 265342 157972 265348 157984
rect 265400 157972 265406 158024
rect 281994 157904 282000 157956
rect 282052 157944 282058 157956
rect 284294 157944 284300 157956
rect 282052 157916 284300 157944
rect 282052 157904 282058 157916
rect 284294 157904 284300 157916
rect 284352 157904 284358 157956
rect 281902 157836 281908 157888
rect 281960 157876 281966 157888
rect 288802 157876 288808 157888
rect 281960 157848 288808 157876
rect 281960 157836 281966 157848
rect 288802 157836 288808 157848
rect 288860 157836 288866 157888
rect 259178 157428 259184 157480
rect 259236 157468 259242 157480
rect 265894 157468 265900 157480
rect 259236 157440 265900 157468
rect 259236 157428 259242 157440
rect 265894 157428 265900 157440
rect 265952 157428 265958 157480
rect 253658 157360 253664 157412
rect 253716 157400 253722 157412
rect 265802 157400 265808 157412
rect 253716 157372 265808 157400
rect 253716 157360 253722 157372
rect 265802 157360 265808 157372
rect 265860 157360 265866 157412
rect 169110 157292 169116 157344
rect 169168 157332 169174 157344
rect 214006 157332 214012 157344
rect 169168 157304 214012 157332
rect 169168 157292 169174 157304
rect 214006 157292 214012 157304
rect 214064 157292 214070 157344
rect 231762 157292 231768 157344
rect 231820 157332 231826 157344
rect 250162 157332 250168 157344
rect 231820 157304 250168 157332
rect 231820 157292 231826 157304
rect 250162 157292 250168 157304
rect 250220 157292 250226 157344
rect 282822 157292 282828 157344
rect 282880 157332 282886 157344
rect 292574 157332 292580 157344
rect 282880 157304 292580 157332
rect 282880 157292 282886 157304
rect 292574 157292 292580 157304
rect 292632 157292 292638 157344
rect 170490 157224 170496 157276
rect 170548 157264 170554 157276
rect 213914 157264 213920 157276
rect 170548 157236 213920 157264
rect 170548 157224 170554 157236
rect 213914 157224 213920 157236
rect 213972 157224 213978 157276
rect 231486 157224 231492 157276
rect 231544 157264 231550 157276
rect 244090 157264 244096 157276
rect 231544 157236 244096 157264
rect 231544 157224 231550 157236
rect 244090 157224 244096 157236
rect 244148 157224 244154 157276
rect 252278 156612 252284 156664
rect 252336 156652 252342 156664
rect 265158 156652 265164 156664
rect 252336 156624 265164 156652
rect 252336 156612 252342 156624
rect 265158 156612 265164 156624
rect 265216 156612 265222 156664
rect 282454 156544 282460 156596
rect 282512 156584 282518 156596
rect 285674 156584 285680 156596
rect 282512 156556 285680 156584
rect 282512 156544 282518 156556
rect 285674 156544 285680 156556
rect 285732 156544 285738 156596
rect 254946 156000 254952 156052
rect 255004 156040 255010 156052
rect 265894 156040 265900 156052
rect 255004 156012 265900 156040
rect 255004 156000 255010 156012
rect 265894 156000 265900 156012
rect 265952 156000 265958 156052
rect 240870 155932 240876 155984
rect 240928 155972 240934 155984
rect 265802 155972 265808 155984
rect 240928 155944 265808 155972
rect 240928 155932 240934 155944
rect 265802 155932 265808 155944
rect 265860 155932 265866 155984
rect 166258 155864 166264 155916
rect 166316 155904 166322 155916
rect 213914 155904 213920 155916
rect 166316 155876 213920 155904
rect 166316 155864 166322 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 230566 155864 230572 155916
rect 230624 155904 230630 155916
rect 250070 155904 250076 155916
rect 230624 155876 250076 155904
rect 230624 155864 230630 155876
rect 250070 155864 250076 155876
rect 250128 155864 250134 155916
rect 282822 155864 282828 155916
rect 282880 155904 282886 155916
rect 291286 155904 291292 155916
rect 282880 155876 291292 155904
rect 282880 155864 282886 155876
rect 291286 155864 291292 155876
rect 291344 155864 291350 155916
rect 170398 155796 170404 155848
rect 170456 155836 170462 155848
rect 214006 155836 214012 155848
rect 170456 155808 214012 155836
rect 170456 155796 170462 155808
rect 214006 155796 214012 155808
rect 214064 155796 214070 155848
rect 230474 155796 230480 155848
rect 230532 155836 230538 155848
rect 232222 155836 232228 155848
rect 230532 155808 232228 155836
rect 230532 155796 230538 155808
rect 232222 155796 232228 155808
rect 232280 155796 232286 155848
rect 282178 155728 282184 155780
rect 282236 155768 282242 155780
rect 283190 155768 283196 155780
rect 282236 155740 283196 155768
rect 282236 155728 282242 155740
rect 283190 155728 283196 155740
rect 283248 155728 283254 155780
rect 230474 155252 230480 155304
rect 230532 155292 230538 155304
rect 232130 155292 232136 155304
rect 230532 155264 232136 155292
rect 230532 155252 230538 155264
rect 232130 155252 232136 155264
rect 232188 155252 232194 155304
rect 260466 154708 260472 154760
rect 260524 154748 260530 154760
rect 265802 154748 265808 154760
rect 260524 154720 265808 154748
rect 260524 154708 260530 154720
rect 265802 154708 265808 154720
rect 265860 154708 265866 154760
rect 261754 154640 261760 154692
rect 261812 154680 261818 154692
rect 265526 154680 265532 154692
rect 261812 154652 265532 154680
rect 261812 154640 261818 154652
rect 265526 154640 265532 154652
rect 265584 154640 265590 154692
rect 250990 154572 250996 154624
rect 251048 154612 251054 154624
rect 265434 154612 265440 154624
rect 251048 154584 265440 154612
rect 251048 154572 251054 154584
rect 265434 154572 265440 154584
rect 265492 154572 265498 154624
rect 282086 154096 282092 154148
rect 282144 154136 282150 154148
rect 286410 154136 286416 154148
rect 282144 154108 286416 154136
rect 282144 154096 282150 154108
rect 286410 154096 286416 154108
rect 286468 154096 286474 154148
rect 230750 153824 230756 153876
rect 230808 153824 230814 153876
rect 230768 153672 230796 153824
rect 230750 153620 230756 153672
rect 230808 153620 230814 153672
rect 255958 153348 255964 153400
rect 256016 153388 256022 153400
rect 265802 153388 265808 153400
rect 256016 153360 265808 153388
rect 256016 153348 256022 153360
rect 265802 153348 265808 153360
rect 265860 153348 265866 153400
rect 166442 153280 166448 153332
rect 166500 153320 166506 153332
rect 214006 153320 214012 153332
rect 166500 153292 214012 153320
rect 166500 153280 166506 153292
rect 214006 153280 214012 153292
rect 214064 153280 214070 153332
rect 249058 153280 249064 153332
rect 249116 153320 249122 153332
rect 265526 153320 265532 153332
rect 249116 153292 265532 153320
rect 249116 153280 249122 153292
rect 265526 153280 265532 153292
rect 265584 153280 265590 153332
rect 282270 153280 282276 153332
rect 282328 153320 282334 153332
rect 286318 153320 286324 153332
rect 282328 153292 286324 153320
rect 282328 153280 282334 153292
rect 286318 153280 286324 153292
rect 286376 153280 286382 153332
rect 166258 153212 166264 153264
rect 166316 153252 166322 153264
rect 213914 153252 213920 153264
rect 166316 153224 213920 153252
rect 166316 153212 166322 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 242342 153212 242348 153264
rect 242400 153252 242406 153264
rect 264514 153252 264520 153264
rect 242400 153224 264520 153252
rect 242400 153212 242406 153224
rect 264514 153212 264520 153224
rect 264572 153212 264578 153264
rect 231762 153144 231768 153196
rect 231820 153184 231826 153196
rect 251450 153184 251456 153196
rect 231820 153156 251456 153184
rect 231820 153144 231826 153156
rect 251450 153144 251456 153156
rect 251508 153144 251514 153196
rect 282086 153144 282092 153196
rect 282144 153184 282150 153196
rect 292758 153184 292764 153196
rect 282144 153156 292764 153184
rect 282144 153144 282150 153156
rect 292758 153144 292764 153156
rect 292816 153144 292822 153196
rect 231118 153076 231124 153128
rect 231176 153116 231182 153128
rect 234890 153116 234896 153128
rect 231176 153088 234896 153116
rect 231176 153076 231182 153088
rect 234890 153076 234896 153088
rect 234948 153076 234954 153128
rect 231302 153008 231308 153060
rect 231360 153048 231366 153060
rect 236638 153048 236644 153060
rect 231360 153020 236644 153048
rect 231360 153008 231366 153020
rect 236638 153008 236644 153020
rect 236696 153008 236702 153060
rect 251910 151852 251916 151904
rect 251968 151892 251974 151904
rect 265250 151892 265256 151904
rect 251968 151864 265256 151892
rect 251968 151852 251974 151864
rect 265250 151852 265256 151864
rect 265308 151852 265314 151904
rect 166350 151784 166356 151836
rect 166408 151824 166414 151836
rect 213914 151824 213920 151836
rect 166408 151796 213920 151824
rect 166408 151784 166414 151796
rect 213914 151784 213920 151796
rect 213972 151784 213978 151836
rect 243630 151784 243636 151836
rect 243688 151824 243694 151836
rect 265802 151824 265808 151836
rect 243688 151796 265808 151824
rect 243688 151784 243694 151796
rect 265802 151784 265808 151796
rect 265860 151784 265866 151836
rect 282270 151716 282276 151768
rect 282328 151756 282334 151768
rect 285030 151756 285036 151768
rect 282328 151728 285036 151756
rect 282328 151716 282334 151728
rect 285030 151716 285036 151728
rect 285088 151716 285094 151768
rect 176010 151036 176016 151088
rect 176068 151076 176074 151088
rect 214834 151076 214840 151088
rect 176068 151048 214840 151076
rect 176068 151036 176074 151048
rect 214834 151036 214840 151048
rect 214892 151036 214898 151088
rect 257338 151036 257344 151088
rect 257396 151076 257402 151088
rect 265894 151076 265900 151088
rect 257396 151048 265900 151076
rect 257396 151036 257402 151048
rect 265894 151036 265900 151048
rect 265952 151036 265958 151088
rect 281626 150968 281632 151020
rect 281684 151008 281690 151020
rect 283558 151008 283564 151020
rect 281684 150980 283564 151008
rect 281684 150968 281690 150980
rect 283558 150968 283564 150980
rect 283616 150968 283622 151020
rect 236730 150560 236736 150612
rect 236788 150600 236794 150612
rect 265802 150600 265808 150612
rect 236788 150572 265808 150600
rect 236788 150560 236794 150572
rect 265802 150560 265808 150572
rect 265860 150560 265866 150612
rect 236822 150492 236828 150544
rect 236880 150532 236886 150544
rect 265342 150532 265348 150544
rect 236880 150504 265348 150532
rect 236880 150492 236886 150504
rect 265342 150492 265348 150504
rect 265400 150492 265406 150544
rect 173158 150424 173164 150476
rect 173216 150464 173222 150476
rect 214006 150464 214012 150476
rect 173216 150436 214012 150464
rect 173216 150424 173222 150436
rect 214006 150424 214012 150436
rect 214064 150424 214070 150476
rect 236638 150424 236644 150476
rect 236696 150464 236702 150476
rect 265066 150464 265072 150476
rect 236696 150436 265072 150464
rect 236696 150424 236702 150436
rect 265066 150424 265072 150436
rect 265124 150424 265130 150476
rect 169018 150356 169024 150408
rect 169076 150396 169082 150408
rect 213914 150396 213920 150408
rect 169076 150368 213920 150396
rect 169076 150356 169082 150368
rect 213914 150356 213920 150368
rect 213972 150356 213978 150408
rect 231762 150356 231768 150408
rect 231820 150396 231826 150408
rect 247126 150396 247132 150408
rect 231820 150368 247132 150396
rect 231820 150356 231826 150368
rect 247126 150356 247132 150368
rect 247184 150356 247190 150408
rect 230750 150288 230756 150340
rect 230808 150328 230814 150340
rect 233510 150328 233516 150340
rect 230808 150300 233516 150328
rect 230808 150288 230814 150300
rect 233510 150288 233516 150300
rect 233568 150288 233574 150340
rect 261662 149200 261668 149252
rect 261720 149240 261726 149252
rect 265342 149240 265348 149252
rect 261720 149212 265348 149240
rect 261720 149200 261726 149212
rect 265342 149200 265348 149212
rect 265400 149200 265406 149252
rect 282822 149200 282828 149252
rect 282880 149240 282886 149252
rect 288434 149240 288440 149252
rect 282880 149212 288440 149240
rect 282880 149200 282886 149212
rect 288434 149200 288440 149212
rect 288492 149200 288498 149252
rect 262858 149132 262864 149184
rect 262916 149172 262922 149184
rect 265802 149172 265808 149184
rect 262916 149144 265808 149172
rect 262916 149132 262922 149144
rect 265802 149132 265808 149144
rect 265860 149132 265866 149184
rect 235258 149064 235264 149116
rect 235316 149104 235322 149116
rect 265526 149104 265532 149116
rect 235316 149076 265532 149104
rect 235316 149064 235322 149076
rect 265526 149064 265532 149076
rect 265584 149064 265590 149116
rect 166626 148996 166632 149048
rect 166684 149036 166690 149048
rect 213914 149036 213920 149048
rect 166684 149008 213920 149036
rect 166684 148996 166690 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 231762 148996 231768 149048
rect 231820 149036 231826 149048
rect 249978 149036 249984 149048
rect 231820 149008 249984 149036
rect 231820 148996 231826 149008
rect 249978 148996 249984 149008
rect 250036 148996 250042 149048
rect 282822 148996 282828 149048
rect 282880 149036 282886 149048
rect 292666 149036 292672 149048
rect 282880 149008 292672 149036
rect 282880 148996 282886 149008
rect 292666 148996 292672 149008
rect 292724 148996 292730 149048
rect 282086 148860 282092 148912
rect 282144 148900 282150 148912
rect 284938 148900 284944 148912
rect 282144 148872 284944 148900
rect 282144 148860 282150 148872
rect 284938 148860 284944 148872
rect 284996 148860 285002 148912
rect 231210 148724 231216 148776
rect 231268 148764 231274 148776
rect 233418 148764 233424 148776
rect 231268 148736 233424 148764
rect 231268 148724 231274 148736
rect 233418 148724 233424 148736
rect 233476 148724 233482 148776
rect 233970 147704 233976 147756
rect 234028 147744 234034 147756
rect 266078 147744 266084 147756
rect 234028 147716 266084 147744
rect 234028 147704 234034 147716
rect 266078 147704 266084 147716
rect 266136 147704 266142 147756
rect 166534 147636 166540 147688
rect 166592 147676 166598 147688
rect 213914 147676 213920 147688
rect 166592 147648 213920 147676
rect 166592 147636 166598 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 233878 147636 233884 147688
rect 233936 147676 233942 147688
rect 265894 147676 265900 147688
rect 233936 147648 265900 147676
rect 233936 147636 233942 147648
rect 265894 147636 265900 147648
rect 265952 147636 265958 147688
rect 231762 147568 231768 147620
rect 231820 147608 231826 147620
rect 251266 147608 251272 147620
rect 231820 147580 251272 147608
rect 231820 147568 231826 147580
rect 251266 147568 251272 147580
rect 251324 147568 251330 147620
rect 230566 147092 230572 147144
rect 230624 147132 230630 147144
rect 232406 147132 232412 147144
rect 230624 147104 232412 147132
rect 230624 147092 230630 147104
rect 232406 147092 232412 147104
rect 232464 147092 232470 147144
rect 245286 146888 245292 146940
rect 245344 146928 245350 146940
rect 265802 146928 265808 146940
rect 245344 146900 265808 146928
rect 245344 146888 245350 146900
rect 265802 146888 265808 146900
rect 265860 146888 265866 146940
rect 258718 146412 258724 146464
rect 258776 146452 258782 146464
rect 265802 146452 265808 146464
rect 258776 146424 265808 146452
rect 258776 146412 258782 146424
rect 265802 146412 265808 146424
rect 265860 146412 265866 146464
rect 178678 146344 178684 146396
rect 178736 146384 178742 146396
rect 213914 146384 213920 146396
rect 178736 146356 213920 146384
rect 178736 146344 178742 146356
rect 213914 146344 213920 146356
rect 213972 146344 213978 146396
rect 254854 146344 254860 146396
rect 254912 146384 254918 146396
rect 265526 146384 265532 146396
rect 254912 146356 265532 146384
rect 254912 146344 254918 146356
rect 265526 146344 265532 146356
rect 265584 146344 265590 146396
rect 177298 146276 177304 146328
rect 177356 146316 177362 146328
rect 214006 146316 214012 146328
rect 177356 146288 214012 146316
rect 177356 146276 177362 146288
rect 214006 146276 214012 146288
rect 214064 146276 214070 146328
rect 232498 146276 232504 146328
rect 232556 146316 232562 146328
rect 265894 146316 265900 146328
rect 232556 146288 265900 146316
rect 232556 146276 232562 146288
rect 265894 146276 265900 146288
rect 265952 146276 265958 146328
rect 231302 146208 231308 146260
rect 231360 146248 231366 146260
rect 234798 146248 234804 146260
rect 231360 146220 234804 146248
rect 231360 146208 231366 146220
rect 234798 146208 234804 146220
rect 234856 146208 234862 146260
rect 231670 145596 231676 145648
rect 231728 145636 231734 145648
rect 241790 145636 241796 145648
rect 231728 145608 241796 145636
rect 231728 145596 231734 145608
rect 241790 145596 241796 145608
rect 241848 145596 241854 145648
rect 232682 145528 232688 145580
rect 232740 145568 232746 145580
rect 265250 145568 265256 145580
rect 232740 145540 265256 145568
rect 232740 145528 232746 145540
rect 265250 145528 265256 145540
rect 265308 145528 265314 145580
rect 256326 145052 256332 145104
rect 256384 145092 256390 145104
rect 265802 145092 265808 145104
rect 256384 145064 265808 145092
rect 256384 145052 256390 145064
rect 265802 145052 265808 145064
rect 265860 145052 265866 145104
rect 282822 145052 282828 145104
rect 282880 145092 282886 145104
rect 288710 145092 288716 145104
rect 282880 145064 288716 145092
rect 282880 145052 282886 145064
rect 288710 145052 288716 145064
rect 288768 145052 288774 145104
rect 184198 144984 184204 145036
rect 184256 145024 184262 145036
rect 214006 145024 214012 145036
rect 184256 144996 214012 145024
rect 184256 144984 184262 144996
rect 214006 144984 214012 144996
rect 214064 144984 214070 145036
rect 231118 144984 231124 145036
rect 231176 145024 231182 145036
rect 233602 145024 233608 145036
rect 231176 144996 233608 145024
rect 231176 144984 231182 144996
rect 233602 144984 233608 144996
rect 233660 144984 233666 145036
rect 250898 144984 250904 145036
rect 250956 145024 250962 145036
rect 265894 145024 265900 145036
rect 250956 144996 265900 145024
rect 250956 144984 250962 144996
rect 265894 144984 265900 144996
rect 265952 144984 265958 145036
rect 174538 144916 174544 144968
rect 174596 144956 174602 144968
rect 213914 144956 213920 144968
rect 174596 144928 213920 144956
rect 174596 144916 174602 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 242618 144916 242624 144968
rect 242676 144956 242682 144968
rect 265158 144956 265164 144968
rect 242676 144928 265164 144956
rect 242676 144916 242682 144928
rect 265158 144916 265164 144928
rect 265216 144916 265222 144968
rect 231302 144848 231308 144900
rect 231360 144888 231366 144900
rect 245102 144888 245108 144900
rect 231360 144860 245108 144888
rect 231360 144848 231366 144860
rect 245102 144848 245108 144860
rect 245160 144848 245166 144900
rect 231762 144780 231768 144832
rect 231820 144820 231826 144832
rect 241146 144820 241152 144832
rect 231820 144792 241152 144820
rect 231820 144780 231826 144792
rect 241146 144780 241152 144792
rect 241204 144780 241210 144832
rect 281902 144440 281908 144492
rect 281960 144480 281966 144492
rect 284386 144480 284392 144492
rect 281960 144452 284392 144480
rect 281960 144440 281966 144452
rect 284386 144440 284392 144452
rect 284444 144440 284450 144492
rect 241238 144168 241244 144220
rect 241296 144208 241302 144220
rect 265250 144208 265256 144220
rect 241296 144180 265256 144208
rect 241296 144168 241302 144180
rect 265250 144168 265256 144180
rect 265308 144168 265314 144220
rect 263134 143624 263140 143676
rect 263192 143664 263198 143676
rect 265802 143664 265808 143676
rect 263192 143636 265808 143664
rect 263192 143624 263198 143636
rect 265802 143624 265808 143636
rect 265860 143624 265866 143676
rect 202138 143556 202144 143608
rect 202196 143596 202202 143608
rect 213914 143596 213920 143608
rect 202196 143568 213920 143596
rect 202196 143556 202202 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 252186 143556 252192 143608
rect 252244 143596 252250 143608
rect 265342 143596 265348 143608
rect 252244 143568 265348 143596
rect 252244 143556 252250 143568
rect 265342 143556 265348 143568
rect 265400 143556 265406 143608
rect 231302 143488 231308 143540
rect 231360 143528 231366 143540
rect 245194 143528 245200 143540
rect 231360 143500 245200 143528
rect 231360 143488 231366 143500
rect 245194 143488 245200 143500
rect 245252 143488 245258 143540
rect 282822 143488 282828 143540
rect 282880 143528 282886 143540
rect 289906 143528 289912 143540
rect 282880 143500 289912 143528
rect 282880 143488 282886 143500
rect 289906 143488 289912 143500
rect 289964 143488 289970 143540
rect 231762 143420 231768 143472
rect 231820 143460 231826 143472
rect 238018 143460 238024 143472
rect 231820 143432 238024 143460
rect 231820 143420 231826 143432
rect 238018 143420 238024 143432
rect 238076 143420 238082 143472
rect 186958 142196 186964 142248
rect 187016 142236 187022 142248
rect 213914 142236 213920 142248
rect 187016 142208 213920 142236
rect 187016 142196 187022 142208
rect 213914 142196 213920 142208
rect 213972 142196 213978 142248
rect 181438 142128 181444 142180
rect 181496 142168 181502 142180
rect 214006 142168 214012 142180
rect 181496 142140 214012 142168
rect 181496 142128 181502 142140
rect 214006 142128 214012 142140
rect 214064 142128 214070 142180
rect 245194 142128 245200 142180
rect 245252 142168 245258 142180
rect 265158 142168 265164 142180
rect 245252 142140 265164 142168
rect 245252 142128 245258 142140
rect 265158 142128 265164 142140
rect 265216 142128 265222 142180
rect 231762 142060 231768 142112
rect 231820 142100 231826 142112
rect 248506 142100 248512 142112
rect 231820 142072 248512 142100
rect 231820 142060 231826 142072
rect 248506 142060 248512 142072
rect 248564 142060 248570 142112
rect 231394 141992 231400 142044
rect 231452 142032 231458 142044
rect 244366 142032 244372 142044
rect 231452 142004 244372 142032
rect 231452 141992 231458 142004
rect 244366 141992 244372 142004
rect 244424 141992 244430 142044
rect 231762 141652 231768 141704
rect 231820 141692 231826 141704
rect 235166 141692 235172 141704
rect 231820 141664 235172 141692
rect 231820 141652 231826 141664
rect 235166 141652 235172 141664
rect 235224 141652 235230 141704
rect 182818 140836 182824 140888
rect 182876 140876 182882 140888
rect 213914 140876 213920 140888
rect 182876 140848 213920 140876
rect 182876 140836 182882 140848
rect 213914 140836 213920 140848
rect 213972 140836 213978 140888
rect 244274 140836 244280 140888
rect 244332 140876 244338 140888
rect 265802 140876 265808 140888
rect 244332 140848 265808 140876
rect 244332 140836 244338 140848
rect 265802 140836 265808 140848
rect 265860 140836 265866 140888
rect 175918 140768 175924 140820
rect 175976 140808 175982 140820
rect 214006 140808 214012 140820
rect 175976 140780 214012 140808
rect 175976 140768 175982 140780
rect 214006 140768 214012 140780
rect 214064 140768 214070 140820
rect 232590 140768 232596 140820
rect 232648 140808 232654 140820
rect 265894 140808 265900 140820
rect 232648 140780 265900 140808
rect 232648 140768 232654 140780
rect 265894 140768 265900 140780
rect 265952 140768 265958 140820
rect 231762 140700 231768 140752
rect 231820 140740 231826 140752
rect 251174 140740 251180 140752
rect 231820 140712 251180 140740
rect 231820 140700 231826 140712
rect 251174 140700 251180 140712
rect 251232 140700 251238 140752
rect 231210 140632 231216 140684
rect 231268 140672 231274 140684
rect 249886 140672 249892 140684
rect 231268 140644 249892 140672
rect 231268 140632 231274 140644
rect 249886 140632 249892 140644
rect 249944 140632 249950 140684
rect 244274 140128 244280 140140
rect 231228 140100 244280 140128
rect 231228 140072 231256 140100
rect 244274 140088 244280 140100
rect 244332 140088 244338 140140
rect 231210 140020 231216 140072
rect 231268 140020 231274 140072
rect 234062 140020 234068 140072
rect 234120 140060 234126 140072
rect 266262 140060 266268 140072
rect 234120 140032 266268 140060
rect 234120 140020 234126 140032
rect 266262 140020 266268 140032
rect 266320 140020 266326 140072
rect 282822 139816 282828 139868
rect 282880 139856 282886 139868
rect 287422 139856 287428 139868
rect 282880 139828 287428 139856
rect 282880 139816 282886 139828
rect 287422 139816 287428 139828
rect 287480 139816 287486 139868
rect 258994 139544 259000 139596
rect 259052 139584 259058 139596
rect 265526 139584 265532 139596
rect 259052 139556 265532 139584
rect 259052 139544 259058 139556
rect 265526 139544 265532 139556
rect 265584 139544 265590 139596
rect 178770 139476 178776 139528
rect 178828 139516 178834 139528
rect 213914 139516 213920 139528
rect 178828 139488 213920 139516
rect 178828 139476 178834 139488
rect 213914 139476 213920 139488
rect 213972 139476 213978 139528
rect 246482 139476 246488 139528
rect 246540 139516 246546 139528
rect 265894 139516 265900 139528
rect 246540 139488 265900 139516
rect 246540 139476 246546 139488
rect 265894 139476 265900 139488
rect 265952 139476 265958 139528
rect 177390 139408 177396 139460
rect 177448 139448 177454 139460
rect 214006 139448 214012 139460
rect 177448 139420 214012 139448
rect 177448 139408 177454 139420
rect 214006 139408 214012 139420
rect 214064 139408 214070 139460
rect 243538 139408 243544 139460
rect 243596 139448 243602 139460
rect 265802 139448 265808 139460
rect 243596 139420 265808 139448
rect 243596 139408 243602 139420
rect 265802 139408 265808 139420
rect 265860 139408 265866 139460
rect 266170 139448 266176 139460
rect 265912 139420 266176 139448
rect 265912 139256 265940 139420
rect 266170 139408 266176 139420
rect 266228 139408 266234 139460
rect 282822 139340 282828 139392
rect 282880 139380 282886 139392
rect 289170 139380 289176 139392
rect 282880 139352 289176 139380
rect 282880 139340 282886 139352
rect 289170 139340 289176 139352
rect 289228 139340 289234 139392
rect 298738 139340 298744 139392
rect 298796 139380 298802 139392
rect 580166 139380 580172 139392
rect 298796 139352 580172 139380
rect 298796 139340 298802 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 265894 139204 265900 139256
rect 265952 139204 265958 139256
rect 231302 138796 231308 138848
rect 231360 138836 231366 138848
rect 234154 138836 234160 138848
rect 231360 138808 234160 138836
rect 231360 138796 231366 138808
rect 234154 138796 234160 138808
rect 234212 138796 234218 138848
rect 231118 138728 231124 138780
rect 231176 138768 231182 138780
rect 254578 138768 254584 138780
rect 231176 138740 254584 138768
rect 231176 138728 231182 138740
rect 254578 138728 254584 138740
rect 254636 138728 254642 138780
rect 238386 138660 238392 138712
rect 238444 138700 238450 138712
rect 261570 138700 261576 138712
rect 238444 138672 261576 138700
rect 238444 138660 238450 138672
rect 261570 138660 261576 138672
rect 261628 138660 261634 138712
rect 253198 138116 253204 138168
rect 253256 138156 253262 138168
rect 265434 138156 265440 138168
rect 253256 138128 265440 138156
rect 253256 138116 253262 138128
rect 265434 138116 265440 138128
rect 265492 138116 265498 138168
rect 252002 138048 252008 138100
rect 252060 138088 252066 138100
rect 265526 138088 265532 138100
rect 252060 138060 265532 138088
rect 252060 138048 252066 138060
rect 265526 138048 265532 138060
rect 265584 138048 265590 138100
rect 242158 137980 242164 138032
rect 242216 138020 242222 138032
rect 265986 138020 265992 138032
rect 242216 137992 265992 138020
rect 242216 137980 242222 137992
rect 265986 137980 265992 137992
rect 266044 137980 266050 138032
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 26878 137952 26884 137964
rect 3292 137924 26884 137952
rect 3292 137912 3298 137924
rect 26878 137912 26884 137924
rect 26936 137912 26942 137964
rect 231670 137912 231676 137964
rect 231728 137952 231734 137964
rect 249794 137952 249800 137964
rect 231728 137924 249800 137952
rect 231728 137912 231734 137924
rect 249794 137912 249800 137924
rect 249852 137912 249858 137964
rect 282270 137912 282276 137964
rect 282328 137952 282334 137964
rect 290182 137952 290188 137964
rect 282328 137924 290188 137952
rect 282328 137912 282334 137924
rect 290182 137912 290188 137924
rect 290240 137912 290246 137964
rect 231762 137844 231768 137896
rect 231820 137884 231826 137896
rect 247034 137884 247040 137896
rect 231820 137856 247040 137884
rect 231820 137844 231826 137856
rect 247034 137844 247040 137856
rect 247092 137844 247098 137896
rect 281626 137844 281632 137896
rect 281684 137884 281690 137896
rect 283466 137884 283472 137896
rect 281684 137856 283472 137884
rect 281684 137844 281690 137856
rect 283466 137844 283472 137856
rect 283524 137844 283530 137896
rect 170674 137232 170680 137284
rect 170732 137272 170738 137284
rect 214742 137272 214748 137284
rect 170732 137244 214748 137272
rect 170732 137232 170738 137244
rect 214742 137232 214748 137244
rect 214800 137232 214806 137284
rect 231302 137232 231308 137284
rect 231360 137272 231366 137284
rect 249518 137272 249524 137284
rect 231360 137244 249524 137272
rect 231360 137232 231366 137244
rect 249518 137232 249524 137244
rect 249576 137232 249582 137284
rect 250438 136756 250444 136808
rect 250496 136796 250502 136808
rect 265526 136796 265532 136808
rect 250496 136768 265532 136796
rect 250496 136756 250502 136768
rect 265526 136756 265532 136768
rect 265584 136756 265590 136808
rect 249334 136688 249340 136740
rect 249392 136728 249398 136740
rect 265986 136728 265992 136740
rect 249392 136700 265992 136728
rect 249392 136688 249398 136700
rect 265986 136688 265992 136700
rect 266044 136688 266050 136740
rect 170398 136620 170404 136672
rect 170456 136660 170462 136672
rect 213914 136660 213920 136672
rect 170456 136632 213920 136660
rect 170456 136620 170462 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 229922 136620 229928 136672
rect 229980 136660 229986 136672
rect 265434 136660 265440 136672
rect 229980 136632 265440 136660
rect 229980 136620 229986 136632
rect 265434 136620 265440 136632
rect 265492 136620 265498 136672
rect 231394 136552 231400 136604
rect 231452 136592 231458 136604
rect 263318 136592 263324 136604
rect 231452 136564 263324 136592
rect 231452 136552 231458 136564
rect 263318 136552 263324 136564
rect 263376 136552 263382 136604
rect 280982 136552 280988 136604
rect 281040 136592 281046 136604
rect 281626 136592 281632 136604
rect 281040 136564 281632 136592
rect 281040 136552 281046 136564
rect 281626 136552 281632 136564
rect 281684 136552 281690 136604
rect 282822 136552 282828 136604
rect 282880 136592 282886 136604
rect 290274 136592 290280 136604
rect 282880 136564 290280 136592
rect 282880 136552 282886 136564
rect 290274 136552 290280 136564
rect 290332 136552 290338 136604
rect 231762 136484 231768 136536
rect 231820 136524 231826 136536
rect 256142 136524 256148 136536
rect 231820 136496 256148 136524
rect 231820 136484 231826 136496
rect 256142 136484 256148 136496
rect 256200 136484 256206 136536
rect 240778 135464 240784 135516
rect 240836 135504 240842 135516
rect 265250 135504 265256 135516
rect 240836 135476 265256 135504
rect 240836 135464 240842 135476
rect 265250 135464 265256 135476
rect 265308 135464 265314 135516
rect 191098 135396 191104 135448
rect 191156 135436 191162 135448
rect 214006 135436 214012 135448
rect 191156 135408 214012 135436
rect 191156 135396 191162 135408
rect 214006 135396 214012 135408
rect 214064 135396 214070 135448
rect 260374 135396 260380 135448
rect 260432 135436 260438 135448
rect 264514 135436 264520 135448
rect 260432 135408 264520 135436
rect 260432 135396 260438 135408
rect 264514 135396 264520 135408
rect 264572 135396 264578 135448
rect 174630 135328 174636 135380
rect 174688 135368 174694 135380
rect 213914 135368 213920 135380
rect 174688 135340 213920 135368
rect 174688 135328 174694 135340
rect 213914 135328 213920 135340
rect 213972 135328 213978 135380
rect 256050 135328 256056 135380
rect 256108 135368 256114 135380
rect 262582 135368 262588 135380
rect 256108 135340 262588 135368
rect 256108 135328 256114 135340
rect 262582 135328 262588 135340
rect 262640 135328 262646 135380
rect 167638 135260 167644 135312
rect 167696 135300 167702 135312
rect 214098 135300 214104 135312
rect 167696 135272 214104 135300
rect 167696 135260 167702 135272
rect 214098 135260 214104 135272
rect 214156 135260 214162 135312
rect 263042 135260 263048 135312
rect 263100 135300 263106 135312
rect 265986 135300 265992 135312
rect 263100 135272 265992 135300
rect 263100 135260 263106 135272
rect 265986 135260 265992 135272
rect 266044 135260 266050 135312
rect 231670 135192 231676 135244
rect 231728 135232 231734 135244
rect 258902 135232 258908 135244
rect 231728 135204 258908 135232
rect 231728 135192 231734 135204
rect 258902 135192 258908 135204
rect 258960 135192 258966 135244
rect 231578 135124 231584 135176
rect 231636 135164 231642 135176
rect 252094 135164 252100 135176
rect 231636 135136 252100 135164
rect 231636 135124 231642 135136
rect 252094 135124 252100 135136
rect 252152 135124 252158 135176
rect 281810 135124 281816 135176
rect 281868 135164 281874 135176
rect 283650 135164 283656 135176
rect 281868 135136 283656 135164
rect 281868 135124 281874 135136
rect 283650 135124 283656 135136
rect 283708 135124 283714 135176
rect 231762 135056 231768 135108
rect 231820 135096 231826 135108
rect 241054 135096 241060 135108
rect 231820 135068 241060 135096
rect 231820 135056 231826 135068
rect 241054 135056 241060 135068
rect 241112 135056 241118 135108
rect 258810 134036 258816 134088
rect 258868 134076 258874 134088
rect 265986 134076 265992 134088
rect 258868 134048 265992 134076
rect 258868 134036 258874 134048
rect 265986 134036 265992 134048
rect 266044 134036 266050 134088
rect 254578 133968 254584 134020
rect 254636 134008 254642 134020
rect 264514 134008 264520 134020
rect 254636 133980 264520 134008
rect 254636 133968 254642 133980
rect 264514 133968 264520 133980
rect 264572 133968 264578 134020
rect 167730 133900 167736 133952
rect 167788 133940 167794 133952
rect 213914 133940 213920 133952
rect 167788 133912 213920 133940
rect 167788 133900 167794 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 214466 133900 214472 133952
rect 214524 133940 214530 133952
rect 214650 133940 214656 133952
rect 214524 133912 214656 133940
rect 214524 133900 214530 133912
rect 214650 133900 214656 133912
rect 214708 133900 214714 133952
rect 229830 133900 229836 133952
rect 229888 133940 229894 133952
rect 265250 133940 265256 133952
rect 229888 133912 265256 133940
rect 229888 133900 229894 133912
rect 265250 133900 265256 133912
rect 265308 133900 265314 133952
rect 231670 133832 231676 133884
rect 231728 133872 231734 133884
rect 256234 133872 256240 133884
rect 231728 133844 256240 133872
rect 231728 133832 231734 133844
rect 256234 133832 256240 133844
rect 256292 133832 256298 133884
rect 282270 133832 282276 133884
rect 282328 133872 282334 133884
rect 286226 133872 286232 133884
rect 282328 133844 286232 133872
rect 282328 133832 282334 133844
rect 286226 133832 286232 133844
rect 286284 133832 286290 133884
rect 231762 133764 231768 133816
rect 231820 133804 231826 133816
rect 253474 133804 253480 133816
rect 231820 133776 253480 133804
rect 231820 133764 231826 133776
rect 253474 133764 253480 133776
rect 253532 133764 253538 133816
rect 230658 133696 230664 133748
rect 230716 133736 230722 133748
rect 250806 133736 250812 133748
rect 230716 133708 250812 133736
rect 230716 133696 230722 133708
rect 250806 133696 250812 133708
rect 250864 133696 250870 133748
rect 214558 133288 214564 133340
rect 214616 133288 214622 133340
rect 214576 133136 214604 133288
rect 214558 133084 214564 133136
rect 214616 133084 214622 133136
rect 261570 132608 261576 132660
rect 261628 132648 261634 132660
rect 265158 132648 265164 132660
rect 261628 132620 265164 132648
rect 261628 132608 261634 132620
rect 265158 132608 265164 132620
rect 265216 132608 265222 132660
rect 169202 132540 169208 132592
rect 169260 132580 169266 132592
rect 213914 132580 213920 132592
rect 169260 132552 213920 132580
rect 169260 132540 169266 132552
rect 213914 132540 213920 132552
rect 213972 132540 213978 132592
rect 257614 132540 257620 132592
rect 257672 132580 257678 132592
rect 265986 132580 265992 132592
rect 257672 132552 265992 132580
rect 257672 132540 257678 132552
rect 265986 132540 265992 132552
rect 266044 132540 266050 132592
rect 169294 132472 169300 132524
rect 169352 132512 169358 132524
rect 214006 132512 214012 132524
rect 169352 132484 214012 132512
rect 169352 132472 169358 132484
rect 214006 132472 214012 132484
rect 214064 132472 214070 132524
rect 242526 132472 242532 132524
rect 242584 132512 242590 132524
rect 266170 132512 266176 132524
rect 242584 132484 266176 132512
rect 242584 132472 242590 132484
rect 266170 132472 266176 132484
rect 266228 132472 266234 132524
rect 231762 132404 231768 132456
rect 231820 132444 231826 132456
rect 251818 132444 251824 132456
rect 231820 132416 251824 132444
rect 231820 132404 231826 132416
rect 251818 132404 251824 132416
rect 251876 132404 251882 132456
rect 282086 132404 282092 132456
rect 282144 132444 282150 132456
rect 291194 132444 291200 132456
rect 282144 132416 291200 132444
rect 282144 132404 282150 132416
rect 291194 132404 291200 132416
rect 291252 132404 291258 132456
rect 231670 132336 231676 132388
rect 231728 132376 231734 132388
rect 250714 132376 250720 132388
rect 231728 132348 250720 132376
rect 231728 132336 231734 132348
rect 250714 132336 250720 132348
rect 250772 132336 250778 132388
rect 282546 132336 282552 132388
rect 282604 132376 282610 132388
rect 285766 132376 285772 132388
rect 282604 132348 285772 132376
rect 282604 132336 282610 132348
rect 285766 132336 285772 132348
rect 285824 132336 285830 132388
rect 231578 132268 231584 132320
rect 231636 132308 231642 132320
rect 249426 132308 249432 132320
rect 231636 132280 249432 132308
rect 231636 132268 231642 132280
rect 249426 132268 249432 132280
rect 249484 132268 249490 132320
rect 250806 131248 250812 131300
rect 250864 131288 250870 131300
rect 265986 131288 265992 131300
rect 250864 131260 265992 131288
rect 250864 131248 250870 131260
rect 265986 131248 265992 131260
rect 266044 131248 266050 131300
rect 169386 131180 169392 131232
rect 169444 131220 169450 131232
rect 214006 131220 214012 131232
rect 169444 131192 214012 131220
rect 169444 131180 169450 131192
rect 214006 131180 214012 131192
rect 214064 131180 214070 131232
rect 253566 131180 253572 131232
rect 253624 131220 253630 131232
rect 266170 131220 266176 131232
rect 253624 131192 266176 131220
rect 253624 131180 253630 131192
rect 266170 131180 266176 131192
rect 266228 131180 266234 131232
rect 169110 131112 169116 131164
rect 169168 131152 169174 131164
rect 213914 131152 213920 131164
rect 169168 131124 213920 131152
rect 169168 131112 169174 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 230934 131044 230940 131096
rect 230992 131084 230998 131096
rect 259086 131084 259092 131096
rect 230992 131056 259092 131084
rect 230992 131044 230998 131056
rect 259086 131044 259092 131056
rect 259144 131044 259150 131096
rect 281902 131044 281908 131096
rect 281960 131084 281966 131096
rect 284478 131084 284484 131096
rect 281960 131056 284484 131084
rect 281960 131044 281966 131056
rect 284478 131044 284484 131056
rect 284536 131044 284542 131096
rect 231486 130976 231492 131028
rect 231544 131016 231550 131028
rect 253382 131016 253388 131028
rect 231544 130988 253388 131016
rect 231544 130976 231550 130988
rect 253382 130976 253388 130988
rect 253440 130976 253446 131028
rect 282086 130976 282092 131028
rect 282144 131016 282150 131028
rect 285122 131016 285128 131028
rect 282144 130988 285128 131016
rect 282144 130976 282150 130988
rect 285122 130976 285128 130988
rect 285180 130976 285186 131028
rect 231026 130772 231032 130824
rect 231084 130812 231090 130824
rect 235626 130812 235632 130824
rect 231084 130784 235632 130812
rect 231084 130772 231090 130784
rect 235626 130772 235632 130784
rect 235684 130772 235690 130824
rect 241054 129888 241060 129940
rect 241112 129928 241118 129940
rect 265986 129928 265992 129940
rect 241112 129900 265992 129928
rect 241112 129888 241118 129900
rect 265986 129888 265992 129900
rect 266044 129888 266050 129940
rect 180150 129820 180156 129872
rect 180208 129860 180214 129872
rect 213914 129860 213920 129872
rect 180208 129832 213920 129860
rect 180208 129820 180214 129832
rect 213914 129820 213920 129832
rect 213972 129820 213978 129872
rect 256234 129820 256240 129872
rect 256292 129860 256298 129872
rect 266170 129860 266176 129872
rect 256292 129832 266176 129860
rect 256292 129820 256298 129832
rect 266170 129820 266176 129832
rect 266228 129820 266234 129872
rect 171778 129752 171784 129804
rect 171836 129792 171842 129804
rect 214006 129792 214012 129804
rect 171836 129764 214012 129792
rect 171836 129752 171842 129764
rect 214006 129752 214012 129764
rect 214064 129752 214070 129804
rect 231762 129684 231768 129736
rect 231820 129724 231826 129736
rect 257522 129724 257528 129736
rect 231820 129696 257528 129724
rect 231820 129684 231826 129696
rect 257522 129684 257528 129696
rect 257580 129684 257586 129736
rect 282086 129616 282092 129668
rect 282144 129656 282150 129668
rect 284846 129656 284852 129668
rect 282144 129628 284852 129656
rect 282144 129616 282150 129628
rect 284846 129616 284852 129628
rect 284904 129616 284910 129668
rect 281902 129548 281908 129600
rect 281960 129588 281966 129600
rect 284662 129588 284668 129600
rect 281960 129560 284668 129588
rect 281960 129548 281966 129560
rect 284662 129548 284668 129560
rect 284720 129548 284726 129600
rect 231670 129480 231676 129532
rect 231728 129520 231734 129532
rect 238294 129520 238300 129532
rect 231728 129492 238300 129520
rect 231728 129480 231734 129492
rect 238294 129480 238300 129492
rect 238352 129480 238358 129532
rect 257430 128460 257436 128512
rect 257488 128500 257494 128512
rect 265986 128500 265992 128512
rect 257488 128472 265992 128500
rect 257488 128460 257494 128472
rect 265986 128460 265992 128472
rect 266044 128460 266050 128512
rect 173250 128392 173256 128444
rect 173308 128432 173314 128444
rect 213914 128432 213920 128444
rect 173308 128404 213920 128432
rect 173308 128392 173314 128404
rect 213914 128392 213920 128404
rect 213972 128392 213978 128444
rect 245102 128392 245108 128444
rect 245160 128432 245166 128444
rect 265342 128432 265348 128444
rect 245160 128404 265348 128432
rect 245160 128392 245166 128404
rect 265342 128392 265348 128404
rect 265400 128392 265406 128444
rect 169018 128324 169024 128376
rect 169076 128364 169082 128376
rect 214006 128364 214012 128376
rect 169076 128336 214012 128364
rect 169076 128324 169082 128336
rect 214006 128324 214012 128336
rect 214064 128324 214070 128376
rect 238202 128324 238208 128376
rect 238260 128364 238266 128376
rect 265526 128364 265532 128376
rect 238260 128336 265532 128364
rect 238260 128324 238266 128336
rect 265526 128324 265532 128336
rect 265584 128324 265590 128376
rect 265986 128324 265992 128376
rect 266044 128364 266050 128376
rect 266170 128364 266176 128376
rect 266044 128336 266176 128364
rect 266044 128324 266050 128336
rect 266170 128324 266176 128336
rect 266228 128324 266234 128376
rect 231578 128256 231584 128308
rect 231636 128296 231642 128308
rect 242434 128296 242440 128308
rect 231636 128268 242440 128296
rect 231636 128256 231642 128268
rect 242434 128256 242440 128268
rect 242492 128256 242498 128308
rect 231670 128188 231676 128240
rect 231728 128228 231734 128240
rect 238478 128228 238484 128240
rect 231728 128200 238484 128228
rect 231728 128188 231734 128200
rect 238478 128188 238484 128200
rect 238536 128188 238542 128240
rect 281902 128188 281908 128240
rect 281960 128228 281966 128240
rect 284570 128228 284576 128240
rect 281960 128200 284576 128228
rect 281960 128188 281966 128200
rect 284570 128188 284576 128200
rect 284628 128188 284634 128240
rect 231762 128120 231768 128172
rect 231820 128160 231826 128172
rect 238110 128160 238116 128172
rect 231820 128132 238116 128160
rect 231820 128120 231826 128132
rect 238110 128120 238116 128132
rect 238168 128120 238174 128172
rect 281902 127644 281908 127696
rect 281960 127684 281966 127696
rect 284754 127684 284760 127696
rect 281960 127656 284760 127684
rect 281960 127644 281966 127656
rect 284754 127644 284760 127656
rect 284812 127644 284818 127696
rect 247678 127100 247684 127152
rect 247736 127140 247742 127152
rect 264146 127140 264152 127152
rect 247736 127112 264152 127140
rect 247736 127100 247742 127112
rect 264146 127100 264152 127112
rect 264204 127100 264210 127152
rect 192478 127032 192484 127084
rect 192536 127072 192542 127084
rect 213914 127072 213920 127084
rect 192536 127044 213920 127072
rect 192536 127032 192542 127044
rect 213914 127032 213920 127044
rect 213972 127032 213978 127084
rect 245010 127032 245016 127084
rect 245068 127072 245074 127084
rect 265526 127072 265532 127084
rect 245068 127044 265532 127072
rect 245068 127032 245074 127044
rect 265526 127032 265532 127044
rect 265584 127032 265590 127084
rect 167822 126964 167828 127016
rect 167880 127004 167886 127016
rect 214006 127004 214012 127016
rect 167880 126976 214012 127004
rect 167880 126964 167886 126976
rect 214006 126964 214012 126976
rect 214064 126964 214070 127016
rect 239398 126964 239404 127016
rect 239456 127004 239462 127016
rect 266170 127004 266176 127016
rect 239456 126976 266176 127004
rect 239456 126964 239462 126976
rect 266170 126964 266176 126976
rect 266228 126964 266234 127016
rect 231578 126896 231584 126948
rect 231636 126936 231642 126948
rect 254670 126936 254676 126948
rect 231636 126908 254676 126936
rect 231636 126896 231642 126908
rect 254670 126896 254676 126908
rect 254728 126896 254734 126948
rect 454678 126896 454684 126948
rect 454736 126936 454742 126948
rect 580166 126936 580172 126948
rect 454736 126908 580172 126936
rect 454736 126896 454742 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 231762 126828 231768 126880
rect 231820 126868 231826 126880
rect 249150 126868 249156 126880
rect 231820 126840 249156 126868
rect 231820 126828 231826 126840
rect 249150 126828 249156 126840
rect 249208 126828 249214 126880
rect 231670 126760 231676 126812
rect 231728 126800 231734 126812
rect 240962 126800 240968 126812
rect 231728 126772 240968 126800
rect 231728 126760 231734 126772
rect 240962 126760 240968 126772
rect 241020 126760 241026 126812
rect 282822 126692 282828 126744
rect 282880 126732 282886 126744
rect 288618 126732 288624 126744
rect 282880 126704 288624 126732
rect 282880 126692 282886 126704
rect 288618 126692 288624 126704
rect 288676 126692 288682 126744
rect 230842 126216 230848 126268
rect 230900 126256 230906 126268
rect 263226 126256 263232 126268
rect 230900 126228 263232 126256
rect 230900 126216 230906 126228
rect 263226 126216 263232 126228
rect 263284 126216 263290 126268
rect 249426 125740 249432 125792
rect 249484 125780 249490 125792
rect 266170 125780 266176 125792
rect 249484 125752 266176 125780
rect 249484 125740 249490 125752
rect 266170 125740 266176 125752
rect 266228 125740 266234 125792
rect 168006 125672 168012 125724
rect 168064 125712 168070 125724
rect 213914 125712 213920 125724
rect 168064 125684 213920 125712
rect 168064 125672 168070 125684
rect 213914 125672 213920 125684
rect 213972 125672 213978 125724
rect 254762 125672 254768 125724
rect 254820 125712 254826 125724
rect 265526 125712 265532 125724
rect 254820 125684 265532 125712
rect 254820 125672 254826 125684
rect 265526 125672 265532 125684
rect 265584 125672 265590 125724
rect 167914 125604 167920 125656
rect 167972 125644 167978 125656
rect 214006 125644 214012 125656
rect 167972 125616 214012 125644
rect 167972 125604 167978 125616
rect 214006 125604 214012 125616
rect 214064 125604 214070 125656
rect 263318 125604 263324 125656
rect 263376 125644 263382 125656
rect 266262 125644 266268 125656
rect 263376 125616 266268 125644
rect 263376 125604 263382 125616
rect 266262 125604 266268 125616
rect 266320 125604 266326 125656
rect 231762 125536 231768 125588
rect 231820 125576 231826 125588
rect 264422 125576 264428 125588
rect 231820 125548 264428 125576
rect 231820 125536 231826 125548
rect 264422 125536 264428 125548
rect 264480 125536 264486 125588
rect 230658 124924 230664 124976
rect 230716 124964 230722 124976
rect 259178 124964 259184 124976
rect 230716 124936 259184 124964
rect 230716 124924 230722 124936
rect 259178 124924 259184 124936
rect 259236 124924 259242 124976
rect 230750 124856 230756 124908
rect 230808 124896 230814 124908
rect 264698 124896 264704 124908
rect 230808 124868 264704 124896
rect 230808 124856 230814 124868
rect 264698 124856 264704 124868
rect 264756 124856 264762 124908
rect 282822 124448 282828 124500
rect 282880 124488 282886 124500
rect 287882 124488 287888 124500
rect 282880 124460 287888 124488
rect 282880 124448 282886 124460
rect 287882 124448 287888 124460
rect 287940 124448 287946 124500
rect 259086 124312 259092 124364
rect 259144 124352 259150 124364
rect 266170 124352 266176 124364
rect 259144 124324 266176 124352
rect 259144 124312 259150 124324
rect 266170 124312 266176 124324
rect 266228 124312 266234 124364
rect 173342 124244 173348 124296
rect 173400 124284 173406 124296
rect 214006 124284 214012 124296
rect 173400 124256 214012 124284
rect 173400 124244 173406 124256
rect 214006 124244 214012 124256
rect 214064 124244 214070 124296
rect 261478 124244 261484 124296
rect 261536 124284 261542 124296
rect 265342 124284 265348 124296
rect 261536 124256 265348 124284
rect 261536 124244 261542 124256
rect 265342 124244 265348 124256
rect 265400 124244 265406 124296
rect 166626 124176 166632 124228
rect 166684 124216 166690 124228
rect 213914 124216 213920 124228
rect 166684 124188 213920 124216
rect 166684 124176 166690 124188
rect 213914 124176 213920 124188
rect 213972 124176 213978 124228
rect 247862 124176 247868 124228
rect 247920 124216 247926 124228
rect 265158 124216 265164 124228
rect 247920 124188 265164 124216
rect 247920 124176 247926 124188
rect 265158 124176 265164 124188
rect 265216 124176 265222 124228
rect 231762 124108 231768 124160
rect 231820 124148 231826 124160
rect 239490 124148 239496 124160
rect 231820 124120 239496 124148
rect 231820 124108 231826 124120
rect 239490 124108 239496 124120
rect 239548 124108 239554 124160
rect 231302 123496 231308 123548
rect 231360 123536 231366 123548
rect 250990 123536 250996 123548
rect 231360 123508 250996 123536
rect 231360 123496 231366 123508
rect 250990 123496 250996 123508
rect 251048 123496 251054 123548
rect 282822 123496 282828 123548
rect 282880 123536 282886 123548
rect 288526 123536 288532 123548
rect 282880 123508 288532 123536
rect 282880 123496 282886 123508
rect 288526 123496 288532 123508
rect 288584 123496 288590 123548
rect 231578 123428 231584 123480
rect 231636 123468 231642 123480
rect 257706 123468 257712 123480
rect 231636 123440 257712 123468
rect 231636 123428 231642 123440
rect 257706 123428 257712 123440
rect 257764 123428 257770 123480
rect 257522 123020 257528 123072
rect 257580 123060 257586 123072
rect 264422 123060 264428 123072
rect 257580 123032 264428 123060
rect 257580 123020 257586 123032
rect 264422 123020 264428 123032
rect 264480 123020 264486 123072
rect 256142 122952 256148 123004
rect 256200 122992 256206 123004
rect 265158 122992 265164 123004
rect 256200 122964 265164 122992
rect 256200 122952 256206 122964
rect 265158 122952 265164 122964
rect 265216 122952 265222 123004
rect 171870 122884 171876 122936
rect 171928 122924 171934 122936
rect 213914 122924 213920 122936
rect 171928 122896 213920 122924
rect 171928 122884 171934 122896
rect 213914 122884 213920 122896
rect 213972 122884 213978 122936
rect 242434 122884 242440 122936
rect 242492 122924 242498 122936
rect 266170 122924 266176 122936
rect 242492 122896 266176 122924
rect 242492 122884 242498 122896
rect 266170 122884 266176 122896
rect 266228 122884 266234 122936
rect 170490 122816 170496 122868
rect 170548 122856 170554 122868
rect 214006 122856 214012 122868
rect 170548 122828 214012 122856
rect 170548 122816 170554 122828
rect 214006 122816 214012 122828
rect 214064 122816 214070 122868
rect 240962 122816 240968 122868
rect 241020 122856 241026 122868
rect 265434 122856 265440 122868
rect 241020 122828 265440 122856
rect 241020 122816 241026 122828
rect 265434 122816 265440 122828
rect 265492 122816 265498 122868
rect 231762 122748 231768 122800
rect 231820 122788 231826 122800
rect 262950 122788 262956 122800
rect 231820 122760 262956 122788
rect 231820 122748 231826 122760
rect 262950 122748 262956 122760
rect 263008 122748 263014 122800
rect 231394 122680 231400 122732
rect 231452 122720 231458 122732
rect 260558 122720 260564 122732
rect 231452 122692 260564 122720
rect 231452 122680 231458 122692
rect 260558 122680 260564 122692
rect 260616 122680 260622 122732
rect 231118 122612 231124 122664
rect 231176 122652 231182 122664
rect 260098 122652 260104 122664
rect 231176 122624 260104 122652
rect 231176 122612 231182 122624
rect 260098 122612 260104 122624
rect 260156 122612 260162 122664
rect 231486 122068 231492 122120
rect 231544 122108 231550 122120
rect 256418 122108 256424 122120
rect 231544 122080 256424 122108
rect 231544 122068 231550 122080
rect 256418 122068 256424 122080
rect 256476 122068 256482 122120
rect 253474 121592 253480 121644
rect 253532 121632 253538 121644
rect 264698 121632 264704 121644
rect 253532 121604 264704 121632
rect 253532 121592 253538 121604
rect 264698 121592 264704 121604
rect 264756 121592 264762 121644
rect 181530 121524 181536 121576
rect 181588 121564 181594 121576
rect 213914 121564 213920 121576
rect 181588 121536 213920 121564
rect 181588 121524 181594 121536
rect 213914 121524 213920 121536
rect 213972 121524 213978 121576
rect 176102 121456 176108 121508
rect 176160 121496 176166 121508
rect 214006 121496 214012 121508
rect 176160 121468 214012 121496
rect 176160 121456 176166 121468
rect 214006 121456 214012 121468
rect 214064 121456 214070 121508
rect 260282 121456 260288 121508
rect 260340 121496 260346 121508
rect 265526 121496 265532 121508
rect 260340 121468 265532 121496
rect 260340 121456 260346 121468
rect 265526 121456 265532 121468
rect 265584 121456 265590 121508
rect 231762 121388 231768 121440
rect 231820 121428 231826 121440
rect 264606 121428 264612 121440
rect 231820 121400 264612 121428
rect 231820 121388 231826 121400
rect 264606 121388 264612 121400
rect 264664 121388 264670 121440
rect 231394 121320 231400 121372
rect 231452 121360 231458 121372
rect 250622 121360 250628 121372
rect 231452 121332 250628 121360
rect 231452 121320 231458 121332
rect 250622 121320 250628 121332
rect 250680 121320 250686 121372
rect 231026 120708 231032 120760
rect 231084 120748 231090 120760
rect 261754 120748 261760 120760
rect 231084 120720 261760 120748
rect 231084 120708 231090 120720
rect 261754 120708 261760 120720
rect 261812 120708 261818 120760
rect 258902 120232 258908 120284
rect 258960 120272 258966 120284
rect 265526 120272 265532 120284
rect 258960 120244 265532 120272
rect 258960 120232 258966 120244
rect 265526 120232 265532 120244
rect 265584 120232 265590 120284
rect 174722 120164 174728 120216
rect 174780 120204 174786 120216
rect 213914 120204 213920 120216
rect 174780 120176 213920 120204
rect 174780 120164 174786 120176
rect 213914 120164 213920 120176
rect 213972 120164 213978 120216
rect 250714 120164 250720 120216
rect 250772 120204 250778 120216
rect 266170 120204 266176 120216
rect 250772 120176 266176 120204
rect 250772 120164 250778 120176
rect 266170 120164 266176 120176
rect 266228 120164 266234 120216
rect 166718 120096 166724 120148
rect 166776 120136 166782 120148
rect 214006 120136 214012 120148
rect 166776 120108 214012 120136
rect 166776 120096 166782 120108
rect 214006 120096 214012 120108
rect 214064 120096 214070 120148
rect 249150 120096 249156 120148
rect 249208 120136 249214 120148
rect 265434 120136 265440 120148
rect 249208 120108 265440 120136
rect 249208 120096 249214 120108
rect 265434 120096 265440 120108
rect 265492 120096 265498 120148
rect 231762 120028 231768 120080
rect 231820 120068 231826 120080
rect 242250 120068 242256 120080
rect 231820 120040 242256 120068
rect 231820 120028 231826 120040
rect 242250 120028 242256 120040
rect 242308 120028 242314 120080
rect 230566 119960 230572 120012
rect 230624 120000 230630 120012
rect 235534 120000 235540 120012
rect 230624 119972 235540 120000
rect 230624 119960 230630 119972
rect 235534 119960 235540 119972
rect 235592 119960 235598 120012
rect 231486 119348 231492 119400
rect 231544 119388 231550 119400
rect 253658 119388 253664 119400
rect 231544 119360 253664 119388
rect 231544 119348 231550 119360
rect 253658 119348 253664 119360
rect 253716 119348 253722 119400
rect 170582 118804 170588 118856
rect 170640 118844 170646 118856
rect 213914 118844 213920 118856
rect 170640 118816 213920 118844
rect 170640 118804 170646 118816
rect 213914 118804 213920 118816
rect 213972 118804 213978 118856
rect 252094 118804 252100 118856
rect 252152 118844 252158 118856
rect 266170 118844 266176 118856
rect 252152 118816 266176 118844
rect 252152 118804 252158 118816
rect 266170 118804 266176 118816
rect 266228 118804 266234 118856
rect 180242 118736 180248 118788
rect 180300 118776 180306 118788
rect 214006 118776 214012 118788
rect 180300 118748 214012 118776
rect 180300 118736 180306 118748
rect 214006 118736 214012 118748
rect 214064 118736 214070 118788
rect 241146 118736 241152 118788
rect 241204 118776 241210 118788
rect 265434 118776 265440 118788
rect 241204 118748 265440 118776
rect 241204 118736 241210 118748
rect 265434 118736 265440 118748
rect 265492 118736 265498 118788
rect 238018 118668 238024 118720
rect 238076 118708 238082 118720
rect 265526 118708 265532 118720
rect 238076 118680 265532 118708
rect 238076 118668 238082 118680
rect 265526 118668 265532 118680
rect 265584 118668 265590 118720
rect 282822 118600 282828 118652
rect 282880 118640 282886 118652
rect 290090 118640 290096 118652
rect 282880 118612 290096 118640
rect 282880 118600 282886 118612
rect 290090 118600 290096 118612
rect 290148 118600 290154 118652
rect 282730 118532 282736 118584
rect 282788 118572 282794 118584
rect 286134 118572 286140 118584
rect 282788 118544 286140 118572
rect 282788 118532 282794 118544
rect 286134 118532 286140 118544
rect 286192 118532 286198 118584
rect 230566 118396 230572 118448
rect 230624 118436 230630 118448
rect 235350 118436 235356 118448
rect 230624 118408 235356 118436
rect 230624 118396 230630 118408
rect 235350 118396 235356 118408
rect 235408 118396 235414 118448
rect 231762 118260 231768 118312
rect 231820 118300 231826 118312
rect 235442 118300 235448 118312
rect 231820 118272 235448 118300
rect 231820 118260 231826 118272
rect 235442 118260 235448 118272
rect 235500 118260 235506 118312
rect 231670 117988 231676 118040
rect 231728 118028 231734 118040
rect 254946 118028 254952 118040
rect 231728 118000 254952 118028
rect 231728 117988 231734 118000
rect 254946 117988 254952 118000
rect 255004 117988 255010 118040
rect 265434 117988 265440 118040
rect 265492 118028 265498 118040
rect 265894 118028 265900 118040
rect 265492 118000 265900 118028
rect 265492 117988 265498 118000
rect 265894 117988 265900 118000
rect 265952 117988 265958 118040
rect 235534 117920 235540 117972
rect 235592 117960 235598 117972
rect 266078 117960 266084 117972
rect 235592 117932 266084 117960
rect 235592 117920 235598 117932
rect 266078 117920 266084 117932
rect 266136 117920 266142 117972
rect 265342 117512 265348 117564
rect 265400 117552 265406 117564
rect 265802 117552 265808 117564
rect 265400 117524 265808 117552
rect 265400 117512 265406 117524
rect 265802 117512 265808 117524
rect 265860 117512 265866 117564
rect 254670 117444 254676 117496
rect 254728 117484 254734 117496
rect 265526 117484 265532 117496
rect 254728 117456 265532 117484
rect 254728 117444 254734 117456
rect 265526 117444 265532 117456
rect 265584 117444 265590 117496
rect 244918 117376 244924 117428
rect 244976 117416 244982 117428
rect 265894 117416 265900 117428
rect 244976 117388 265900 117416
rect 244976 117376 244982 117388
rect 265894 117376 265900 117388
rect 265952 117376 265958 117428
rect 178862 117308 178868 117360
rect 178920 117348 178926 117360
rect 213914 117348 213920 117360
rect 178920 117320 213920 117348
rect 178920 117308 178926 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 229738 117308 229744 117360
rect 229796 117348 229802 117360
rect 265802 117348 265808 117360
rect 229796 117320 265808 117348
rect 229796 117308 229802 117320
rect 265802 117308 265808 117320
rect 265860 117308 265866 117360
rect 231762 117240 231768 117292
rect 231820 117280 231826 117292
rect 252278 117280 252284 117292
rect 231820 117252 252284 117280
rect 231820 117240 231826 117252
rect 252278 117240 252284 117252
rect 252336 117240 252342 117292
rect 282822 117240 282828 117292
rect 282880 117280 282886 117292
rect 289078 117280 289084 117292
rect 282880 117252 289084 117280
rect 282880 117240 282886 117252
rect 289078 117240 289084 117252
rect 289136 117240 289142 117292
rect 231118 116628 231124 116680
rect 231176 116668 231182 116680
rect 245194 116668 245200 116680
rect 231176 116640 245200 116668
rect 231176 116628 231182 116640
rect 245194 116628 245200 116640
rect 245252 116628 245258 116680
rect 234246 116560 234252 116612
rect 234304 116600 234310 116612
rect 265434 116600 265440 116612
rect 234304 116572 265440 116600
rect 234304 116560 234310 116572
rect 265434 116560 265440 116572
rect 265492 116560 265498 116612
rect 282822 116424 282828 116476
rect 282880 116464 282886 116476
rect 287790 116464 287796 116476
rect 282880 116436 287796 116464
rect 282880 116424 282886 116436
rect 287790 116424 287796 116436
rect 287848 116424 287854 116476
rect 238294 116152 238300 116204
rect 238352 116192 238358 116204
rect 265894 116192 265900 116204
rect 238352 116164 265900 116192
rect 238352 116152 238358 116164
rect 265894 116152 265900 116164
rect 265952 116152 265958 116204
rect 260098 116084 260104 116136
rect 260156 116124 260162 116136
rect 265802 116124 265808 116136
rect 260156 116096 265808 116124
rect 260156 116084 260162 116096
rect 265802 116084 265808 116096
rect 265860 116084 265866 116136
rect 173434 116016 173440 116068
rect 173492 116056 173498 116068
rect 213914 116056 213920 116068
rect 173492 116028 213920 116056
rect 173492 116016 173498 116028
rect 213914 116016 213920 116028
rect 213972 116016 213978 116068
rect 251818 116016 251824 116068
rect 251876 116056 251882 116068
rect 264606 116056 264612 116068
rect 251876 116028 264612 116056
rect 251876 116016 251882 116028
rect 264606 116016 264612 116028
rect 264664 116016 264670 116068
rect 166810 115948 166816 116000
rect 166868 115988 166874 116000
rect 214006 115988 214012 116000
rect 166868 115960 214012 115988
rect 166868 115948 166874 115960
rect 214006 115948 214012 115960
rect 214064 115948 214070 116000
rect 262950 115948 262956 116000
rect 263008 115988 263014 116000
rect 266078 115988 266084 116000
rect 263008 115960 266084 115988
rect 263008 115948 263014 115960
rect 266078 115948 266084 115960
rect 266136 115948 266142 116000
rect 231762 115880 231768 115932
rect 231820 115920 231826 115932
rect 240870 115920 240876 115932
rect 231820 115892 240876 115920
rect 231820 115880 231826 115892
rect 240870 115880 240876 115892
rect 240928 115880 240934 115932
rect 230934 115812 230940 115864
rect 230992 115852 230998 115864
rect 234062 115852 234068 115864
rect 230992 115824 234068 115852
rect 230992 115812 230998 115824
rect 234062 115812 234068 115824
rect 234120 115812 234126 115864
rect 234154 115200 234160 115252
rect 234212 115240 234218 115252
rect 265342 115240 265348 115252
rect 234212 115212 265348 115240
rect 234212 115200 234218 115212
rect 265342 115200 265348 115212
rect 265400 115200 265406 115252
rect 282822 114792 282828 114844
rect 282880 114832 282886 114844
rect 287330 114832 287336 114844
rect 282880 114804 287336 114832
rect 282880 114792 282886 114804
rect 287330 114792 287336 114804
rect 287388 114792 287394 114844
rect 174814 114588 174820 114640
rect 174872 114628 174878 114640
rect 214006 114628 214012 114640
rect 174872 114600 214012 114628
rect 174872 114588 174878 114600
rect 214006 114588 214012 114600
rect 214064 114588 214070 114640
rect 243722 114588 243728 114640
rect 243780 114628 243786 114640
rect 265802 114628 265808 114640
rect 243780 114600 265808 114628
rect 243780 114588 243786 114600
rect 265802 114588 265808 114600
rect 265860 114588 265866 114640
rect 170766 114520 170772 114572
rect 170824 114560 170830 114572
rect 213914 114560 213920 114572
rect 170824 114532 213920 114560
rect 170824 114520 170830 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 239490 114520 239496 114572
rect 239548 114560 239554 114572
rect 265894 114560 265900 114572
rect 239548 114532 265900 114560
rect 239548 114520 239554 114532
rect 265894 114520 265900 114532
rect 265952 114520 265958 114572
rect 231486 114452 231492 114504
rect 231544 114492 231550 114504
rect 260466 114492 260472 114504
rect 231544 114464 260472 114492
rect 231544 114452 231550 114464
rect 260466 114452 260472 114464
rect 260524 114452 260530 114504
rect 231762 114384 231768 114436
rect 231820 114424 231826 114436
rect 245286 114424 245292 114436
rect 231820 114396 245292 114424
rect 231820 114384 231826 114396
rect 245286 114384 245292 114396
rect 245344 114384 245350 114436
rect 282730 114316 282736 114368
rect 282788 114356 282794 114368
rect 286042 114356 286048 114368
rect 282788 114328 286048 114356
rect 282788 114316 282794 114328
rect 286042 114316 286048 114328
rect 286100 114316 286106 114368
rect 282822 113432 282828 113484
rect 282880 113472 282886 113484
rect 287606 113472 287612 113484
rect 282880 113444 287612 113472
rect 282880 113432 282886 113444
rect 287606 113432 287612 113444
rect 287664 113432 287670 113484
rect 246390 113296 246396 113348
rect 246448 113336 246454 113348
rect 265802 113336 265808 113348
rect 246448 113308 265808 113336
rect 246448 113296 246454 113308
rect 265802 113296 265808 113308
rect 265860 113296 265866 113348
rect 172054 113228 172060 113280
rect 172112 113268 172118 113280
rect 214006 113268 214012 113280
rect 172112 113240 214012 113268
rect 172112 113228 172118 113240
rect 214006 113228 214012 113240
rect 214064 113228 214070 113280
rect 245194 113228 245200 113280
rect 245252 113268 245258 113280
rect 265894 113268 265900 113280
rect 245252 113240 265900 113268
rect 245252 113228 245258 113240
rect 265894 113228 265900 113240
rect 265952 113228 265958 113280
rect 169478 113160 169484 113212
rect 169536 113200 169542 113212
rect 213914 113200 213920 113212
rect 169536 113172 213920 113200
rect 169536 113160 169542 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 235350 113160 235356 113212
rect 235408 113200 235414 113212
rect 265802 113200 265808 113212
rect 235408 113172 265808 113200
rect 235408 113160 235414 113172
rect 265802 113160 265808 113172
rect 265860 113160 265866 113212
rect 231762 113092 231768 113144
rect 231820 113132 231826 113144
rect 249058 113132 249064 113144
rect 231820 113104 249064 113132
rect 231820 113092 231826 113104
rect 249058 113092 249064 113104
rect 249116 113092 249122 113144
rect 231670 113024 231676 113076
rect 231728 113064 231734 113076
rect 242342 113064 242348 113076
rect 231728 113036 242348 113064
rect 231728 113024 231734 113036
rect 242342 113024 242348 113036
rect 242400 113024 242406 113076
rect 282822 112684 282828 112736
rect 282880 112724 282886 112736
rect 286502 112724 286508 112736
rect 282880 112696 286508 112724
rect 282880 112684 282886 112696
rect 286502 112684 286508 112696
rect 286560 112684 286566 112736
rect 168098 112412 168104 112464
rect 168156 112452 168162 112464
rect 215110 112452 215116 112464
rect 168156 112424 215116 112452
rect 168156 112412 168162 112424
rect 215110 112412 215116 112424
rect 215168 112412 215174 112464
rect 231578 112412 231584 112464
rect 231636 112452 231642 112464
rect 251910 112452 251916 112464
rect 231636 112424 251916 112452
rect 231636 112412 231642 112424
rect 251910 112412 251916 112424
rect 251968 112412 251974 112464
rect 252278 111936 252284 111988
rect 252336 111976 252342 111988
rect 265802 111976 265808 111988
rect 252336 111948 265808 111976
rect 252336 111936 252342 111948
rect 265802 111936 265808 111948
rect 265860 111936 265866 111988
rect 171962 111868 171968 111920
rect 172020 111908 172026 111920
rect 213914 111908 213920 111920
rect 172020 111880 213920 111908
rect 172020 111868 172026 111880
rect 213914 111868 213920 111880
rect 213972 111868 213978 111920
rect 250990 111868 250996 111920
rect 251048 111908 251054 111920
rect 265526 111908 265532 111920
rect 251048 111880 265532 111908
rect 251048 111868 251054 111880
rect 265526 111868 265532 111880
rect 265584 111868 265590 111920
rect 170858 111800 170864 111852
rect 170916 111840 170922 111852
rect 214006 111840 214012 111852
rect 170916 111812 214012 111840
rect 170916 111800 170922 111812
rect 214006 111800 214012 111812
rect 214064 111800 214070 111852
rect 242250 111800 242256 111852
rect 242308 111840 242314 111852
rect 265894 111840 265900 111852
rect 242308 111812 265900 111840
rect 242308 111800 242314 111812
rect 265894 111800 265900 111812
rect 265952 111800 265958 111852
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 25498 111772 25504 111784
rect 3476 111744 25504 111772
rect 3476 111732 3482 111744
rect 25498 111732 25504 111744
rect 25556 111732 25562 111784
rect 168282 111732 168288 111784
rect 168340 111772 168346 111784
rect 170674 111772 170680 111784
rect 168340 111744 170680 111772
rect 168340 111732 168346 111744
rect 170674 111732 170680 111744
rect 170732 111732 170738 111784
rect 231486 111732 231492 111784
rect 231544 111772 231550 111784
rect 257338 111772 257344 111784
rect 231544 111744 257344 111772
rect 231544 111732 231550 111744
rect 257338 111732 257344 111744
rect 257396 111732 257402 111784
rect 231762 111664 231768 111716
rect 231820 111704 231826 111716
rect 255958 111704 255964 111716
rect 231820 111676 255964 111704
rect 231820 111664 231826 111676
rect 255958 111664 255964 111676
rect 256016 111664 256022 111716
rect 282822 111120 282828 111172
rect 282880 111160 282886 111172
rect 287698 111160 287704 111172
rect 282880 111132 287704 111160
rect 282880 111120 282886 111132
rect 287698 111120 287704 111132
rect 287756 111120 287762 111172
rect 281994 111052 282000 111104
rect 282052 111092 282058 111104
rect 287238 111092 287244 111104
rect 282052 111064 287244 111092
rect 282052 111052 282058 111064
rect 287238 111052 287244 111064
rect 287296 111052 287302 111104
rect 260466 110576 260472 110628
rect 260524 110616 260530 110628
rect 265158 110616 265164 110628
rect 260524 110588 265164 110616
rect 260524 110576 260530 110588
rect 265158 110576 265164 110588
rect 265216 110576 265222 110628
rect 256418 110508 256424 110560
rect 256476 110548 256482 110560
rect 265802 110548 265808 110560
rect 256476 110520 265808 110548
rect 256476 110508 256482 110520
rect 265802 110508 265808 110520
rect 265860 110508 265866 110560
rect 173526 110440 173532 110492
rect 173584 110480 173590 110492
rect 213914 110480 213920 110492
rect 173584 110452 213920 110480
rect 173584 110440 173590 110452
rect 213914 110440 213920 110452
rect 213972 110440 213978 110492
rect 240870 110440 240876 110492
rect 240928 110480 240934 110492
rect 265894 110480 265900 110492
rect 240928 110452 265900 110480
rect 240928 110440 240934 110452
rect 265894 110440 265900 110452
rect 265952 110440 265958 110492
rect 167546 110372 167552 110424
rect 167604 110412 167610 110424
rect 173158 110412 173164 110424
rect 167604 110384 173164 110412
rect 167604 110372 167610 110384
rect 173158 110372 173164 110384
rect 173216 110372 173222 110424
rect 231762 110372 231768 110424
rect 231820 110412 231826 110424
rect 243630 110412 243636 110424
rect 231820 110384 243636 110412
rect 231820 110372 231826 110384
rect 243630 110372 243636 110384
rect 243688 110372 243694 110424
rect 230934 110168 230940 110220
rect 230992 110208 230998 110220
rect 236730 110208 236736 110220
rect 230992 110180 236736 110208
rect 230992 110168 230998 110180
rect 236730 110168 236736 110180
rect 236788 110168 236794 110220
rect 282822 110032 282828 110084
rect 282880 110072 282886 110084
rect 287054 110072 287060 110084
rect 282880 110044 287060 110072
rect 282880 110032 282886 110044
rect 287054 110032 287060 110044
rect 287112 110032 287118 110084
rect 282270 109896 282276 109948
rect 282328 109936 282334 109948
rect 287146 109936 287152 109948
rect 282328 109908 287152 109936
rect 282328 109896 282334 109908
rect 287146 109896 287152 109908
rect 287204 109896 287210 109948
rect 231762 109420 231768 109472
rect 231820 109460 231826 109472
rect 236822 109460 236828 109472
rect 231820 109432 236828 109460
rect 231820 109420 231826 109432
rect 236822 109420 236828 109432
rect 236880 109420 236886 109472
rect 253382 109148 253388 109200
rect 253440 109188 253446 109200
rect 265802 109188 265808 109200
rect 253440 109160 265808 109188
rect 253440 109148 253446 109160
rect 265802 109148 265808 109160
rect 265860 109148 265866 109200
rect 177482 109080 177488 109132
rect 177540 109120 177546 109132
rect 213914 109120 213920 109132
rect 177540 109092 213920 109120
rect 177540 109080 177546 109092
rect 213914 109080 213920 109092
rect 213972 109080 213978 109132
rect 246298 109080 246304 109132
rect 246356 109120 246362 109132
rect 265894 109120 265900 109132
rect 246356 109092 265900 109120
rect 246356 109080 246362 109092
rect 265894 109080 265900 109092
rect 265952 109080 265958 109132
rect 174906 109012 174912 109064
rect 174964 109052 174970 109064
rect 214006 109052 214012 109064
rect 174964 109024 214012 109052
rect 174964 109012 174970 109024
rect 214006 109012 214012 109024
rect 214064 109012 214070 109064
rect 242342 109012 242348 109064
rect 242400 109052 242406 109064
rect 265342 109052 265348 109064
rect 242400 109024 265348 109052
rect 242400 109012 242406 109024
rect 265342 109012 265348 109024
rect 265400 109012 265406 109064
rect 167546 108944 167552 108996
rect 167604 108984 167610 108996
rect 176010 108984 176016 108996
rect 167604 108956 176016 108984
rect 167604 108944 167610 108956
rect 176010 108944 176016 108956
rect 176068 108944 176074 108996
rect 231762 108944 231768 108996
rect 231820 108984 231826 108996
rect 261662 108984 261668 108996
rect 231820 108956 261668 108984
rect 231820 108944 231826 108956
rect 261662 108944 261668 108956
rect 261720 108944 261726 108996
rect 282362 108944 282368 108996
rect 282420 108984 282426 108996
rect 288986 108984 288992 108996
rect 282420 108956 288992 108984
rect 282420 108944 282426 108956
rect 288986 108944 288992 108956
rect 289044 108944 289050 108996
rect 231670 108876 231676 108928
rect 231728 108916 231734 108928
rect 236638 108916 236644 108928
rect 231728 108888 236644 108916
rect 231728 108876 231734 108888
rect 236638 108876 236644 108888
rect 236696 108876 236702 108928
rect 281534 108604 281540 108656
rect 281592 108644 281598 108656
rect 283374 108644 283380 108656
rect 281592 108616 283380 108644
rect 281592 108604 281598 108616
rect 283374 108604 283380 108616
rect 283432 108604 283438 108656
rect 231026 108536 231032 108588
rect 231084 108576 231090 108588
rect 235258 108576 235264 108588
rect 231084 108548 235264 108576
rect 231084 108536 231090 108548
rect 235258 108536 235264 108548
rect 235316 108536 235322 108588
rect 249058 107856 249064 107908
rect 249116 107896 249122 107908
rect 265802 107896 265808 107908
rect 249116 107868 265808 107896
rect 249116 107856 249122 107868
rect 265802 107856 265808 107868
rect 265860 107856 265866 107908
rect 257706 107788 257712 107840
rect 257764 107828 257770 107840
rect 265526 107828 265532 107840
rect 257764 107800 265532 107828
rect 257764 107788 257770 107800
rect 265526 107788 265532 107800
rect 265584 107788 265590 107840
rect 255958 107720 255964 107772
rect 256016 107760 256022 107772
rect 265802 107760 265808 107772
rect 256016 107732 265808 107760
rect 256016 107720 256022 107732
rect 265802 107720 265808 107732
rect 265860 107720 265866 107772
rect 182910 107652 182916 107704
rect 182968 107692 182974 107704
rect 213914 107692 213920 107704
rect 182968 107664 213920 107692
rect 182968 107652 182974 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 231762 107584 231768 107636
rect 231820 107624 231826 107636
rect 262858 107624 262864 107636
rect 231820 107596 262864 107624
rect 231820 107584 231826 107596
rect 262858 107584 262864 107596
rect 262916 107584 262922 107636
rect 281718 107584 281724 107636
rect 281776 107624 281782 107636
rect 289814 107624 289820 107636
rect 281776 107596 289820 107624
rect 281776 107584 281782 107596
rect 289814 107584 289820 107596
rect 289872 107584 289878 107636
rect 231210 107516 231216 107568
rect 231268 107556 231274 107568
rect 233878 107556 233884 107568
rect 231268 107528 233884 107556
rect 231268 107516 231274 107528
rect 233878 107516 233884 107528
rect 233936 107516 233942 107568
rect 231486 107176 231492 107228
rect 231544 107216 231550 107228
rect 233970 107216 233976 107228
rect 231544 107188 233976 107216
rect 231544 107176 231550 107188
rect 233970 107176 233976 107188
rect 234028 107176 234034 107228
rect 230934 106904 230940 106956
rect 230992 106944 230998 106956
rect 258718 106944 258724 106956
rect 230992 106916 258724 106944
rect 230992 106904 230998 106916
rect 258718 106904 258724 106916
rect 258776 106904 258782 106956
rect 251910 106428 251916 106480
rect 251968 106468 251974 106480
rect 265802 106468 265808 106480
rect 251968 106440 265808 106468
rect 251968 106428 251974 106440
rect 265802 106428 265808 106440
rect 265860 106428 265866 106480
rect 176010 106360 176016 106412
rect 176068 106400 176074 106412
rect 214006 106400 214012 106412
rect 176068 106372 214012 106400
rect 176068 106360 176074 106372
rect 214006 106360 214012 106372
rect 214064 106360 214070 106412
rect 259270 106360 259276 106412
rect 259328 106400 259334 106412
rect 265434 106400 265440 106412
rect 259328 106372 265440 106400
rect 259328 106360 259334 106372
rect 265434 106360 265440 106372
rect 265492 106360 265498 106412
rect 173158 106292 173164 106344
rect 173216 106332 173222 106344
rect 213914 106332 213920 106344
rect 173216 106304 213920 106332
rect 173216 106292 173222 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 263226 106292 263232 106344
rect 263284 106332 263290 106344
rect 265894 106332 265900 106344
rect 263284 106304 265900 106332
rect 263284 106292 263290 106304
rect 265894 106292 265900 106304
rect 265952 106292 265958 106344
rect 231762 106156 231768 106208
rect 231820 106196 231826 106208
rect 241238 106196 241244 106208
rect 231820 106168 241244 106196
rect 231820 106156 231826 106168
rect 241238 106156 241244 106168
rect 241296 106156 241302 106208
rect 231670 106088 231676 106140
rect 231728 106128 231734 106140
rect 254854 106128 254860 106140
rect 231728 106100 254860 106128
rect 231728 106088 231734 106100
rect 254854 106088 254860 106100
rect 254912 106088 254918 106140
rect 230750 106020 230756 106072
rect 230808 106060 230814 106072
rect 232682 106060 232688 106072
rect 230808 106032 232688 106060
rect 230808 106020 230814 106032
rect 232682 106020 232688 106032
rect 232740 106020 232746 106072
rect 230566 105544 230572 105596
rect 230624 105584 230630 105596
rect 256326 105584 256332 105596
rect 230624 105556 256332 105584
rect 230624 105544 230630 105556
rect 256326 105544 256332 105556
rect 256384 105544 256390 105596
rect 282822 105068 282828 105120
rect 282880 105108 282886 105120
rect 288894 105108 288900 105120
rect 282880 105080 288900 105108
rect 282880 105068 282886 105080
rect 288894 105068 288900 105080
rect 288952 105068 288958 105120
rect 170674 105000 170680 105052
rect 170732 105040 170738 105052
rect 213914 105040 213920 105052
rect 170732 105012 213920 105040
rect 170732 105000 170738 105012
rect 213914 105000 213920 105012
rect 213972 105000 213978 105052
rect 250622 105000 250628 105052
rect 250680 105040 250686 105052
rect 265802 105040 265808 105052
rect 250680 105012 265808 105040
rect 250680 105000 250686 105012
rect 265802 105000 265808 105012
rect 265860 105000 265866 105052
rect 168190 104932 168196 104984
rect 168248 104972 168254 104984
rect 214006 104972 214012 104984
rect 168248 104944 214012 104972
rect 168248 104932 168254 104944
rect 214006 104932 214012 104944
rect 214064 104932 214070 104984
rect 166902 104864 166908 104916
rect 166960 104904 166966 104916
rect 214098 104904 214104 104916
rect 166960 104876 214104 104904
rect 166960 104864 166966 104876
rect 214098 104864 214104 104876
rect 214156 104864 214162 104916
rect 260558 104864 260564 104916
rect 260616 104904 260622 104916
rect 265434 104904 265440 104916
rect 260616 104876 265440 104904
rect 260616 104864 260622 104876
rect 265434 104864 265440 104876
rect 265492 104864 265498 104916
rect 231762 104796 231768 104848
rect 231820 104836 231826 104848
rect 250898 104836 250904 104848
rect 231820 104808 250904 104836
rect 231820 104796 231826 104808
rect 250898 104796 250904 104808
rect 250956 104796 250962 104848
rect 281534 104796 281540 104848
rect 281592 104836 281598 104848
rect 283742 104836 283748 104848
rect 281592 104808 283748 104836
rect 281592 104796 281598 104808
rect 283742 104796 283748 104808
rect 283800 104796 283806 104848
rect 230750 104660 230756 104712
rect 230808 104700 230814 104712
rect 232498 104700 232504 104712
rect 230808 104672 232504 104700
rect 230808 104660 230814 104672
rect 232498 104660 232504 104672
rect 232556 104660 232562 104712
rect 281534 104524 281540 104576
rect 281592 104564 281598 104576
rect 283282 104564 283288 104576
rect 281592 104536 283288 104564
rect 281592 104524 281598 104536
rect 283282 104524 283288 104536
rect 283340 104524 283346 104576
rect 230658 104116 230664 104168
rect 230716 104156 230722 104168
rect 263134 104156 263140 104168
rect 230716 104128 263140 104156
rect 230716 104116 230722 104128
rect 263134 104116 263140 104128
rect 263192 104116 263198 104168
rect 258718 103708 258724 103760
rect 258776 103748 258782 103760
rect 265158 103748 265164 103760
rect 258776 103720 265164 103748
rect 258776 103708 258782 103720
rect 265158 103708 265164 103720
rect 265216 103708 265222 103760
rect 263410 103572 263416 103624
rect 263468 103612 263474 103624
rect 265802 103612 265808 103624
rect 263468 103584 265808 103612
rect 263468 103572 263474 103584
rect 265802 103572 265808 103584
rect 265860 103572 265866 103624
rect 168282 103504 168288 103556
rect 168340 103544 168346 103556
rect 213914 103544 213920 103556
rect 168340 103516 213920 103544
rect 168340 103504 168346 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 235258 103504 235264 103556
rect 235316 103544 235322 103556
rect 265342 103544 265348 103556
rect 235316 103516 265348 103544
rect 235316 103504 235322 103516
rect 265342 103504 265348 103516
rect 265400 103504 265406 103556
rect 231486 103436 231492 103488
rect 231544 103476 231550 103488
rect 252186 103476 252192 103488
rect 231544 103448 252192 103476
rect 231544 103436 231550 103448
rect 252186 103436 252192 103448
rect 252244 103436 252250 103488
rect 282822 103436 282828 103488
rect 282880 103476 282886 103488
rect 289998 103476 290004 103488
rect 282880 103448 290004 103476
rect 282880 103436 282886 103448
rect 289998 103436 290004 103448
rect 290056 103436 290062 103488
rect 231762 103368 231768 103420
rect 231820 103408 231826 103420
rect 242618 103408 242624 103420
rect 231820 103380 242624 103408
rect 231820 103368 231826 103380
rect 242618 103368 242624 103380
rect 242676 103368 242682 103420
rect 281994 103232 282000 103284
rect 282052 103272 282058 103284
rect 289262 103272 289268 103284
rect 282052 103244 289268 103272
rect 282052 103232 282058 103244
rect 289262 103232 289268 103244
rect 289320 103232 289326 103284
rect 65702 102416 65708 102468
rect 65760 102456 65766 102468
rect 65978 102456 65984 102468
rect 65760 102428 65984 102456
rect 65760 102416 65766 102428
rect 65978 102416 65984 102428
rect 66036 102416 66042 102468
rect 246574 102348 246580 102400
rect 246632 102388 246638 102400
rect 265434 102388 265440 102400
rect 246632 102360 265440 102388
rect 246632 102348 246638 102360
rect 265434 102348 265440 102360
rect 265492 102348 265498 102400
rect 169754 102212 169760 102264
rect 169812 102252 169818 102264
rect 214006 102252 214012 102264
rect 169812 102224 214012 102252
rect 169812 102212 169818 102224
rect 214006 102212 214012 102224
rect 214064 102212 214070 102264
rect 257338 102212 257344 102264
rect 257396 102252 257402 102264
rect 265802 102252 265808 102264
rect 257396 102224 265808 102252
rect 257396 102212 257402 102224
rect 265802 102212 265808 102224
rect 265860 102212 265866 102264
rect 168374 102144 168380 102196
rect 168432 102184 168438 102196
rect 213914 102184 213920 102196
rect 168432 102156 213920 102184
rect 168432 102144 168438 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 231762 102076 231768 102128
rect 231820 102116 231826 102128
rect 258994 102116 259000 102128
rect 231820 102088 259000 102116
rect 231820 102076 231826 102088
rect 258994 102076 259000 102088
rect 259052 102076 259058 102128
rect 214282 101056 214288 101108
rect 214340 101096 214346 101108
rect 214926 101096 214932 101108
rect 214340 101068 214932 101096
rect 214340 101056 214346 101068
rect 214926 101056 214932 101068
rect 214984 101056 214990 101108
rect 259178 100852 259184 100904
rect 259236 100892 259242 100904
rect 265526 100892 265532 100904
rect 259236 100864 265532 100892
rect 259236 100852 259242 100864
rect 265526 100852 265532 100864
rect 265584 100852 265590 100904
rect 65794 100784 65800 100836
rect 65852 100824 65858 100836
rect 66162 100824 66168 100836
rect 65852 100796 66168 100824
rect 65852 100784 65858 100796
rect 66162 100784 66168 100796
rect 66220 100784 66226 100836
rect 263134 100784 263140 100836
rect 263192 100824 263198 100836
rect 265894 100824 265900 100836
rect 263192 100796 265900 100824
rect 263192 100784 263198 100796
rect 265894 100784 265900 100796
rect 265952 100784 265958 100836
rect 249518 100716 249524 100768
rect 249576 100756 249582 100768
rect 265802 100756 265808 100768
rect 249576 100728 265808 100756
rect 249576 100716 249582 100728
rect 265802 100716 265808 100728
rect 265860 100716 265866 100768
rect 565078 100648 565084 100700
rect 565136 100688 565142 100700
rect 580166 100688 580172 100700
rect 565136 100660 580172 100688
rect 565136 100648 565142 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 231670 100580 231676 100632
rect 231728 100620 231734 100632
rect 234246 100620 234252 100632
rect 231728 100592 234252 100620
rect 231728 100580 231734 100592
rect 234246 100580 234252 100592
rect 234304 100580 234310 100632
rect 282270 100240 282276 100292
rect 282328 100280 282334 100292
rect 285950 100280 285956 100292
rect 282328 100252 285956 100280
rect 282328 100240 282334 100252
rect 285950 100240 285956 100252
rect 286008 100240 286014 100292
rect 230842 100104 230848 100156
rect 230900 100144 230906 100156
rect 235534 100144 235540 100156
rect 230900 100116 235540 100144
rect 230900 100104 230906 100116
rect 235534 100104 235540 100116
rect 235592 100104 235598 100156
rect 231762 99900 231768 99952
rect 231820 99940 231826 99952
rect 238386 99940 238392 99952
rect 231820 99912 238392 99940
rect 231820 99900 231826 99912
rect 238386 99900 238392 99912
rect 238444 99900 238450 99952
rect 230750 99832 230756 99884
rect 230808 99872 230814 99884
rect 232590 99872 232596 99884
rect 230808 99844 232596 99872
rect 230808 99832 230814 99844
rect 232590 99832 232596 99844
rect 232648 99832 232654 99884
rect 254854 99492 254860 99544
rect 254912 99532 254918 99544
rect 265802 99532 265808 99544
rect 254912 99504 265808 99532
rect 254912 99492 254918 99504
rect 265802 99492 265808 99504
rect 265860 99492 265866 99544
rect 238110 99424 238116 99476
rect 238168 99464 238174 99476
rect 265526 99464 265532 99476
rect 238168 99436 265532 99464
rect 238168 99424 238174 99436
rect 265526 99424 265532 99436
rect 265584 99424 265590 99476
rect 233970 99356 233976 99408
rect 234028 99396 234034 99408
rect 265894 99396 265900 99408
rect 234028 99368 265900 99396
rect 234028 99356 234034 99368
rect 265894 99356 265900 99368
rect 265952 99356 265958 99408
rect 231026 99288 231032 99340
rect 231084 99328 231090 99340
rect 249242 99328 249248 99340
rect 231084 99300 249248 99328
rect 231084 99288 231090 99300
rect 249242 99288 249248 99300
rect 249300 99288 249306 99340
rect 166074 98812 166080 98864
rect 166132 98852 166138 98864
rect 166626 98852 166632 98864
rect 166132 98824 166632 98852
rect 166132 98812 166138 98824
rect 166626 98812 166632 98824
rect 166684 98812 166690 98864
rect 166626 98676 166632 98728
rect 166684 98716 166690 98728
rect 166902 98716 166908 98728
rect 166684 98688 166908 98716
rect 166684 98676 166690 98688
rect 166902 98676 166908 98688
rect 166960 98676 166966 98728
rect 233878 98608 233884 98660
rect 233936 98648 233942 98660
rect 266078 98648 266084 98660
rect 233936 98620 266084 98648
rect 233936 98608 233942 98620
rect 266078 98608 266084 98620
rect 266136 98608 266142 98660
rect 262858 98064 262864 98116
rect 262916 98104 262922 98116
rect 265710 98104 265716 98116
rect 262916 98076 265716 98104
rect 262916 98064 262922 98076
rect 265710 98064 265716 98076
rect 265768 98064 265774 98116
rect 169570 97996 169576 98048
rect 169628 98036 169634 98048
rect 213914 98036 213920 98048
rect 169628 98008 213920 98036
rect 169628 97996 169634 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 231118 97996 231124 98048
rect 231176 98036 231182 98048
rect 265802 98036 265808 98048
rect 231176 98008 265808 98036
rect 231176 97996 231182 98008
rect 265802 97996 265808 98008
rect 265860 97996 265866 98048
rect 3418 97588 3424 97640
rect 3476 97628 3482 97640
rect 7558 97628 7564 97640
rect 3476 97600 7564 97628
rect 3476 97588 3482 97600
rect 7558 97588 7564 97600
rect 7616 97588 7622 97640
rect 231578 97588 231584 97640
rect 231636 97628 231642 97640
rect 234154 97628 234160 97640
rect 231636 97600 234160 97628
rect 231636 97588 231642 97600
rect 234154 97588 234160 97600
rect 234212 97588 234218 97640
rect 231762 97316 231768 97368
rect 231820 97356 231826 97368
rect 248414 97356 248420 97368
rect 231820 97328 248420 97356
rect 231820 97316 231826 97328
rect 248414 97316 248420 97328
rect 248472 97356 248478 97368
rect 267550 97356 267556 97368
rect 248472 97328 267556 97356
rect 248472 97316 248478 97328
rect 267550 97316 267556 97328
rect 267608 97316 267614 97368
rect 231302 97248 231308 97300
rect 231360 97288 231366 97300
rect 237282 97288 237288 97300
rect 231360 97260 237288 97288
rect 231360 97248 231366 97260
rect 237282 97248 237288 97260
rect 237340 97288 237346 97300
rect 267274 97288 267280 97300
rect 237340 97260 267280 97288
rect 237340 97248 237346 97260
rect 267274 97248 267280 97260
rect 267332 97248 267338 97300
rect 256326 96772 256332 96824
rect 256384 96812 256390 96824
rect 265526 96812 265532 96824
rect 256384 96784 265532 96812
rect 256384 96772 256390 96784
rect 265526 96772 265532 96784
rect 265584 96772 265590 96824
rect 236638 96704 236644 96756
rect 236696 96744 236702 96756
rect 265618 96744 265624 96756
rect 236696 96716 265624 96744
rect 236696 96704 236702 96716
rect 265618 96704 265624 96716
rect 265676 96704 265682 96756
rect 165522 96636 165528 96688
rect 165580 96676 165586 96688
rect 213914 96676 213920 96688
rect 165580 96648 213920 96676
rect 165580 96636 165586 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 232590 96636 232596 96688
rect 232648 96676 232654 96688
rect 265894 96676 265900 96688
rect 232648 96648 265900 96676
rect 232648 96636 232654 96648
rect 265894 96636 265900 96648
rect 265952 96636 265958 96688
rect 247770 96364 247776 96416
rect 247828 96404 247834 96416
rect 279418 96404 279424 96416
rect 247828 96376 279424 96404
rect 247828 96364 247834 96376
rect 279418 96364 279424 96376
rect 279476 96364 279482 96416
rect 250530 96296 250536 96348
rect 250588 96336 250594 96348
rect 279326 96336 279332 96348
rect 250588 96308 279332 96336
rect 250588 96296 250594 96308
rect 279326 96296 279332 96308
rect 279384 96296 279390 96348
rect 265710 96228 265716 96280
rect 265768 96268 265774 96280
rect 279234 96268 279240 96280
rect 265768 96240 279240 96268
rect 265768 96228 265774 96240
rect 279234 96228 279240 96240
rect 279292 96228 279298 96280
rect 166166 96092 166172 96144
rect 166224 96132 166230 96144
rect 214098 96132 214104 96144
rect 166224 96104 214104 96132
rect 166224 96092 166230 96104
rect 214098 96092 214104 96104
rect 214156 96092 214162 96144
rect 267090 96092 267096 96144
rect 267148 96132 267154 96144
rect 279510 96132 279516 96144
rect 267148 96104 279516 96132
rect 267148 96092 267154 96104
rect 279510 96092 279516 96104
rect 279568 96092 279574 96144
rect 165338 96024 165344 96076
rect 165396 96064 165402 96076
rect 214006 96064 214012 96076
rect 165396 96036 214012 96064
rect 165396 96024 165402 96036
rect 214006 96024 214012 96036
rect 214064 96024 214070 96076
rect 165062 95956 165068 96008
rect 165120 95996 165126 96008
rect 214650 95996 214656 96008
rect 165120 95968 214656 95996
rect 165120 95956 165126 95968
rect 214650 95956 214656 95968
rect 214708 95956 214714 96008
rect 165430 95888 165436 95940
rect 165488 95928 165494 95940
rect 214190 95928 214196 95940
rect 165488 95900 214196 95928
rect 165488 95888 165494 95900
rect 214190 95888 214196 95900
rect 214248 95888 214254 95940
rect 230566 95276 230572 95328
rect 230624 95316 230630 95328
rect 232498 95316 232504 95328
rect 230624 95288 232504 95316
rect 230624 95276 230630 95288
rect 232498 95276 232504 95288
rect 232556 95276 232562 95328
rect 165982 95208 165988 95260
rect 166040 95248 166046 95260
rect 213914 95248 213920 95260
rect 166040 95220 213920 95248
rect 166040 95208 166046 95220
rect 213914 95208 213920 95220
rect 213972 95208 213978 95260
rect 228358 95208 228364 95260
rect 228416 95248 228422 95260
rect 265710 95248 265716 95260
rect 228416 95220 265716 95248
rect 228416 95208 228422 95220
rect 265710 95208 265716 95220
rect 265768 95208 265774 95260
rect 267274 95140 267280 95192
rect 267332 95180 267338 95192
rect 270954 95180 270960 95192
rect 267332 95152 270960 95180
rect 267332 95140 267338 95152
rect 270954 95140 270960 95152
rect 271012 95140 271018 95192
rect 265434 95072 265440 95124
rect 265492 95112 265498 95124
rect 281534 95112 281540 95124
rect 265492 95084 281540 95112
rect 265492 95072 265498 95084
rect 281534 95072 281540 95084
rect 281592 95072 281598 95124
rect 65886 95004 65892 95056
rect 65944 95044 65950 95056
rect 169754 95044 169760 95056
rect 65944 95016 169760 95044
rect 65944 95004 65950 95016
rect 169754 95004 169760 95016
rect 169812 95004 169818 95056
rect 194502 95004 194508 95056
rect 194560 95044 194566 95056
rect 281626 95044 281632 95056
rect 194560 95016 281632 95044
rect 194560 95004 194566 95016
rect 281626 95004 281632 95016
rect 281684 95004 281690 95056
rect 66070 94936 66076 94988
rect 66128 94976 66134 94988
rect 170674 94976 170680 94988
rect 66128 94948 170680 94976
rect 66128 94936 66134 94948
rect 170674 94936 170680 94948
rect 170732 94936 170738 94988
rect 65610 94868 65616 94920
rect 65668 94908 65674 94920
rect 168374 94908 168380 94920
rect 65668 94880 168380 94908
rect 65668 94868 65674 94880
rect 168374 94868 168380 94880
rect 168432 94868 168438 94920
rect 65702 94800 65708 94852
rect 65760 94840 65766 94852
rect 168282 94840 168288 94852
rect 65760 94812 168288 94840
rect 65760 94800 65766 94812
rect 168282 94800 168288 94812
rect 168340 94800 168346 94852
rect 65794 94732 65800 94784
rect 65852 94772 65858 94784
rect 168190 94772 168196 94784
rect 65852 94744 168196 94772
rect 65852 94732 65858 94744
rect 168190 94732 168196 94744
rect 168248 94732 168254 94784
rect 128722 94528 128728 94580
rect 128780 94568 128786 94580
rect 214374 94568 214380 94580
rect 128780 94540 214380 94568
rect 128780 94528 128786 94540
rect 214374 94528 214380 94540
rect 214432 94528 214438 94580
rect 110322 94460 110328 94512
rect 110380 94500 110386 94512
rect 215018 94500 215024 94512
rect 110380 94472 215024 94500
rect 110380 94460 110386 94472
rect 215018 94460 215024 94472
rect 215076 94460 215082 94512
rect 151722 94120 151728 94172
rect 151780 94160 151786 94172
rect 166442 94160 166448 94172
rect 151780 94132 166448 94160
rect 151780 94120 151786 94132
rect 166442 94120 166448 94132
rect 166500 94120 166506 94172
rect 173342 94160 173348 94172
rect 171106 94132 173348 94160
rect 124122 94052 124128 94104
rect 124180 94092 124186 94104
rect 171106 94092 171134 94132
rect 173342 94120 173348 94132
rect 173400 94120 173406 94172
rect 124180 94064 171134 94092
rect 124180 94052 124186 94064
rect 117130 93984 117136 94036
rect 117188 94024 117194 94036
rect 166718 94024 166724 94036
rect 117188 93996 166724 94024
rect 117188 93984 117194 93996
rect 166718 93984 166724 93996
rect 166776 93984 166782 94036
rect 122098 93916 122104 93968
rect 122156 93956 122162 93968
rect 177390 93956 177396 93968
rect 122156 93928 177396 93956
rect 122156 93916 122162 93928
rect 177390 93916 177396 93928
rect 177448 93916 177454 93968
rect 118234 93848 118240 93900
rect 118292 93888 118298 93900
rect 181530 93888 181536 93900
rect 118292 93860 181536 93888
rect 118292 93848 118298 93860
rect 181530 93848 181536 93860
rect 181588 93848 181594 93900
rect 151538 93780 151544 93832
rect 151596 93820 151602 93832
rect 166350 93820 166356 93832
rect 151596 93792 166356 93820
rect 151596 93780 151602 93792
rect 166350 93780 166356 93792
rect 166408 93780 166414 93832
rect 166442 93780 166448 93832
rect 166500 93820 166506 93832
rect 214558 93820 214564 93832
rect 166500 93792 214564 93820
rect 166500 93780 166506 93792
rect 214558 93780 214564 93792
rect 214616 93780 214622 93832
rect 267550 93780 267556 93832
rect 267608 93820 267614 93832
rect 276934 93820 276940 93832
rect 267608 93792 276940 93820
rect 267608 93780 267614 93792
rect 276934 93780 276940 93792
rect 276992 93780 276998 93832
rect 119706 93712 119712 93764
rect 119764 93752 119770 93764
rect 176102 93752 176108 93764
rect 119764 93724 176108 93752
rect 119764 93712 119770 93724
rect 176102 93712 176108 93724
rect 176160 93712 176166 93764
rect 109218 93644 109224 93696
rect 109276 93684 109282 93696
rect 166810 93684 166816 93696
rect 109276 93656 166816 93684
rect 109276 93644 109282 93656
rect 166810 93644 166816 93656
rect 166868 93644 166874 93696
rect 107746 93576 107752 93628
rect 107804 93616 107810 93628
rect 173434 93616 173440 93628
rect 107804 93588 173440 93616
rect 107804 93576 107810 93588
rect 173434 93576 173440 93588
rect 173492 93576 173498 93628
rect 105538 93508 105544 93560
rect 105596 93548 105602 93560
rect 170766 93548 170772 93560
rect 105596 93520 170772 93548
rect 105596 93508 105602 93520
rect 170766 93508 170772 93520
rect 170824 93508 170830 93560
rect 102962 93440 102968 93492
rect 103020 93480 103026 93492
rect 169478 93480 169484 93492
rect 103020 93452 169484 93480
rect 103020 93440 103026 93452
rect 169478 93440 169484 93452
rect 169536 93440 169542 93492
rect 106458 93372 106464 93424
rect 106516 93412 106522 93424
rect 174814 93412 174820 93424
rect 106516 93384 174820 93412
rect 106516 93372 106522 93384
rect 174814 93372 174820 93384
rect 174872 93372 174878 93424
rect 104250 93304 104256 93356
rect 104308 93344 104314 93356
rect 172054 93344 172060 93356
rect 104308 93316 172060 93344
rect 104308 93304 104314 93316
rect 172054 93304 172060 93316
rect 172112 93304 172118 93356
rect 101858 93236 101864 93288
rect 101916 93276 101922 93288
rect 170858 93276 170864 93288
rect 101916 93248 170864 93276
rect 101916 93236 101922 93248
rect 170858 93236 170864 93248
rect 170916 93236 170922 93288
rect 90266 93168 90272 93220
rect 90324 93208 90330 93220
rect 166626 93208 166632 93220
rect 90324 93180 166632 93208
rect 90324 93168 90330 93180
rect 166626 93168 166632 93180
rect 166684 93168 166690 93220
rect 111794 93100 111800 93152
rect 111852 93140 111858 93152
rect 214926 93140 214932 93152
rect 111852 93112 214932 93140
rect 111852 93100 111858 93112
rect 214926 93100 214932 93112
rect 214984 93100 214990 93152
rect 125410 93032 125416 93084
rect 125468 93072 125474 93084
rect 168006 93072 168012 93084
rect 125468 93044 168012 93072
rect 125468 93032 125474 93044
rect 168006 93032 168012 93044
rect 168064 93032 168070 93084
rect 135714 92964 135720 93016
rect 135772 93004 135778 93016
rect 166534 93004 166540 93016
rect 135772 92976 166540 93004
rect 135772 92964 135778 92976
rect 166534 92964 166540 92976
rect 166592 92964 166598 93016
rect 151630 92896 151636 92948
rect 151688 92936 151694 92948
rect 166258 92936 166264 92948
rect 151688 92908 166264 92936
rect 151688 92896 151694 92908
rect 166258 92896 166264 92908
rect 166316 92896 166322 92948
rect 118050 92420 118056 92472
rect 118108 92460 118114 92472
rect 126054 92460 126060 92472
rect 118108 92432 126060 92460
rect 118108 92420 118114 92432
rect 126054 92420 126060 92432
rect 126112 92420 126118 92472
rect 84378 92352 84384 92404
rect 84436 92392 84442 92404
rect 128722 92392 128728 92404
rect 84436 92364 128728 92392
rect 84436 92352 84442 92364
rect 128722 92352 128728 92364
rect 128780 92352 128786 92404
rect 153102 92352 153108 92404
rect 153160 92392 153166 92404
rect 166442 92392 166448 92404
rect 153160 92364 166448 92392
rect 153160 92352 153166 92364
rect 166442 92352 166448 92364
rect 166500 92352 166506 92404
rect 88058 92284 88064 92336
rect 88116 92324 88122 92336
rect 166166 92324 166172 92336
rect 88116 92296 166172 92324
rect 88116 92284 88122 92296
rect 166166 92284 166172 92296
rect 166224 92284 166230 92336
rect 100018 92216 100024 92268
rect 100076 92256 100082 92268
rect 110322 92256 110328 92268
rect 100076 92228 110328 92256
rect 100076 92216 100082 92228
rect 110322 92216 110328 92228
rect 110380 92216 110386 92268
rect 114370 92216 114376 92268
rect 114428 92256 114434 92268
rect 191098 92256 191104 92268
rect 114428 92228 191104 92256
rect 114428 92216 114434 92228
rect 191098 92216 191104 92228
rect 191156 92216 191162 92268
rect 89070 92148 89076 92200
rect 89128 92188 89134 92200
rect 165430 92188 165436 92200
rect 89128 92160 165436 92188
rect 89128 92148 89134 92160
rect 165430 92148 165436 92160
rect 165488 92148 165494 92200
rect 105722 92080 105728 92132
rect 105780 92120 105786 92132
rect 169386 92120 169392 92132
rect 105780 92092 169392 92120
rect 105780 92080 105786 92092
rect 169386 92080 169392 92092
rect 169444 92080 169450 92132
rect 111978 92012 111984 92064
rect 112036 92052 112042 92064
rect 174630 92052 174636 92064
rect 112036 92024 174636 92052
rect 112036 92012 112042 92024
rect 174630 92012 174636 92024
rect 174688 92012 174694 92064
rect 108114 91944 108120 91996
rect 108172 91984 108178 91996
rect 169294 91984 169300 91996
rect 108172 91956 169300 91984
rect 108172 91944 108178 91956
rect 169294 91944 169300 91956
rect 169352 91944 169358 91996
rect 125778 91876 125784 91928
rect 125836 91916 125842 91928
rect 186958 91916 186964 91928
rect 125836 91888 186964 91916
rect 125836 91876 125842 91888
rect 186958 91876 186964 91888
rect 187016 91876 187022 91928
rect 109954 91808 109960 91860
rect 110012 91848 110018 91860
rect 168098 91848 168104 91860
rect 110012 91820 168104 91848
rect 110012 91808 110018 91820
rect 168098 91808 168104 91820
rect 168156 91808 168162 91860
rect 129458 91740 129464 91792
rect 129516 91780 129522 91792
rect 165062 91780 165068 91792
rect 129516 91752 165068 91780
rect 129516 91740 129522 91752
rect 165062 91740 165068 91752
rect 165120 91740 165126 91792
rect 169018 91740 169024 91792
rect 169076 91780 169082 91792
rect 266078 91780 266084 91792
rect 169076 91752 266084 91780
rect 169076 91740 169082 91752
rect 266078 91740 266084 91752
rect 266136 91740 266142 91792
rect 120258 91672 120264 91724
rect 120316 91712 120322 91724
rect 178770 91712 178776 91724
rect 120316 91684 178776 91712
rect 120316 91672 120322 91684
rect 178770 91672 178776 91684
rect 178828 91672 178834 91724
rect 134426 91604 134432 91656
rect 134484 91644 134490 91656
rect 177298 91644 177304 91656
rect 134484 91616 177304 91644
rect 134484 91604 134490 91616
rect 177298 91604 177304 91616
rect 177356 91604 177362 91656
rect 86678 91536 86684 91588
rect 86736 91576 86742 91588
rect 165338 91576 165344 91588
rect 86736 91548 165344 91576
rect 86736 91536 86742 91548
rect 165338 91536 165344 91548
rect 165396 91536 165402 91588
rect 94958 91468 94964 91520
rect 95016 91508 95022 91520
rect 214282 91508 214288 91520
rect 95016 91480 214288 91508
rect 95016 91468 95022 91480
rect 214282 91468 214288 91480
rect 214340 91468 214346 91520
rect 112346 90992 112352 91044
rect 112404 91032 112410 91044
rect 213178 91032 213184 91044
rect 112404 91004 213184 91032
rect 112404 90992 112410 91004
rect 213178 90992 213184 91004
rect 213236 90992 213242 91044
rect 91462 90924 91468 90976
rect 91520 90964 91526 90976
rect 173158 90964 173164 90976
rect 91520 90936 173164 90964
rect 91520 90924 91526 90936
rect 173158 90924 173164 90936
rect 173216 90924 173222 90976
rect 110138 90856 110144 90908
rect 110196 90896 110202 90908
rect 178862 90896 178868 90908
rect 110196 90868 178868 90896
rect 110196 90856 110202 90868
rect 178862 90856 178868 90868
rect 178920 90856 178926 90908
rect 113358 90788 113364 90840
rect 113416 90828 113422 90840
rect 180242 90828 180248 90840
rect 113416 90800 180248 90828
rect 113416 90788 113422 90800
rect 180242 90788 180248 90800
rect 180300 90788 180306 90840
rect 115842 90720 115848 90772
rect 115900 90760 115906 90772
rect 174722 90760 174728 90772
rect 115900 90732 174728 90760
rect 115900 90720 115906 90732
rect 174722 90720 174728 90732
rect 174780 90720 174786 90772
rect 110966 90652 110972 90704
rect 111024 90692 111030 90704
rect 167730 90692 167736 90704
rect 111024 90664 167736 90692
rect 111024 90652 111030 90664
rect 167730 90652 167736 90664
rect 167788 90652 167794 90704
rect 115198 90584 115204 90636
rect 115256 90624 115262 90636
rect 170582 90624 170588 90636
rect 115256 90596 170588 90624
rect 115256 90584 115262 90596
rect 170582 90584 170588 90596
rect 170640 90584 170646 90636
rect 132402 90516 132408 90568
rect 132460 90556 132466 90568
rect 184198 90556 184204 90568
rect 132460 90528 184204 90556
rect 132460 90516 132466 90528
rect 184198 90516 184204 90528
rect 184256 90516 184262 90568
rect 121178 90448 121184 90500
rect 121236 90488 121242 90500
rect 171870 90488 171876 90500
rect 121236 90460 171876 90488
rect 121236 90448 121242 90460
rect 171870 90448 171876 90460
rect 171928 90448 171934 90500
rect 115934 90380 115940 90432
rect 115992 90420 115998 90432
rect 259086 90420 259092 90432
rect 115992 90392 259092 90420
rect 115992 90380 115998 90392
rect 259086 90380 259092 90392
rect 259144 90380 259150 90432
rect 7558 90312 7564 90364
rect 7616 90352 7622 90364
rect 230658 90352 230664 90364
rect 7616 90324 230664 90352
rect 7616 90312 7622 90324
rect 230658 90312 230664 90324
rect 230716 90312 230722 90364
rect 121914 90244 121920 90296
rect 121972 90284 121978 90296
rect 170490 90284 170496 90296
rect 121972 90256 170496 90284
rect 121972 90244 121978 90256
rect 170490 90244 170496 90256
rect 170548 90244 170554 90296
rect 122834 90176 122840 90228
rect 122892 90216 122898 90228
rect 166074 90216 166080 90228
rect 122892 90188 166080 90216
rect 122892 90176 122898 90188
rect 166074 90176 166080 90188
rect 166132 90176 166138 90228
rect 126606 90108 126612 90160
rect 126664 90148 126670 90160
rect 167914 90148 167920 90160
rect 126664 90120 167920 90148
rect 126664 90108 126670 90120
rect 167914 90108 167920 90120
rect 167972 90108 167978 90160
rect 97810 89632 97816 89684
rect 97868 89672 97874 89684
rect 192478 89672 192484 89684
rect 97868 89644 192484 89672
rect 97868 89632 97874 89644
rect 192478 89632 192484 89644
rect 192536 89632 192542 89684
rect 75730 89564 75736 89616
rect 75788 89604 75794 89616
rect 165982 89604 165988 89616
rect 75788 89576 165988 89604
rect 75788 89564 75794 89576
rect 165982 89564 165988 89576
rect 166040 89564 166046 89616
rect 95050 89496 95056 89548
rect 95108 89536 95114 89548
rect 182910 89536 182916 89548
rect 95108 89508 182916 89536
rect 95108 89496 95114 89508
rect 182910 89496 182916 89508
rect 182968 89496 182974 89548
rect 93210 89428 93216 89480
rect 93268 89468 93274 89480
rect 176010 89468 176016 89480
rect 93268 89440 176016 89468
rect 93268 89428 93274 89440
rect 176010 89428 176016 89440
rect 176068 89428 176074 89480
rect 96338 89360 96344 89412
rect 96396 89400 96402 89412
rect 177482 89400 177488 89412
rect 96396 89372 177488 89400
rect 96396 89360 96402 89372
rect 177482 89360 177488 89372
rect 177540 89360 177546 89412
rect 97534 89292 97540 89344
rect 97592 89332 97598 89344
rect 174906 89332 174912 89344
rect 97592 89304 174912 89332
rect 97592 89292 97598 89304
rect 174906 89292 174912 89304
rect 174964 89292 174970 89344
rect 99282 89224 99288 89276
rect 99340 89264 99346 89276
rect 173526 89264 173532 89276
rect 99340 89236 173532 89264
rect 99340 89224 99346 89236
rect 173526 89224 173532 89236
rect 173584 89224 173590 89276
rect 100570 89156 100576 89208
rect 100628 89196 100634 89208
rect 171962 89196 171968 89208
rect 100628 89168 171968 89196
rect 100628 89156 100634 89168
rect 171962 89156 171968 89168
rect 172020 89156 172026 89208
rect 115474 89088 115480 89140
rect 115532 89128 115538 89140
rect 170398 89128 170404 89140
rect 115532 89100 170404 89128
rect 115532 89088 115538 89100
rect 170398 89088 170404 89100
rect 170456 89088 170462 89140
rect 122834 89020 122840 89072
rect 122892 89060 122898 89072
rect 263318 89060 263324 89072
rect 122892 89032 263324 89060
rect 122892 89020 122898 89032
rect 263318 89020 263324 89032
rect 263376 89020 263382 89072
rect 51074 88952 51080 89004
rect 51132 88992 51138 89004
rect 263410 88992 263416 89004
rect 51132 88964 263416 88992
rect 51132 88952 51138 88964
rect 263410 88952 263416 88964
rect 263468 88952 263474 89004
rect 113174 88884 113180 88936
rect 113232 88924 113238 88936
rect 167638 88924 167644 88936
rect 113232 88896 167644 88924
rect 113232 88884 113238 88896
rect 167638 88884 167644 88896
rect 167696 88884 167702 88936
rect 125318 88816 125324 88868
rect 125376 88856 125382 88868
rect 175918 88856 175924 88868
rect 125376 88828 175924 88856
rect 125376 88816 125382 88828
rect 175918 88816 175924 88828
rect 175976 88816 175982 88868
rect 86770 88272 86776 88324
rect 86828 88312 86834 88324
rect 169570 88312 169576 88324
rect 86828 88284 169576 88312
rect 86828 88272 86834 88284
rect 169570 88272 169576 88284
rect 169628 88272 169634 88324
rect 99098 88204 99104 88256
rect 99156 88244 99162 88256
rect 173250 88244 173256 88256
rect 99156 88216 173256 88244
rect 99156 88204 99162 88216
rect 173250 88204 173256 88216
rect 173308 88204 173314 88256
rect 128170 88136 128176 88188
rect 128228 88176 128234 88188
rect 202138 88176 202144 88188
rect 128228 88148 202144 88176
rect 128228 88136 128234 88148
rect 202138 88136 202144 88148
rect 202196 88136 202202 88188
rect 104618 88068 104624 88120
rect 104676 88108 104682 88120
rect 169110 88108 169116 88120
rect 104676 88080 169116 88108
rect 104676 88068 104682 88080
rect 169110 88068 169116 88080
rect 169168 88068 169174 88120
rect 123570 88000 123576 88052
rect 123628 88040 123634 88052
rect 182818 88040 182824 88052
rect 123628 88012 182824 88040
rect 123628 88000 123634 88012
rect 182818 88000 182824 88012
rect 182876 88000 182882 88052
rect 126698 87932 126704 87984
rect 126756 87972 126762 87984
rect 181438 87972 181444 87984
rect 126756 87944 181444 87972
rect 126756 87932 126762 87944
rect 181438 87932 181444 87944
rect 181496 87932 181502 87984
rect 133322 87864 133328 87916
rect 133380 87904 133386 87916
rect 178678 87904 178684 87916
rect 133380 87876 178684 87904
rect 133380 87864 133386 87876
rect 178678 87864 178684 87876
rect 178736 87864 178742 87916
rect 130746 87796 130752 87848
rect 130804 87836 130810 87848
rect 174538 87836 174544 87848
rect 130804 87808 174544 87836
rect 130804 87796 130810 87808
rect 174538 87796 174544 87808
rect 174596 87796 174602 87848
rect 60734 87660 60740 87712
rect 60792 87700 60798 87712
rect 264790 87700 264796 87712
rect 60792 87672 264796 87700
rect 60792 87660 60798 87672
rect 264790 87660 264796 87672
rect 264848 87660 264854 87712
rect 49694 87592 49700 87644
rect 49752 87632 49758 87644
rect 256234 87632 256240 87644
rect 49752 87604 256240 87632
rect 49752 87592 49758 87604
rect 256234 87592 256240 87604
rect 256292 87592 256298 87644
rect 195698 86912 195704 86964
rect 195756 86952 195762 86964
rect 580166 86952 580172 86964
rect 195756 86924 580172 86952
rect 195756 86912 195762 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 63494 86300 63500 86352
rect 63552 86340 63558 86352
rect 257614 86340 257620 86352
rect 63552 86312 257620 86340
rect 63552 86300 63558 86312
rect 257614 86300 257620 86312
rect 257672 86300 257678 86352
rect 64874 86232 64880 86284
rect 64932 86272 64938 86284
rect 260558 86272 260564 86284
rect 64932 86244 260564 86272
rect 64932 86232 64938 86244
rect 260558 86232 260564 86244
rect 260616 86232 260622 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 47578 85524 47584 85536
rect 3200 85496 47584 85524
rect 3200 85484 3206 85496
rect 47578 85484 47584 85496
rect 47636 85484 47642 85536
rect 67634 84872 67640 84924
rect 67692 84912 67698 84924
rect 261570 84912 261576 84924
rect 67692 84884 261576 84912
rect 67692 84872 67698 84884
rect 261570 84872 261576 84884
rect 261628 84872 261634 84924
rect 46934 84804 46940 84856
rect 46992 84844 46998 84856
rect 264698 84844 264704 84856
rect 46992 84816 264704 84844
rect 46992 84804 46998 84816
rect 264698 84804 264704 84816
rect 264756 84804 264762 84856
rect 70394 83512 70400 83564
rect 70452 83552 70458 83564
rect 242526 83552 242532 83564
rect 70452 83524 242532 83552
rect 70452 83512 70458 83524
rect 242526 83512 242532 83524
rect 242584 83512 242590 83564
rect 71774 83444 71780 83496
rect 71832 83484 71838 83496
rect 263226 83484 263232 83496
rect 71832 83456 263232 83484
rect 71832 83444 71838 83456
rect 263226 83444 263232 83456
rect 263284 83444 263290 83496
rect 78674 82152 78680 82204
rect 78732 82192 78738 82204
rect 259270 82192 259276 82204
rect 78732 82164 259276 82192
rect 78732 82152 78738 82164
rect 259270 82152 259276 82164
rect 259328 82152 259334 82204
rect 56594 82084 56600 82136
rect 56652 82124 56658 82136
rect 250806 82124 250812 82136
rect 56652 82096 250812 82124
rect 56652 82084 56658 82096
rect 250806 82084 250812 82096
rect 250864 82084 250870 82136
rect 89714 80724 89720 80776
rect 89772 80764 89778 80776
rect 257706 80764 257712 80776
rect 89772 80736 257712 80764
rect 89772 80724 89778 80736
rect 257706 80724 257712 80736
rect 257764 80724 257770 80776
rect 9674 80656 9680 80708
rect 9732 80696 9738 80708
rect 249426 80696 249432 80708
rect 9732 80668 249432 80696
rect 9732 80656 9738 80668
rect 249426 80656 249432 80668
rect 249484 80656 249490 80708
rect 93854 79364 93860 79416
rect 93912 79404 93918 79416
rect 264606 79404 264612 79416
rect 93912 79376 264612 79404
rect 93912 79364 93918 79376
rect 264606 79364 264612 79376
rect 264664 79364 264670 79416
rect 52454 79296 52460 79348
rect 52512 79336 52518 79348
rect 253566 79336 253572 79348
rect 52512 79308 253572 79336
rect 52512 79296 52518 79308
rect 253566 79296 253572 79308
rect 253624 79296 253630 79348
rect 107654 78004 107660 78056
rect 107712 78044 107718 78056
rect 256418 78044 256424 78056
rect 107712 78016 256424 78044
rect 107712 78004 107718 78016
rect 256418 78004 256424 78016
rect 256476 78004 256482 78056
rect 44174 77936 44180 77988
rect 44232 77976 44238 77988
rect 238294 77976 238300 77988
rect 44232 77948 238300 77976
rect 44232 77936 44238 77948
rect 238294 77936 238300 77948
rect 238352 77936 238358 77988
rect 110414 76576 110420 76628
rect 110472 76616 110478 76628
rect 260466 76616 260472 76628
rect 110472 76588 260472 76616
rect 110472 76576 110478 76588
rect 260466 76576 260472 76588
rect 260524 76576 260530 76628
rect 34514 76508 34520 76560
rect 34572 76548 34578 76560
rect 239490 76548 239496 76560
rect 34572 76520 239496 76548
rect 34572 76508 34578 76520
rect 239490 76508 239496 76520
rect 239548 76508 239554 76560
rect 85574 75216 85580 75268
rect 85632 75256 85638 75268
rect 263042 75256 263048 75268
rect 85632 75228 263048 75256
rect 85632 75216 85638 75228
rect 263042 75216 263048 75228
rect 263100 75216 263106 75268
rect 16574 75148 16580 75200
rect 16632 75188 16638 75200
rect 254854 75188 254860 75200
rect 16632 75160 254860 75188
rect 16632 75148 16638 75160
rect 254854 75148 254860 75160
rect 254912 75148 254918 75200
rect 118694 73856 118700 73908
rect 118752 73896 118758 73908
rect 252278 73896 252284 73908
rect 118752 73868 252284 73896
rect 118752 73856 118758 73868
rect 252278 73856 252284 73868
rect 252336 73856 252342 73908
rect 27614 73788 27620 73840
rect 27672 73828 27678 73840
rect 243722 73828 243728 73840
rect 27672 73800 243728 73828
rect 27672 73788 27678 73800
rect 243722 73788 243728 73800
rect 243780 73788 243786 73840
rect 253290 73108 253296 73160
rect 253348 73148 253354 73160
rect 579982 73148 579988 73160
rect 253348 73120 579988 73148
rect 253348 73108 253354 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 121454 72496 121460 72548
rect 121512 72536 121518 72548
rect 250990 72536 250996 72548
rect 121512 72508 250996 72536
rect 121512 72496 121518 72508
rect 250990 72496 250996 72508
rect 251048 72496 251054 72548
rect 22094 72428 22100 72480
rect 22152 72468 22158 72480
rect 245194 72468 245200 72480
rect 22152 72440 245200 72468
rect 22152 72428 22158 72440
rect 245194 72428 245200 72440
rect 245252 72428 245258 72480
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 195238 71720 195244 71732
rect 3476 71692 195244 71720
rect 3476 71680 3482 71692
rect 195238 71680 195244 71692
rect 195296 71680 195302 71732
rect 118786 71000 118792 71052
rect 118844 71040 118850 71052
rect 254762 71040 254768 71052
rect 118844 71012 254768 71040
rect 118844 71000 118850 71012
rect 254762 71000 254768 71012
rect 254820 71000 254826 71052
rect 88334 69708 88340 69760
rect 88392 69748 88398 69760
rect 260374 69748 260380 69760
rect 88392 69720 260380 69748
rect 88392 69708 88398 69720
rect 260374 69708 260380 69720
rect 260432 69708 260438 69760
rect 26234 69640 26240 69692
rect 26292 69680 26298 69692
rect 249518 69680 249524 69692
rect 26292 69652 249524 69680
rect 26292 69640 26298 69652
rect 249518 69640 249524 69652
rect 249576 69640 249582 69692
rect 106274 68348 106280 68400
rect 106332 68388 106338 68400
rect 229922 68388 229928 68400
rect 106332 68360 229928 68388
rect 106332 68348 106338 68360
rect 229922 68348 229928 68360
rect 229980 68348 229986 68400
rect 28994 68280 29000 68332
rect 29052 68320 29058 68332
rect 259178 68320 259184 68332
rect 29052 68292 259184 68320
rect 29052 68280 29058 68292
rect 259178 68280 259184 68292
rect 259236 68280 259242 68332
rect 110506 66920 110512 66972
rect 110564 66960 110570 66972
rect 252002 66960 252008 66972
rect 110564 66932 252008 66960
rect 110564 66920 110570 66932
rect 252002 66920 252008 66932
rect 252060 66920 252066 66972
rect 33134 66852 33140 66904
rect 33192 66892 33198 66904
rect 263134 66892 263140 66904
rect 33192 66864 263140 66892
rect 33192 66852 33198 66864
rect 263134 66852 263140 66864
rect 263192 66852 263198 66904
rect 120074 65560 120080 65612
rect 120132 65600 120138 65612
rect 243538 65600 243544 65612
rect 120132 65572 243544 65600
rect 120132 65560 120138 65572
rect 243538 65560 243544 65572
rect 243596 65560 243602 65612
rect 40034 65492 40040 65544
rect 40092 65532 40098 65544
rect 261662 65532 261668 65544
rect 40092 65504 261668 65532
rect 40092 65492 40098 65504
rect 261662 65492 261668 65504
rect 261720 65492 261726 65544
rect 124214 64200 124220 64252
rect 124272 64240 124278 64252
rect 246482 64240 246488 64252
rect 124272 64212 246488 64240
rect 124272 64200 124278 64212
rect 246482 64200 246488 64212
rect 246540 64200 246546 64252
rect 2774 64132 2780 64184
rect 2832 64172 2838 64184
rect 256326 64172 256332 64184
rect 2832 64144 256332 64172
rect 2832 64132 2838 64144
rect 256326 64132 256332 64144
rect 256384 64132 256390 64184
rect 99374 62840 99380 62892
rect 99432 62880 99438 62892
rect 249334 62880 249340 62892
rect 99432 62852 249340 62880
rect 99432 62840 99438 62852
rect 249334 62840 249340 62852
rect 249392 62840 249398 62892
rect 62114 62772 62120 62824
rect 62172 62812 62178 62824
rect 241146 62812 241152 62824
rect 62172 62784 241152 62812
rect 62172 62772 62178 62784
rect 241146 62772 241152 62784
rect 241204 62772 241210 62824
rect 69014 61412 69020 61464
rect 69072 61452 69078 61464
rect 252094 61452 252100 61464
rect 69072 61424 252100 61452
rect 69072 61412 69078 61424
rect 252094 61412 252100 61424
rect 252152 61412 252158 61464
rect 42794 61344 42800 61396
rect 42852 61384 42858 61396
rect 241054 61384 241060 61396
rect 42852 61356 241060 61384
rect 42852 61344 42858 61356
rect 241054 61344 241060 61356
rect 241112 61344 241118 61396
rect 209774 60664 209780 60716
rect 209832 60704 209838 60716
rect 580166 60704 580172 60716
rect 209832 60676 580172 60704
rect 209832 60664 209838 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 111794 60052 111800 60104
rect 111852 60092 111858 60104
rect 247862 60092 247868 60104
rect 111852 60064 247868 60092
rect 111852 60052 111858 60064
rect 247862 60052 247868 60064
rect 247920 60052 247926 60104
rect 24854 59984 24860 60036
rect 24912 60024 24918 60036
rect 265894 60024 265900 60036
rect 24912 59996 265900 60024
rect 24912 59984 24918 59996
rect 265894 59984 265900 59996
rect 265952 59984 265958 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 188338 59344 188344 59356
rect 3108 59316 188344 59344
rect 3108 59304 3114 59316
rect 188338 59304 188344 59316
rect 188396 59304 188402 59356
rect 60826 58624 60832 58676
rect 60884 58664 60890 58676
rect 264514 58664 264520 58676
rect 60884 58636 264520 58664
rect 60884 58624 60890 58636
rect 264514 58624 264520 58636
rect 264572 58624 264578 58676
rect 80054 57264 80060 57316
rect 80112 57304 80118 57316
rect 258902 57304 258908 57316
rect 80112 57276 258908 57304
rect 80112 57264 80118 57276
rect 258902 57264 258908 57276
rect 258960 57264 258966 57316
rect 38654 57196 38660 57248
rect 38712 57236 38718 57248
rect 238202 57236 238208 57248
rect 38712 57208 238208 57236
rect 38712 57196 38718 57208
rect 238202 57196 238208 57208
rect 238260 57196 238266 57248
rect 93946 55904 93952 55956
rect 94004 55944 94010 55956
rect 256142 55944 256148 55956
rect 94004 55916 256148 55944
rect 94004 55904 94010 55916
rect 256142 55904 256148 55916
rect 256200 55904 256206 55956
rect 31754 55836 31760 55888
rect 31812 55876 31818 55888
rect 257430 55876 257436 55888
rect 31812 55848 257436 55876
rect 31812 55836 31818 55848
rect 257430 55836 257436 55848
rect 257488 55836 257494 55888
rect 97994 54544 98000 54596
rect 98052 54584 98058 54596
rect 257522 54584 257528 54596
rect 98052 54556 257528 54584
rect 98052 54544 98058 54556
rect 257522 54544 257528 54556
rect 257580 54544 257586 54596
rect 35894 54476 35900 54528
rect 35952 54516 35958 54528
rect 245102 54516 245108 54528
rect 35952 54488 245108 54516
rect 35952 54476 35958 54488
rect 245102 54476 245108 54488
rect 245160 54476 245166 54528
rect 104894 53116 104900 53168
rect 104952 53156 104958 53168
rect 242434 53156 242440 53168
rect 104952 53128 242440 53156
rect 104952 53116 104958 53128
rect 242434 53116 242440 53128
rect 242492 53116 242498 53168
rect 74534 53048 74540 53100
rect 74592 53088 74598 53100
rect 258810 53088 258816 53100
rect 74592 53060 258816 53088
rect 74592 53048 74598 53060
rect 258810 53048 258816 53060
rect 258868 53048 258874 53100
rect 81434 51756 81440 51808
rect 81492 51796 81498 51808
rect 229830 51796 229836 51808
rect 81492 51768 229836 51796
rect 81492 51756 81498 51768
rect 229830 51756 229836 51768
rect 229888 51756 229894 51808
rect 109034 51688 109040 51740
rect 109092 51728 109098 51740
rect 261478 51728 261484 51740
rect 109092 51700 261484 51728
rect 109092 51688 109098 51700
rect 261478 51688 261484 51700
rect 261536 51688 261542 51740
rect 102134 50396 102140 50448
rect 102192 50436 102198 50448
rect 240962 50436 240968 50448
rect 102192 50408 240968 50436
rect 102192 50396 102198 50408
rect 240962 50396 240968 50408
rect 241020 50396 241026 50448
rect 13814 50328 13820 50380
rect 13872 50368 13878 50380
rect 245010 50368 245016 50380
rect 13872 50340 245016 50368
rect 13872 50328 13878 50340
rect 245010 50328 245016 50340
rect 245068 50328 245074 50380
rect 91094 49036 91100 49088
rect 91152 49076 91158 49088
rect 264422 49076 264428 49088
rect 91152 49048 264428 49076
rect 91152 49036 91158 49048
rect 264422 49036 264428 49048
rect 264480 49036 264486 49088
rect 11054 48968 11060 49020
rect 11112 49008 11118 49020
rect 236638 49008 236644 49020
rect 11112 48980 236644 49008
rect 11112 48968 11118 48980
rect 236638 48968 236644 48980
rect 236696 48968 236702 49020
rect 86954 47608 86960 47660
rect 87012 47648 87018 47660
rect 253474 47648 253480 47660
rect 87012 47620 253480 47648
rect 87012 47608 87018 47620
rect 253474 47608 253480 47620
rect 253532 47608 253538 47660
rect 15194 47540 15200 47592
rect 15252 47580 15258 47592
rect 232590 47580 232596 47592
rect 15252 47552 232596 47580
rect 15252 47540 15258 47552
rect 232590 47540 232596 47552
rect 232648 47540 232654 47592
rect 84194 46180 84200 46232
rect 84252 46220 84258 46232
rect 260282 46220 260288 46232
rect 84252 46192 260288 46220
rect 84252 46180 84258 46192
rect 260282 46180 260288 46192
rect 260340 46180 260346 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 209038 45540 209044 45552
rect 3476 45512 209044 45540
rect 3476 45500 3482 45512
rect 209038 45500 209044 45512
rect 209096 45500 209102 45552
rect 92474 44820 92480 44872
rect 92532 44860 92538 44872
rect 256050 44860 256056 44872
rect 92532 44832 256056 44860
rect 92532 44820 92538 44832
rect 256050 44820 256056 44832
rect 256108 44820 256114 44872
rect 12434 43392 12440 43444
rect 12492 43432 12498 43444
rect 235350 43432 235356 43444
rect 12492 43404 235356 43432
rect 12492 43392 12498 43404
rect 235350 43392 235356 43404
rect 235408 43392 235414 43444
rect 77294 42032 77300 42084
rect 77352 42072 77358 42084
rect 250714 42072 250720 42084
rect 77352 42044 250720 42072
rect 77352 42032 77358 42044
rect 250714 42032 250720 42044
rect 250772 42032 250778 42084
rect 44266 40672 44272 40724
rect 44324 40712 44330 40724
rect 246574 40712 246580 40724
rect 44324 40684 246580 40712
rect 44324 40672 44330 40684
rect 246574 40672 246580 40684
rect 246632 40672 246638 40724
rect 96614 39380 96620 39432
rect 96672 39420 96678 39432
rect 242342 39420 242348 39432
rect 96672 39392 242348 39420
rect 96672 39380 96678 39392
rect 242342 39380 242348 39392
rect 242400 39380 242406 39432
rect 45554 39312 45560 39364
rect 45612 39352 45618 39364
rect 264330 39352 264336 39364
rect 45612 39324 264336 39352
rect 45612 39312 45618 39324
rect 264330 39312 264336 39324
rect 264388 39312 264394 39364
rect 73154 37884 73160 37936
rect 73212 37924 73218 37936
rect 249150 37924 249156 37936
rect 73212 37896 249156 37924
rect 73212 37884 73218 37896
rect 249150 37884 249156 37896
rect 249208 37884 249214 37936
rect 66254 36524 66260 36576
rect 66312 36564 66318 36576
rect 238018 36564 238024 36576
rect 66312 36536 238024 36564
rect 66312 36524 66318 36536
rect 238018 36524 238024 36536
rect 238076 36524 238082 36576
rect 59354 35164 59360 35216
rect 59412 35204 59418 35216
rect 254670 35204 254676 35216
rect 59412 35176 254676 35204
rect 59412 35164 59418 35176
rect 254670 35164 254676 35176
rect 254728 35164 254734 35216
rect 20714 33736 20720 33788
rect 20772 33776 20778 33788
rect 233970 33776 233976 33788
rect 20772 33748 233976 33776
rect 20772 33736 20778 33748
rect 233970 33736 233976 33748
rect 234028 33736 234034 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 15838 33096 15844 33108
rect 3568 33068 15844 33096
rect 3568 33056 3574 33068
rect 15838 33056 15844 33068
rect 15896 33056 15902 33108
rect 206278 33056 206284 33108
rect 206336 33096 206342 33108
rect 580166 33096 580172 33108
rect 206336 33068 580172 33096
rect 206336 33056 206342 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 17954 32376 17960 32428
rect 18012 32416 18018 32428
rect 246390 32416 246396 32428
rect 18012 32388 246396 32416
rect 18012 32376 18018 32388
rect 246390 32376 246396 32388
rect 246448 32376 246454 32428
rect 55214 31016 55220 31068
rect 55272 31056 55278 31068
rect 244918 31056 244924 31068
rect 55272 31028 244924 31056
rect 55272 31016 55278 31028
rect 244918 31016 244924 31028
rect 244976 31016 244982 31068
rect 48314 29588 48320 29640
rect 48372 29628 48378 29640
rect 262950 29628 262956 29640
rect 48372 29600 262956 29628
rect 48372 29588 48378 29600
rect 262950 29588 262956 29600
rect 263008 29588 263014 29640
rect 35986 28228 35992 28280
rect 36044 28268 36050 28280
rect 257338 28268 257344 28280
rect 36044 28240 257344 28268
rect 36044 28228 36050 28240
rect 257338 28228 257344 28240
rect 257396 28228 257402 28280
rect 8294 26868 8300 26920
rect 8352 26908 8358 26920
rect 242250 26908 242256 26920
rect 8352 26880 242256 26908
rect 8352 26868 8358 26880
rect 242250 26868 242256 26880
rect 242308 26868 242314 26920
rect 114554 25576 114560 25628
rect 114612 25616 114618 25628
rect 240870 25616 240876 25628
rect 114612 25588 240876 25616
rect 114612 25576 114618 25588
rect 240870 25576 240876 25588
rect 240928 25576 240934 25628
rect 41414 25508 41420 25560
rect 41472 25548 41478 25560
rect 251818 25548 251824 25560
rect 41472 25520 251824 25548
rect 41472 25508 41478 25520
rect 251818 25508 251824 25520
rect 251876 25508 251882 25560
rect 103514 24148 103520 24200
rect 103572 24188 103578 24200
rect 246298 24188 246304 24200
rect 103572 24160 246304 24188
rect 103572 24148 103578 24160
rect 246298 24148 246304 24160
rect 246356 24148 246362 24200
rect 19334 24080 19340 24132
rect 19392 24120 19398 24132
rect 247678 24120 247684 24132
rect 19392 24092 247684 24120
rect 19392 24080 19398 24092
rect 247678 24080 247684 24092
rect 247736 24080 247742 24132
rect 100754 22788 100760 22840
rect 100812 22828 100818 22840
rect 253382 22828 253388 22840
rect 100812 22800 253388 22828
rect 100812 22788 100818 22800
rect 253382 22788 253388 22800
rect 253440 22788 253446 22840
rect 23474 22720 23480 22772
rect 23532 22760 23538 22772
rect 239398 22760 239404 22772
rect 23532 22732 239404 22760
rect 23532 22720 23538 22732
rect 239398 22720 239404 22732
rect 239456 22720 239462 22772
rect 11146 21360 11152 21412
rect 11204 21400 11210 21412
rect 238110 21400 238116 21412
rect 11204 21372 238116 21400
rect 11204 21360 11210 21372
rect 238110 21360 238116 21372
rect 238168 21360 238174 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 196618 20652 196624 20664
rect 3476 20624 196624 20652
rect 3476 20612 3482 20624
rect 196618 20612 196624 20624
rect 196676 20612 196682 20664
rect 260190 20612 260196 20664
rect 260248 20652 260254 20664
rect 579982 20652 579988 20664
rect 260248 20624 579988 20652
rect 260248 20612 260254 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 77386 19932 77392 19984
rect 77444 19972 77450 19984
rect 254578 19972 254584 19984
rect 77444 19944 254584 19972
rect 77444 19932 77450 19944
rect 254578 19932 254584 19944
rect 254636 19932 254642 19984
rect 75914 18572 75920 18624
rect 75972 18612 75978 18624
rect 251910 18612 251916 18624
rect 75972 18584 251916 18612
rect 75972 18572 75978 18584
rect 251910 18572 251916 18584
rect 251968 18572 251974 18624
rect 85666 17280 85672 17332
rect 85724 17320 85730 17332
rect 249058 17320 249064 17332
rect 85724 17292 249064 17320
rect 85724 17280 85730 17292
rect 249058 17280 249064 17292
rect 249116 17280 249122 17332
rect 4154 17212 4160 17264
rect 4212 17252 4218 17264
rect 228358 17252 228364 17264
rect 4212 17224 228364 17252
rect 4212 17212 4218 17224
rect 228358 17212 228364 17224
rect 228416 17212 228422 17264
rect 83274 15920 83280 15972
rect 83332 15960 83338 15972
rect 255958 15960 255964 15972
rect 83332 15932 255964 15960
rect 83332 15920 83338 15932
rect 255958 15920 255964 15932
rect 256016 15920 256022 15972
rect 20162 15852 20168 15904
rect 20220 15892 20226 15904
rect 231118 15892 231124 15904
rect 20220 15864 231124 15892
rect 20220 15852 20226 15864
rect 231118 15852 231124 15864
rect 231176 15852 231182 15904
rect 54938 14424 54944 14476
rect 54996 14464 55002 14476
rect 258718 14464 258724 14476
rect 54996 14436 258724 14464
rect 54996 14424 55002 14436
rect 258718 14424 258724 14436
rect 258776 14424 258782 14476
rect 69106 13064 69112 13116
rect 69164 13104 69170 13116
rect 250622 13104 250628 13116
rect 69164 13076 250628 13104
rect 69164 13064 69170 13076
rect 250622 13064 250628 13076
rect 250680 13064 250686 13116
rect 103330 11772 103336 11824
rect 103388 11812 103394 11824
rect 250438 11812 250444 11824
rect 103388 11784 250444 11812
rect 103388 11772 103394 11784
rect 250438 11772 250444 11784
rect 250496 11772 250502 11824
rect 58434 11704 58440 11756
rect 58492 11744 58498 11756
rect 235258 11744 235264 11756
rect 58492 11716 235264 11744
rect 58492 11704 58498 11716
rect 235258 11704 235264 11716
rect 235316 11704 235322 11756
rect 117314 10344 117320 10396
rect 117372 10384 117378 10396
rect 242158 10384 242164 10396
rect 117372 10356 242164 10384
rect 117372 10344 117378 10356
rect 242158 10344 242164 10356
rect 242216 10344 242222 10396
rect 7466 10276 7472 10328
rect 7524 10316 7530 10328
rect 262858 10316 262864 10328
rect 7524 10288 262864 10316
rect 7524 10276 7530 10288
rect 262858 10276 262864 10288
rect 262916 10276 262922 10328
rect 114002 8984 114008 9036
rect 114060 9024 114066 9036
rect 253198 9024 253204 9036
rect 114060 8996 253204 9024
rect 114060 8984 114066 8996
rect 253198 8984 253204 8996
rect 253256 8984 253262 9036
rect 2866 8916 2872 8968
rect 2924 8956 2930 8968
rect 264238 8956 264244 8968
rect 2924 8928 264244 8956
rect 2924 8916 2930 8928
rect 264238 8916 264244 8928
rect 264296 8916 264302 8968
rect 96246 7624 96252 7676
rect 96304 7664 96310 7676
rect 240778 7664 240784 7676
rect 96304 7636 240784 7664
rect 96304 7624 96310 7636
rect 240778 7624 240784 7636
rect 240836 7624 240842 7676
rect 3970 7556 3976 7608
rect 4028 7596 4034 7608
rect 230750 7596 230756 7608
rect 4028 7568 230756 7596
rect 4028 7556 4034 7568
rect 230750 7556 230756 7568
rect 230808 7556 230814 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 58618 6848 58624 6860
rect 3476 6820 58624 6848
rect 3476 6808 3482 6820
rect 58618 6808 58624 6820
rect 58676 6808 58682 6860
rect 266998 6808 267004 6860
rect 267056 6848 267062 6860
rect 580166 6848 580172 6860
rect 267056 6820 580172 6848
rect 267056 6808 267062 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 38378 6128 38384 6180
rect 38436 6168 38442 6180
rect 260098 6168 260104 6180
rect 38436 6140 260104 6168
rect 38436 6128 38442 6140
rect 260098 6128 260104 6140
rect 260156 6128 260162 6180
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 265802 4808 265808 4820
rect 6512 4780 265808 4808
rect 6512 4768 6518 4780
rect 265802 4768 265808 4780
rect 265860 4768 265866 4820
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 7558 4128 7564 4140
rect 624 4100 7564 4128
rect 624 4088 630 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 125870 3612 125876 3664
rect 125928 3652 125934 3664
rect 180058 3652 180064 3664
rect 125928 3624 180064 3652
rect 125928 3612 125934 3624
rect 180058 3612 180064 3624
rect 180116 3612 180122 3664
rect 28902 3544 28908 3596
rect 28960 3584 28966 3596
rect 169018 3584 169024 3596
rect 28960 3556 169024 3584
rect 28960 3544 28966 3556
rect 169018 3544 169024 3556
rect 169076 3544 169082 3596
rect 44174 3476 44180 3528
rect 44232 3516 44238 3528
rect 45094 3516 45100 3528
rect 44232 3488 45100 3516
rect 44232 3476 44238 3488
rect 45094 3476 45100 3488
rect 45152 3476 45158 3528
rect 52546 3476 52552 3528
rect 52604 3516 52610 3528
rect 229738 3516 229744 3528
rect 52604 3488 229744 3516
rect 52604 3476 52610 3488
rect 229738 3476 229744 3488
rect 229796 3476 229802 3528
rect 232498 3476 232504 3528
rect 232556 3516 232562 3528
rect 235810 3516 235816 3528
rect 232556 3488 235816 3516
rect 232556 3476 232562 3488
rect 235810 3476 235816 3488
rect 235868 3476 235874 3528
rect 31294 3408 31300 3460
rect 31352 3448 31358 3460
rect 233878 3448 233884 3460
rect 31352 3420 233884 3448
rect 31352 3408 31358 3420
rect 233878 3408 233884 3420
rect 233936 3408 233942 3460
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 69014 3340 69020 3392
rect 69072 3380 69078 3392
rect 69934 3380 69940 3392
rect 69072 3352 69940 3380
rect 69072 3340 69078 3352
rect 69934 3340 69940 3352
rect 69992 3340 69998 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 3970 3040 3976 3052
rect 1728 3012 3976 3040
rect 1728 3000 1734 3012
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 251824 700680 251876 700732
rect 267648 700680 267700 700732
rect 195796 700612 195848 700664
rect 300124 700612 300176 700664
rect 198648 700544 198700 700596
rect 332508 700544 332560 700596
rect 235540 700476 235592 700528
rect 413652 700476 413704 700528
rect 197268 700408 197320 700460
rect 397460 700408 397512 700460
rect 234620 700340 234672 700392
rect 478512 700340 478564 700392
rect 529204 700340 529256 700392
rect 559656 700340 559708 700392
rect 40500 700272 40552 700324
rect 50344 700272 50396 700324
rect 195888 700272 195940 700324
rect 218980 700272 219032 700324
rect 247684 700272 247736 700324
rect 543464 700272 543516 700324
rect 154120 700068 154172 700120
rect 155224 700068 155276 700120
rect 105452 699728 105504 699780
rect 108304 699728 108356 699780
rect 24308 699660 24360 699712
rect 26884 699660 26936 699712
rect 347044 699660 347096 699712
rect 348792 699660 348844 699712
rect 422944 699660 422996 699712
rect 429844 699660 429896 699712
rect 526444 699660 526496 699712
rect 527180 699660 527232 699712
rect 212908 696940 212960 696992
rect 580172 696940 580224 696992
rect 253204 696192 253256 696244
rect 283840 696192 283892 696244
rect 3424 683136 3476 683188
rect 246212 683136 246264 683188
rect 295984 683136 296036 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 156604 670692 156656 670744
rect 223028 670692 223080 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 233884 656888 233936 656940
rect 249064 643084 249116 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 28264 632068 28316 632120
rect 260104 630640 260156 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 29644 618264 29696 618316
rect 255964 616836 256016 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 224224 605820 224276 605872
rect 3332 579640 3384 579692
rect 240784 579640 240836 579692
rect 225972 563048 226024 563100
rect 579896 563048 579948 563100
rect 3332 553392 3384 553444
rect 25504 553392 25556 553444
rect 250444 536800 250496 536852
rect 580172 536800 580224 536852
rect 2964 527144 3016 527196
rect 10324 527144 10376 527196
rect 294604 524424 294656 524476
rect 580172 524424 580224 524476
rect 198556 510620 198608 510672
rect 580172 510620 580224 510672
rect 3332 500964 3384 501016
rect 244924 500964 244976 501016
rect 286324 484372 286376 484424
rect 580172 484372 580224 484424
rect 3056 474716 3108 474768
rect 86224 474716 86276 474768
rect 258724 470568 258776 470620
rect 580172 470568 580224 470620
rect 3332 462340 3384 462392
rect 175924 462340 175976 462392
rect 197176 456764 197228 456816
rect 580172 456764 580224 456816
rect 3332 448536 3384 448588
rect 204904 448536 204956 448588
rect 251916 430584 251968 430636
rect 580172 430584 580224 430636
rect 3148 422288 3200 422340
rect 15844 422288 15896 422340
rect 213460 418140 213512 418192
rect 580172 418140 580224 418192
rect 200120 404336 200172 404388
rect 579988 404336 580040 404388
rect 3332 397468 3384 397520
rect 195336 397468 195388 397520
rect 305644 378156 305696 378208
rect 580172 378156 580224 378208
rect 3332 371220 3384 371272
rect 196716 371220 196768 371272
rect 3332 357416 3384 357468
rect 226984 357416 227036 357468
rect 209964 351908 210016 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 232504 345040 232556 345092
rect 250628 324300 250680 324352
rect 579620 324300 579672 324352
rect 3332 318792 3384 318844
rect 214564 318792 214616 318844
rect 234712 312536 234764 312588
rect 246856 312536 246908 312588
rect 316684 311856 316736 311908
rect 580172 311856 580224 311908
rect 3056 298732 3108 298784
rect 244372 298732 244424 298784
rect 250720 298120 250772 298172
rect 580172 298120 580224 298172
rect 88340 297372 88392 297424
rect 232780 297372 232832 297424
rect 218612 295944 218664 295996
rect 347044 295944 347096 295996
rect 71780 294584 71832 294636
rect 240508 294584 240560 294636
rect 201500 293224 201552 293276
rect 244280 293224 244332 293276
rect 3332 292544 3384 292596
rect 11704 292544 11756 292596
rect 15844 291796 15896 291848
rect 209044 291796 209096 291848
rect 214564 291796 214616 291848
rect 241428 291796 241480 291848
rect 233884 289144 233936 289196
rect 245660 289144 245712 289196
rect 198372 289076 198424 289128
rect 422944 289076 422996 289128
rect 224500 288736 224552 288788
rect 251364 288736 251416 288788
rect 222476 288668 222528 288720
rect 250076 288668 250128 288720
rect 216220 288600 216272 288652
rect 247132 288600 247184 288652
rect 220084 288532 220136 288584
rect 251272 288532 251324 288584
rect 214380 288464 214432 288516
rect 249892 288464 249944 288516
rect 235172 288396 235224 288448
rect 287060 288396 287112 288448
rect 204904 288328 204956 288380
rect 208124 288328 208176 288380
rect 224224 288328 224276 288380
rect 225420 288328 225472 288380
rect 226984 288328 227036 288380
rect 228364 288328 228416 288380
rect 201316 287920 201368 287972
rect 287336 287920 287388 287972
rect 202236 287852 202288 287904
rect 289820 287852 289872 287904
rect 220636 287784 220688 287836
rect 247224 287784 247276 287836
rect 86224 287716 86276 287768
rect 246120 287716 246172 287768
rect 26884 287648 26936 287700
rect 218244 287648 218296 287700
rect 232504 287648 232556 287700
rect 243636 287648 243688 287700
rect 231308 287580 231360 287632
rect 251180 287580 251232 287632
rect 217324 287512 217376 287564
rect 248604 287512 248656 287564
rect 216772 287444 216824 287496
rect 248696 287444 248748 287496
rect 239588 287376 239640 287428
rect 291200 287376 291252 287428
rect 232228 287308 232280 287360
rect 292580 287308 292632 287360
rect 222108 287240 222160 287292
rect 287152 287240 287204 287292
rect 211988 287172 212040 287224
rect 287244 287172 287296 287224
rect 230756 287104 230808 287156
rect 249984 287104 250036 287156
rect 229284 287036 229336 287088
rect 249800 287036 249852 287088
rect 209412 286560 209464 286612
rect 280896 286560 280948 286612
rect 219164 286492 219216 286544
rect 248788 286492 248840 286544
rect 208492 286424 208544 286476
rect 283196 286424 283248 286476
rect 156604 286356 156656 286408
rect 202788 286356 202840 286408
rect 207572 286356 207624 286408
rect 283656 286356 283708 286408
rect 155224 286288 155276 286340
rect 204260 286288 204312 286340
rect 215300 286288 215352 286340
rect 248512 286288 248564 286340
rect 210884 286220 210936 286272
rect 247040 286220 247092 286272
rect 195428 286152 195480 286204
rect 207020 286152 207072 286204
rect 236092 286152 236144 286204
rect 278044 286152 278096 286204
rect 195612 286084 195664 286136
rect 203708 286084 203760 286136
rect 205180 286084 205232 286136
rect 247776 286084 247828 286136
rect 3700 286016 3752 286068
rect 206100 286016 206152 286068
rect 237564 286016 237616 286068
rect 285864 286016 285916 286068
rect 197084 285948 197136 286000
rect 217692 285948 217744 286000
rect 228916 285948 228968 286000
rect 280804 285948 280856 286000
rect 194416 285880 194468 285932
rect 204628 285880 204680 285932
rect 211436 285880 211488 285932
rect 265624 285880 265676 285932
rect 196992 285812 197044 285864
rect 203156 285812 203208 285864
rect 234252 285812 234304 285864
rect 244096 285812 244148 285864
rect 196900 285744 196952 285796
rect 210516 285744 210568 285796
rect 227812 285744 227864 285796
rect 243912 285744 243964 285796
rect 195520 285676 195572 285728
rect 205548 285676 205600 285728
rect 226524 285676 226576 285728
rect 250536 285676 250588 285728
rect 196624 285200 196676 285252
rect 242900 285200 242952 285252
rect 229836 285132 229888 285184
rect 250168 285132 250220 285184
rect 201684 285064 201736 285116
rect 249156 285064 249208 285116
rect 214748 284996 214800 285048
rect 256056 284996 256108 285048
rect 231676 284928 231728 284980
rect 284300 284928 284352 284980
rect 223580 284860 223632 284912
rect 247316 284860 247368 284912
rect 225052 284792 225104 284844
rect 251548 284792 251600 284844
rect 212356 284724 212408 284776
rect 244004 284724 244056 284776
rect 192484 284656 192536 284708
rect 223948 284656 224000 284708
rect 238116 284656 238168 284708
rect 283104 284656 283156 284708
rect 195244 284588 195296 284640
rect 230388 284588 230440 284640
rect 241980 284588 242032 284640
rect 288716 284588 288768 284640
rect 236644 284520 236696 284572
rect 252008 284520 252060 284572
rect 239956 284452 240008 284504
rect 289268 284452 289320 284504
rect 188344 284384 188396 284436
rect 227444 284384 227496 284436
rect 233148 284384 233200 284436
rect 249248 284384 249300 284436
rect 18604 284316 18656 284368
rect 213828 284316 213880 284368
rect 240876 284316 240928 284368
rect 298744 284316 298796 284368
rect 242624 284044 242676 284096
rect 283748 284044 283800 284096
rect 238576 283976 238628 284028
rect 251456 283976 251508 284028
rect 237288 283908 237340 283960
rect 244464 283908 244516 283960
rect 243912 283840 243964 283892
rect 282184 283840 282236 283892
rect 244096 283568 244148 283620
rect 282368 283568 282420 283620
rect 245936 282820 245988 282872
rect 305644 282820 305696 282872
rect 58624 281528 58676 281580
rect 197360 281528 197412 281580
rect 245660 280236 245712 280288
rect 287428 280236 287480 280288
rect 193128 280168 193180 280220
rect 197360 280168 197412 280220
rect 245936 280168 245988 280220
rect 289912 280168 289964 280220
rect 193036 278740 193088 278792
rect 197360 278740 197412 278792
rect 245660 278740 245712 278792
rect 454684 278740 454736 278792
rect 194324 276020 194376 276072
rect 197452 276020 197504 276072
rect 29644 275952 29696 276004
rect 197360 275952 197412 276004
rect 246120 275952 246172 276004
rect 526444 275952 526496 276004
rect 245752 275884 245804 275936
rect 258724 275884 258776 275936
rect 245752 273232 245804 273284
rect 285772 273232 285824 273284
rect 169760 273164 169812 273216
rect 197360 273164 197412 273216
rect 245752 271940 245804 271992
rect 288532 271940 288584 271992
rect 194508 271872 194560 271924
rect 197452 271872 197504 271924
rect 258724 271872 258776 271924
rect 580172 271872 580224 271924
rect 15844 269084 15896 269136
rect 197360 269084 197412 269136
rect 245752 269084 245804 269136
rect 288624 269084 288676 269136
rect 3424 269016 3476 269068
rect 197452 269016 197504 269068
rect 6920 268948 6972 269000
rect 197360 268948 197412 269000
rect 245660 267792 245712 267844
rect 291292 267792 291344 267844
rect 245752 267724 245804 267776
rect 291936 267724 291988 267776
rect 28264 267656 28316 267708
rect 197360 267656 197412 267708
rect 245660 266704 245712 266756
rect 245936 266704 245988 266756
rect 3332 266568 3384 266620
rect 7564 266568 7616 266620
rect 245752 266432 245804 266484
rect 284392 266432 284444 266484
rect 192944 266364 192996 266416
rect 197452 266364 197504 266416
rect 245936 266364 245988 266416
rect 565084 266364 565136 266416
rect 246120 266296 246172 266348
rect 316684 266296 316736 266348
rect 192852 265004 192904 265056
rect 197360 265004 197412 265056
rect 17224 264936 17276 264988
rect 197452 264936 197504 264988
rect 25504 264868 25556 264920
rect 197360 264868 197412 264920
rect 196440 263576 196492 263628
rect 197360 263576 197412 263628
rect 10324 262148 10376 262200
rect 197360 262148 197412 262200
rect 245936 259428 245988 259480
rect 286508 259428 286560 259480
rect 244096 259360 244148 259412
rect 580172 259360 580224 259412
rect 245844 259292 245896 259344
rect 245844 259020 245896 259072
rect 195152 258612 195204 258664
rect 197452 258612 197504 258664
rect 246488 258136 246540 258188
rect 288808 258136 288860 258188
rect 26884 258068 26936 258120
rect 197360 258068 197412 258120
rect 245752 258068 245804 258120
rect 292672 258068 292724 258120
rect 246212 256912 246264 256964
rect 246488 256912 246540 256964
rect 246028 256776 246080 256828
rect 246212 256776 246264 256828
rect 194232 256708 194284 256760
rect 197360 256708 197412 256760
rect 246028 256640 246080 256692
rect 286324 256640 286376 256692
rect 245752 255280 245804 255332
rect 267096 255280 267148 255332
rect 195704 253988 195756 254040
rect 197452 253988 197504 254040
rect 47584 253920 47636 253972
rect 197360 253920 197412 253972
rect 3424 253172 3476 253224
rect 191104 253172 191156 253224
rect 194140 252560 194192 252612
rect 197360 252560 197412 252612
rect 246028 252560 246080 252612
rect 280988 252560 281040 252612
rect 246488 252084 246540 252136
rect 246672 252084 246724 252136
rect 246028 251200 246080 251252
rect 291844 251200 291896 251252
rect 136640 251132 136692 251184
rect 197360 251132 197412 251184
rect 246028 249772 246080 249824
rect 284484 249772 284536 249824
rect 196348 248480 196400 248532
rect 197544 248480 197596 248532
rect 245660 248344 245712 248396
rect 251916 248344 251968 248396
rect 246028 248140 246080 248192
rect 250628 248140 250680 248192
rect 196532 247052 196584 247104
rect 198004 247052 198056 247104
rect 3608 246984 3660 247036
rect 197360 246984 197412 247036
rect 246028 246984 246080 247036
rect 255964 246984 256016 247036
rect 246028 245624 246080 245676
rect 280160 245624 280212 245676
rect 248972 244264 249024 244316
rect 579804 244264 579856 244316
rect 11704 244196 11756 244248
rect 197360 244196 197412 244248
rect 245660 244196 245712 244248
rect 295984 244196 296036 244248
rect 195796 244128 195848 244180
rect 197452 244128 197504 244180
rect 246028 242904 246080 242956
rect 292764 242904 292816 242956
rect 249432 242156 249484 242208
rect 580356 242156 580408 242208
rect 195796 241476 195848 241528
rect 198004 241476 198056 241528
rect 246028 241408 246080 241460
rect 294604 241408 294656 241460
rect 245292 240864 245344 240916
rect 462320 240864 462372 240916
rect 243912 240252 243964 240304
rect 3056 240116 3108 240168
rect 201408 240116 201460 240168
rect 242900 240116 242952 240168
rect 243820 240116 243872 240168
rect 580264 240796 580316 240848
rect 244280 240728 244332 240780
rect 580448 240728 580500 240780
rect 7564 240048 7616 240100
rect 212724 240048 212776 240100
rect 238860 240048 238912 240100
rect 529204 240048 529256 240100
rect 175924 239980 175976 240032
rect 232964 239980 233016 240032
rect 235916 239980 235968 240032
rect 201408 239912 201460 239964
rect 225236 239912 225288 239964
rect 249064 239912 249116 239964
rect 216588 239844 216640 239896
rect 243544 239844 243596 239896
rect 243820 239844 243872 239896
rect 244280 239844 244332 239896
rect 245292 239844 245344 239896
rect 248972 239844 249024 239896
rect 196716 239776 196768 239828
rect 221924 239776 221976 239828
rect 227628 239776 227680 239828
rect 251824 239776 251876 239828
rect 233516 239708 233568 239760
rect 243452 239708 243504 239760
rect 243544 239708 243596 239760
rect 250720 239708 250772 239760
rect 221372 239640 221424 239692
rect 364340 239640 364392 239692
rect 232596 239572 232648 239624
rect 494060 239572 494112 239624
rect 198188 239504 198240 239556
rect 231952 239504 232004 239556
rect 243452 239504 243504 239556
rect 250444 239504 250496 239556
rect 199292 239436 199344 239488
rect 281724 239436 281776 239488
rect 3516 239368 3568 239420
rect 233148 239368 233200 239420
rect 239220 239368 239272 239420
rect 245292 239368 245344 239420
rect 228180 239300 228232 239352
rect 247684 239300 247736 239352
rect 50344 238688 50396 238740
rect 219532 238688 219584 238740
rect 240692 238688 240744 238740
rect 243912 238688 243964 238740
rect 108304 238620 108356 238672
rect 214564 238620 214616 238672
rect 239772 238620 239824 238672
rect 253204 238620 253256 238672
rect 202052 238552 202104 238604
rect 243820 238552 243872 238604
rect 204444 238484 204496 238536
rect 243728 238484 243780 238536
rect 191104 238416 191156 238468
rect 231492 238416 231544 238468
rect 236460 238416 236512 238468
rect 249432 238416 249484 238468
rect 195336 238348 195388 238400
rect 209228 238348 209280 238400
rect 215668 238348 215720 238400
rect 229744 238348 229796 238400
rect 233148 238348 233200 238400
rect 242716 238348 242768 238400
rect 195888 238280 195940 238332
rect 208860 238280 208912 238332
rect 215116 238280 215168 238332
rect 234620 238280 234672 238332
rect 218980 238212 219032 238264
rect 290096 238212 290148 238264
rect 213092 238144 213144 238196
rect 290004 238144 290056 238196
rect 207388 238076 207440 238128
rect 290188 238076 290240 238128
rect 200580 238008 200632 238060
rect 287520 238008 287572 238060
rect 234988 237940 235040 237992
rect 260104 237940 260156 237992
rect 240876 237396 240928 237448
rect 244464 237396 244516 237448
rect 216036 237328 216088 237380
rect 258724 237328 258776 237380
rect 197636 237124 197688 237176
rect 229560 237124 229612 237176
rect 230572 237124 230624 237176
rect 231860 237124 231912 237176
rect 209044 236988 209096 237040
rect 229652 236988 229704 237040
rect 199660 236852 199712 236904
rect 230756 236852 230808 236904
rect 199568 236784 199620 236836
rect 231216 236784 231268 236836
rect 212172 236716 212224 236768
rect 267004 236716 267056 236768
rect 25504 236648 25556 236700
rect 230204 236648 230256 236700
rect 238024 236648 238076 236700
rect 245752 236648 245804 236700
rect 240784 236036 240836 236088
rect 245844 236036 245896 236088
rect 204996 235968 205048 236020
rect 206284 235968 206336 236020
rect 239404 235968 239456 236020
rect 243268 235968 243320 236020
rect 238116 235424 238168 235476
rect 245660 235424 245712 235476
rect 236644 235356 236696 235408
rect 246120 235356 246172 235408
rect 199476 235288 199528 235340
rect 230664 235288 230716 235340
rect 197728 235220 197780 235272
rect 281816 235220 281868 235272
rect 237288 234608 237340 234660
rect 238300 234608 238352 234660
rect 199384 233928 199436 233980
rect 230572 233928 230624 233980
rect 7564 233860 7616 233912
rect 210332 233860 210384 233912
rect 235264 233656 235316 233708
rect 237932 233656 237984 233708
rect 291936 233180 291988 233232
rect 579988 233180 580040 233232
rect 180064 229712 180116 229764
rect 245936 229712 245988 229764
rect 256056 219376 256108 219428
rect 580172 219376 580224 219428
rect 3332 215228 3384 215280
rect 17224 215228 17276 215280
rect 249248 206932 249300 206984
rect 579804 206932 579856 206984
rect 3056 202784 3108 202836
rect 238116 202784 238168 202836
rect 235356 199384 235408 199436
rect 580264 199384 580316 199436
rect 208308 197956 208360 198008
rect 286324 197956 286376 198008
rect 249156 193128 249208 193180
rect 580172 193128 580224 193180
rect 214196 191088 214248 191140
rect 286416 191088 286468 191140
rect 3424 188980 3476 189032
rect 192484 188980 192536 189032
rect 206468 188368 206520 188420
rect 229468 188368 229520 188420
rect 229100 188300 229152 188352
rect 284576 188300 284628 188352
rect 204076 187076 204128 187128
rect 233424 187076 233476 187128
rect 222292 187008 222344 187060
rect 285680 187008 285732 187060
rect 205916 186940 205968 186992
rect 284668 186940 284720 186992
rect 218060 184356 218112 184408
rect 233516 184356 233568 184408
rect 237380 184356 237432 184408
rect 286232 184356 286284 184408
rect 224316 184288 224368 184340
rect 282000 184288 282052 184340
rect 226708 184220 226760 184272
rect 285956 184220 286008 184272
rect 211252 184152 211304 184204
rect 284944 184152 284996 184204
rect 213644 182996 213696 183048
rect 229284 182996 229336 183048
rect 203524 182928 203576 182980
rect 281080 182928 281132 182980
rect 201500 182860 201552 182912
rect 290280 182860 290332 182912
rect 194140 182792 194192 182844
rect 289176 182792 289228 182844
rect 211804 181636 211856 181688
rect 232136 181636 232188 181688
rect 236828 181636 236880 181688
rect 284852 181636 284904 181688
rect 226156 181568 226208 181620
rect 283288 181568 283340 181620
rect 218428 181500 218480 181552
rect 280344 181500 280396 181552
rect 217508 181432 217560 181484
rect 285128 181432 285180 181484
rect 199200 180752 199252 180804
rect 230940 180752 230992 180804
rect 196900 180684 196952 180736
rect 233976 180684 234028 180736
rect 196808 180616 196860 180668
rect 233700 180616 233752 180668
rect 194416 180548 194468 180600
rect 232320 180548 232372 180600
rect 195428 180480 195480 180532
rect 229376 180480 229428 180532
rect 195520 180412 195572 180464
rect 234896 180412 234948 180464
rect 193036 180344 193088 180396
rect 233792 180344 233844 180396
rect 246672 180344 246724 180396
rect 279148 180344 279200 180396
rect 228732 180276 228784 180328
rect 285036 180276 285088 180328
rect 221004 180208 221056 180260
rect 286048 180208 286100 180260
rect 205364 180140 205416 180192
rect 284760 180140 284812 180192
rect 200212 180072 200264 180124
rect 282920 180072 282972 180124
rect 201132 180004 201184 180056
rect 229836 180004 229888 180056
rect 223396 179936 223448 179988
rect 232228 179936 232280 179988
rect 222844 179460 222896 179512
rect 229100 179460 229152 179512
rect 252008 179324 252060 179376
rect 579988 179324 580040 179376
rect 223764 178916 223816 178968
rect 232412 178916 232464 178968
rect 220452 178848 220504 178900
rect 229560 178848 229612 178900
rect 199936 178780 199988 178832
rect 230848 178780 230900 178832
rect 241244 178780 241296 178832
rect 280528 178780 280580 178832
rect 200028 178712 200080 178764
rect 231032 178712 231084 178764
rect 243636 178712 243688 178764
rect 283380 178712 283432 178764
rect 202972 178644 203024 178696
rect 283564 178644 283616 178696
rect 114008 178440 114060 178492
rect 169300 178440 169352 178492
rect 114376 178372 114428 178424
rect 170588 178372 170640 178424
rect 110696 178304 110748 178356
rect 169208 178304 169260 178356
rect 112628 178236 112680 178288
rect 173256 178236 173308 178288
rect 148232 178168 148284 178220
rect 213184 178168 213236 178220
rect 97816 178100 97868 178152
rect 170404 178100 170456 178152
rect 110052 178032 110104 178084
rect 192484 178032 192536 178084
rect 196440 177964 196492 178016
rect 234712 177964 234764 178016
rect 196348 177896 196400 177948
rect 234160 177896 234212 177948
rect 196992 177828 197044 177880
rect 235172 177828 235224 177880
rect 246580 177828 246632 177880
rect 283472 177828 283524 177880
rect 195796 177760 195848 177812
rect 234804 177760 234856 177812
rect 240324 177760 240376 177812
rect 283012 177760 283064 177812
rect 195612 177692 195664 177744
rect 235080 177692 235132 177744
rect 244188 177692 244240 177744
rect 287888 177692 287940 177744
rect 196532 177624 196584 177676
rect 233240 177624 233292 177676
rect 234068 177624 234120 177676
rect 288992 177624 289044 177676
rect 199844 177556 199896 177608
rect 134524 177488 134576 177540
rect 165160 177488 165212 177540
rect 224868 177556 224920 177608
rect 229192 177556 229244 177608
rect 232044 177556 232096 177608
rect 287796 177556 287848 177608
rect 230480 177488 230532 177540
rect 233884 177488 233936 177540
rect 286140 177488 286192 177540
rect 133144 177420 133196 177472
rect 165252 177420 165304 177472
rect 219900 177420 219952 177472
rect 281540 177420 281592 177472
rect 103336 177352 103388 177404
rect 129740 177352 129792 177404
rect 130936 177352 130988 177404
rect 165712 177352 165764 177404
rect 202604 177352 202656 177404
rect 281632 177352 281684 177404
rect 127992 177284 128044 177336
rect 165344 177284 165396 177336
rect 192944 177284 192996 177336
rect 287704 177284 287756 177336
rect 129464 177216 129516 177268
rect 165804 177216 165856 177268
rect 206836 177216 206888 177268
rect 233608 177216 233660 177268
rect 124496 177148 124548 177200
rect 166356 177148 166408 177200
rect 217140 177148 217192 177200
rect 234988 177148 235040 177200
rect 122288 177080 122340 177132
rect 169392 177080 169444 177132
rect 227260 177080 227312 177132
rect 233884 177080 233936 177132
rect 120816 177012 120868 177064
rect 170680 177012 170732 177064
rect 118424 176944 118476 176996
rect 174636 176944 174688 176996
rect 107016 176876 107068 176928
rect 167828 176876 167880 176928
rect 108120 176808 108172 176860
rect 174544 176808 174596 176860
rect 116952 176740 117004 176792
rect 191104 176740 191156 176792
rect 115848 176672 115900 176724
rect 202144 176672 202196 176724
rect 125692 176604 125744 176656
rect 166540 176604 166592 176656
rect 193128 176604 193180 176656
rect 278780 176604 278832 176656
rect 135720 176536 135772 176588
rect 213920 176536 213972 176588
rect 123116 176468 123168 176520
rect 166448 176468 166500 176520
rect 197084 176468 197136 176520
rect 227720 176468 227772 176520
rect 119436 176400 119488 176452
rect 167736 176400 167788 176452
rect 104624 176332 104676 176384
rect 167644 176332 167696 176384
rect 98368 176264 98420 176316
rect 166264 176264 166316 176316
rect 100760 176196 100812 176248
rect 170496 176196 170548 176248
rect 99472 176128 99524 176180
rect 169116 176128 169168 176180
rect 105728 176060 105780 176112
rect 175924 176060 175976 176112
rect 246304 176060 246356 176112
rect 280712 176060 280764 176112
rect 129740 175992 129792 176044
rect 214564 175992 214616 176044
rect 230756 175992 230808 176044
rect 231308 175992 231360 176044
rect 246488 175992 246540 176044
rect 280620 175992 280672 176044
rect 102048 175924 102100 175976
rect 173164 175924 173216 175976
rect 194324 175924 194376 175976
rect 288440 175924 288492 175976
rect 128176 175856 128228 175908
rect 165436 175856 165488 175908
rect 280436 175856 280488 175908
rect 281080 175856 281132 175908
rect 132040 175788 132092 175840
rect 165528 175788 165580 175840
rect 278044 175788 278096 175840
rect 282092 175788 282144 175840
rect 158904 175720 158956 175772
rect 166632 175720 166684 175772
rect 165160 175176 165212 175228
rect 213920 175176 213972 175228
rect 165252 175108 165304 175160
rect 214012 175108 214064 175160
rect 231768 175108 231820 175160
rect 242900 175108 242952 175160
rect 230756 175040 230808 175092
rect 244648 175040 244700 175092
rect 165344 174496 165396 174548
rect 214656 174496 214708 174548
rect 249248 174496 249300 174548
rect 265900 174496 265952 174548
rect 229376 174156 229428 174208
rect 229836 174156 229888 174208
rect 258908 174020 258960 174072
rect 265808 174020 265860 174072
rect 256148 173952 256200 174004
rect 265992 173952 266044 174004
rect 241060 173884 241112 173936
rect 264428 173884 264480 173936
rect 165528 173816 165580 173868
rect 213920 173816 213972 173868
rect 231124 173816 231176 173868
rect 251548 173816 251600 173868
rect 165712 173748 165764 173800
rect 214012 173748 214064 173800
rect 231492 173748 231544 173800
rect 244740 173748 244792 173800
rect 263324 172864 263376 172916
rect 266084 172864 266136 172916
rect 253480 172660 253532 172712
rect 265808 172660 265860 172712
rect 252100 172592 252152 172644
rect 265992 172592 266044 172644
rect 250812 172524 250864 172576
rect 265900 172524 265952 172576
rect 165436 172456 165488 172508
rect 214012 172456 214064 172508
rect 231768 172456 231820 172508
rect 244832 172456 244884 172508
rect 165804 172388 165856 172440
rect 213920 172388 213972 172440
rect 231492 172388 231544 172440
rect 245016 172388 245068 172440
rect 231676 172320 231728 172372
rect 239404 172320 239456 172372
rect 231400 171300 231452 171352
rect 231676 171300 231728 171352
rect 256240 171232 256292 171284
rect 265256 171232 265308 171284
rect 251824 171164 251876 171216
rect 265440 171164 265492 171216
rect 250720 171096 250772 171148
rect 265532 171096 265584 171148
rect 166540 171028 166592 171080
rect 213920 171028 213972 171080
rect 231768 171028 231820 171080
rect 248788 171028 248840 171080
rect 231032 170688 231084 170740
rect 231124 170484 231176 170536
rect 231216 170484 231268 170536
rect 233240 170484 233292 170536
rect 167828 170348 167880 170400
rect 214748 170348 214800 170400
rect 229744 170076 229796 170128
rect 230756 170076 230808 170128
rect 253388 169872 253440 169924
rect 265808 169872 265860 169924
rect 249432 169804 249484 169856
rect 265532 169804 265584 169856
rect 235632 169736 235684 169788
rect 265164 169736 265216 169788
rect 166448 169668 166500 169720
rect 214012 169668 214064 169720
rect 231768 169668 231820 169720
rect 247224 169668 247276 169720
rect 166356 169600 166408 169652
rect 213920 169600 213972 169652
rect 259092 168512 259144 168564
rect 265900 168512 265952 168564
rect 257528 168444 257580 168496
rect 265808 168444 265860 168496
rect 238300 168376 238352 168428
rect 265992 168376 266044 168428
rect 169392 168308 169444 168360
rect 213920 168308 213972 168360
rect 231768 168308 231820 168360
rect 248696 168308 248748 168360
rect 170680 168240 170732 168292
rect 214012 168240 214064 168292
rect 231492 168240 231544 168292
rect 247316 168240 247368 168292
rect 231400 168172 231452 168224
rect 244004 168172 244056 168224
rect 280896 167560 280948 167612
rect 282552 167560 282604 167612
rect 242440 167084 242492 167136
rect 265808 167084 265860 167136
rect 238116 167016 238168 167068
rect 265348 167016 265400 167068
rect 167736 166948 167788 167000
rect 213920 166948 213972 167000
rect 291844 166948 291896 167000
rect 580172 166948 580224 167000
rect 174636 166880 174688 166932
rect 214012 166880 214064 166932
rect 191104 166812 191156 166864
rect 214104 166812 214156 166864
rect 231308 166676 231360 166728
rect 235264 166676 235316 166728
rect 231768 166608 231820 166660
rect 234712 166608 234764 166660
rect 240968 166268 241020 166320
rect 265164 166268 265216 166320
rect 231768 165724 231820 165776
rect 234988 165724 235040 165776
rect 249156 165724 249208 165776
rect 265808 165724 265860 165776
rect 254676 165656 254728 165708
rect 265440 165656 265492 165708
rect 170588 165520 170640 165572
rect 214012 165520 214064 165572
rect 231768 165520 231820 165572
rect 240876 165520 240928 165572
rect 202144 165452 202196 165504
rect 213920 165452 213972 165504
rect 231768 164908 231820 164960
rect 234620 164908 234672 164960
rect 231400 164772 231452 164824
rect 233792 164772 233844 164824
rect 263232 164364 263284 164416
rect 265808 164364 265860 164416
rect 254584 164296 254636 164348
rect 265900 164296 265952 164348
rect 249524 164228 249576 164280
rect 265440 164228 265492 164280
rect 3240 164160 3292 164212
rect 18604 164160 18656 164212
rect 169300 164160 169352 164212
rect 213920 164160 213972 164212
rect 231492 164160 231544 164212
rect 244924 164160 244976 164212
rect 173256 164092 173308 164144
rect 214012 164092 214064 164144
rect 231400 163820 231452 163872
rect 233976 163820 234028 163872
rect 231768 163412 231820 163464
rect 235080 163412 235132 163464
rect 239496 163072 239548 163124
rect 265164 163072 265216 163124
rect 260104 162936 260156 162988
rect 265808 162936 265860 162988
rect 169208 162800 169260 162852
rect 213920 162800 213972 162852
rect 280804 162800 280856 162852
rect 281540 162800 281592 162852
rect 192484 162732 192536 162784
rect 214012 162732 214064 162784
rect 260564 161712 260616 161764
rect 265440 161712 265492 161764
rect 256424 161440 256476 161492
rect 265808 161440 265860 161492
rect 174544 161372 174596 161424
rect 213920 161372 213972 161424
rect 231768 161372 231820 161424
rect 248604 161372 248656 161424
rect 282184 161168 282236 161220
rect 285864 161168 285916 161220
rect 231768 160556 231820 160608
rect 234436 160556 234488 160608
rect 257712 160216 257764 160268
rect 265532 160216 265584 160268
rect 250628 160148 250680 160200
rect 265992 160148 266044 160200
rect 241152 160080 241204 160132
rect 242164 160080 242216 160132
rect 242256 160080 242308 160132
rect 265900 160080 265952 160132
rect 167644 160012 167696 160064
rect 214012 160012 214064 160064
rect 175924 159944 175976 159996
rect 213920 159944 213972 159996
rect 231216 159944 231268 159996
rect 240784 159944 240836 159996
rect 231768 159876 231820 159928
rect 244556 159876 244608 159928
rect 230664 159740 230716 159792
rect 232320 159740 232372 159792
rect 264612 159264 264664 159316
rect 266268 159264 266320 159316
rect 282828 159128 282880 159180
rect 287520 159128 287572 159180
rect 235356 158788 235408 158840
rect 265440 158788 265492 158840
rect 235540 158720 235592 158772
rect 265900 158720 265952 158772
rect 173164 158652 173216 158704
rect 213920 158652 213972 158704
rect 231768 158652 231820 158704
rect 251364 158652 251416 158704
rect 231032 158312 231084 158364
rect 233700 158312 233752 158364
rect 238484 158040 238536 158092
rect 266084 158040 266136 158092
rect 235448 157972 235500 158024
rect 265348 157972 265400 158024
rect 282000 157904 282052 157956
rect 284300 157904 284352 157956
rect 281908 157836 281960 157888
rect 288808 157836 288860 157888
rect 259184 157428 259236 157480
rect 265900 157428 265952 157480
rect 253664 157360 253716 157412
rect 265808 157360 265860 157412
rect 169116 157292 169168 157344
rect 214012 157292 214064 157344
rect 231768 157292 231820 157344
rect 250168 157292 250220 157344
rect 282828 157292 282880 157344
rect 292580 157292 292632 157344
rect 170496 157224 170548 157276
rect 213920 157224 213972 157276
rect 231492 157224 231544 157276
rect 244096 157224 244148 157276
rect 252284 156612 252336 156664
rect 265164 156612 265216 156664
rect 282460 156544 282512 156596
rect 285680 156544 285732 156596
rect 254952 156000 255004 156052
rect 265900 156000 265952 156052
rect 240876 155932 240928 155984
rect 265808 155932 265860 155984
rect 166264 155864 166316 155916
rect 213920 155864 213972 155916
rect 230572 155864 230624 155916
rect 250076 155864 250128 155916
rect 282828 155864 282880 155916
rect 291292 155864 291344 155916
rect 170404 155796 170456 155848
rect 214012 155796 214064 155848
rect 230480 155796 230532 155848
rect 232228 155796 232280 155848
rect 282184 155728 282236 155780
rect 283196 155728 283248 155780
rect 230480 155252 230532 155304
rect 232136 155252 232188 155304
rect 260472 154708 260524 154760
rect 265808 154708 265860 154760
rect 261760 154640 261812 154692
rect 265532 154640 265584 154692
rect 250996 154572 251048 154624
rect 265440 154572 265492 154624
rect 282092 154096 282144 154148
rect 286416 154096 286468 154148
rect 230756 153824 230808 153876
rect 230756 153620 230808 153672
rect 255964 153348 256016 153400
rect 265808 153348 265860 153400
rect 166448 153280 166500 153332
rect 214012 153280 214064 153332
rect 249064 153280 249116 153332
rect 265532 153280 265584 153332
rect 282276 153280 282328 153332
rect 286324 153280 286376 153332
rect 166264 153212 166316 153264
rect 213920 153212 213972 153264
rect 242348 153212 242400 153264
rect 264520 153212 264572 153264
rect 231768 153144 231820 153196
rect 251456 153144 251508 153196
rect 282092 153144 282144 153196
rect 292764 153144 292816 153196
rect 231124 153076 231176 153128
rect 234896 153076 234948 153128
rect 231308 153008 231360 153060
rect 236644 153008 236696 153060
rect 251916 151852 251968 151904
rect 265256 151852 265308 151904
rect 166356 151784 166408 151836
rect 213920 151784 213972 151836
rect 243636 151784 243688 151836
rect 265808 151784 265860 151836
rect 282276 151716 282328 151768
rect 285036 151716 285088 151768
rect 176016 151036 176068 151088
rect 214840 151036 214892 151088
rect 257344 151036 257396 151088
rect 265900 151036 265952 151088
rect 281632 150968 281684 151020
rect 283564 150968 283616 151020
rect 236736 150560 236788 150612
rect 265808 150560 265860 150612
rect 236828 150492 236880 150544
rect 265348 150492 265400 150544
rect 173164 150424 173216 150476
rect 214012 150424 214064 150476
rect 236644 150424 236696 150476
rect 265072 150424 265124 150476
rect 169024 150356 169076 150408
rect 213920 150356 213972 150408
rect 231768 150356 231820 150408
rect 247132 150356 247184 150408
rect 230756 150288 230808 150340
rect 233516 150288 233568 150340
rect 261668 149200 261720 149252
rect 265348 149200 265400 149252
rect 282828 149200 282880 149252
rect 288440 149200 288492 149252
rect 262864 149132 262916 149184
rect 265808 149132 265860 149184
rect 235264 149064 235316 149116
rect 265532 149064 265584 149116
rect 166632 148996 166684 149048
rect 213920 148996 213972 149048
rect 231768 148996 231820 149048
rect 249984 148996 250036 149048
rect 282828 148996 282880 149048
rect 292672 148996 292724 149048
rect 282092 148860 282144 148912
rect 284944 148860 284996 148912
rect 231216 148724 231268 148776
rect 233424 148724 233476 148776
rect 233976 147704 234028 147756
rect 266084 147704 266136 147756
rect 166540 147636 166592 147688
rect 213920 147636 213972 147688
rect 233884 147636 233936 147688
rect 265900 147636 265952 147688
rect 231768 147568 231820 147620
rect 251272 147568 251324 147620
rect 230572 147092 230624 147144
rect 232412 147092 232464 147144
rect 245292 146888 245344 146940
rect 265808 146888 265860 146940
rect 258724 146412 258776 146464
rect 265808 146412 265860 146464
rect 178684 146344 178736 146396
rect 213920 146344 213972 146396
rect 254860 146344 254912 146396
rect 265532 146344 265584 146396
rect 177304 146276 177356 146328
rect 214012 146276 214064 146328
rect 232504 146276 232556 146328
rect 265900 146276 265952 146328
rect 231308 146208 231360 146260
rect 234804 146208 234856 146260
rect 231676 145596 231728 145648
rect 241796 145596 241848 145648
rect 232688 145528 232740 145580
rect 265256 145528 265308 145580
rect 256332 145052 256384 145104
rect 265808 145052 265860 145104
rect 282828 145052 282880 145104
rect 288716 145052 288768 145104
rect 184204 144984 184256 145036
rect 214012 144984 214064 145036
rect 231124 144984 231176 145036
rect 233608 144984 233660 145036
rect 250904 144984 250956 145036
rect 265900 144984 265952 145036
rect 174544 144916 174596 144968
rect 213920 144916 213972 144968
rect 242624 144916 242676 144968
rect 265164 144916 265216 144968
rect 231308 144848 231360 144900
rect 245108 144848 245160 144900
rect 231768 144780 231820 144832
rect 241152 144780 241204 144832
rect 281908 144440 281960 144492
rect 284392 144440 284444 144492
rect 241244 144168 241296 144220
rect 265256 144168 265308 144220
rect 263140 143624 263192 143676
rect 265808 143624 265860 143676
rect 202144 143556 202196 143608
rect 213920 143556 213972 143608
rect 252192 143556 252244 143608
rect 265348 143556 265400 143608
rect 231308 143488 231360 143540
rect 245200 143488 245252 143540
rect 282828 143488 282880 143540
rect 289912 143488 289964 143540
rect 231768 143420 231820 143472
rect 238024 143420 238076 143472
rect 186964 142196 187016 142248
rect 213920 142196 213972 142248
rect 181444 142128 181496 142180
rect 214012 142128 214064 142180
rect 245200 142128 245252 142180
rect 265164 142128 265216 142180
rect 231768 142060 231820 142112
rect 248512 142060 248564 142112
rect 231400 141992 231452 142044
rect 244372 141992 244424 142044
rect 231768 141652 231820 141704
rect 235172 141652 235224 141704
rect 182824 140836 182876 140888
rect 213920 140836 213972 140888
rect 244280 140836 244332 140888
rect 265808 140836 265860 140888
rect 175924 140768 175976 140820
rect 214012 140768 214064 140820
rect 232596 140768 232648 140820
rect 265900 140768 265952 140820
rect 231768 140700 231820 140752
rect 251180 140700 251232 140752
rect 231216 140632 231268 140684
rect 249892 140632 249944 140684
rect 244280 140088 244332 140140
rect 231216 140020 231268 140072
rect 234068 140020 234120 140072
rect 266268 140020 266320 140072
rect 282828 139816 282880 139868
rect 287428 139816 287480 139868
rect 259000 139544 259052 139596
rect 265532 139544 265584 139596
rect 178776 139476 178828 139528
rect 213920 139476 213972 139528
rect 246488 139476 246540 139528
rect 265900 139476 265952 139528
rect 177396 139408 177448 139460
rect 214012 139408 214064 139460
rect 243544 139408 243596 139460
rect 265808 139408 265860 139460
rect 266176 139408 266228 139460
rect 282828 139340 282880 139392
rect 289176 139340 289228 139392
rect 298744 139340 298796 139392
rect 580172 139340 580224 139392
rect 265900 139204 265952 139256
rect 231308 138796 231360 138848
rect 234160 138796 234212 138848
rect 231124 138728 231176 138780
rect 254584 138728 254636 138780
rect 238392 138660 238444 138712
rect 261576 138660 261628 138712
rect 253204 138116 253256 138168
rect 265440 138116 265492 138168
rect 252008 138048 252060 138100
rect 265532 138048 265584 138100
rect 242164 137980 242216 138032
rect 265992 137980 266044 138032
rect 3240 137912 3292 137964
rect 26884 137912 26936 137964
rect 231676 137912 231728 137964
rect 249800 137912 249852 137964
rect 282276 137912 282328 137964
rect 290188 137912 290240 137964
rect 231768 137844 231820 137896
rect 247040 137844 247092 137896
rect 281632 137844 281684 137896
rect 283472 137844 283524 137896
rect 170680 137232 170732 137284
rect 214748 137232 214800 137284
rect 231308 137232 231360 137284
rect 249524 137232 249576 137284
rect 250444 136756 250496 136808
rect 265532 136756 265584 136808
rect 249340 136688 249392 136740
rect 265992 136688 266044 136740
rect 170404 136620 170456 136672
rect 213920 136620 213972 136672
rect 229928 136620 229980 136672
rect 265440 136620 265492 136672
rect 231400 136552 231452 136604
rect 263324 136552 263376 136604
rect 280988 136552 281040 136604
rect 281632 136552 281684 136604
rect 282828 136552 282880 136604
rect 290280 136552 290332 136604
rect 231768 136484 231820 136536
rect 256148 136484 256200 136536
rect 240784 135464 240836 135516
rect 265256 135464 265308 135516
rect 191104 135396 191156 135448
rect 214012 135396 214064 135448
rect 260380 135396 260432 135448
rect 264520 135396 264572 135448
rect 174636 135328 174688 135380
rect 213920 135328 213972 135380
rect 256056 135328 256108 135380
rect 262588 135328 262640 135380
rect 167644 135260 167696 135312
rect 214104 135260 214156 135312
rect 263048 135260 263100 135312
rect 265992 135260 266044 135312
rect 231676 135192 231728 135244
rect 258908 135192 258960 135244
rect 231584 135124 231636 135176
rect 252100 135124 252152 135176
rect 281816 135124 281868 135176
rect 283656 135124 283708 135176
rect 231768 135056 231820 135108
rect 241060 135056 241112 135108
rect 258816 134036 258868 134088
rect 265992 134036 266044 134088
rect 254584 133968 254636 134020
rect 264520 133968 264572 134020
rect 167736 133900 167788 133952
rect 213920 133900 213972 133952
rect 214472 133900 214524 133952
rect 214656 133900 214708 133952
rect 229836 133900 229888 133952
rect 265256 133900 265308 133952
rect 231676 133832 231728 133884
rect 256240 133832 256292 133884
rect 282276 133832 282328 133884
rect 286232 133832 286284 133884
rect 231768 133764 231820 133816
rect 253480 133764 253532 133816
rect 230664 133696 230716 133748
rect 250812 133696 250864 133748
rect 214564 133288 214616 133340
rect 214564 133084 214616 133136
rect 261576 132608 261628 132660
rect 265164 132608 265216 132660
rect 169208 132540 169260 132592
rect 213920 132540 213972 132592
rect 257620 132540 257672 132592
rect 265992 132540 266044 132592
rect 169300 132472 169352 132524
rect 214012 132472 214064 132524
rect 242532 132472 242584 132524
rect 266176 132472 266228 132524
rect 231768 132404 231820 132456
rect 251824 132404 251876 132456
rect 282092 132404 282144 132456
rect 291200 132404 291252 132456
rect 231676 132336 231728 132388
rect 250720 132336 250772 132388
rect 282552 132336 282604 132388
rect 285772 132336 285824 132388
rect 231584 132268 231636 132320
rect 249432 132268 249484 132320
rect 250812 131248 250864 131300
rect 265992 131248 266044 131300
rect 169392 131180 169444 131232
rect 214012 131180 214064 131232
rect 253572 131180 253624 131232
rect 266176 131180 266228 131232
rect 169116 131112 169168 131164
rect 213920 131112 213972 131164
rect 230940 131044 230992 131096
rect 259092 131044 259144 131096
rect 281908 131044 281960 131096
rect 284484 131044 284536 131096
rect 231492 130976 231544 131028
rect 253388 130976 253440 131028
rect 282092 130976 282144 131028
rect 285128 130976 285180 131028
rect 231032 130772 231084 130824
rect 235632 130772 235684 130824
rect 241060 129888 241112 129940
rect 265992 129888 266044 129940
rect 180156 129820 180208 129872
rect 213920 129820 213972 129872
rect 256240 129820 256292 129872
rect 266176 129820 266228 129872
rect 171784 129752 171836 129804
rect 214012 129752 214064 129804
rect 231768 129684 231820 129736
rect 257528 129684 257580 129736
rect 282092 129616 282144 129668
rect 284852 129616 284904 129668
rect 281908 129548 281960 129600
rect 284668 129548 284720 129600
rect 231676 129480 231728 129532
rect 238300 129480 238352 129532
rect 257436 128460 257488 128512
rect 265992 128460 266044 128512
rect 173256 128392 173308 128444
rect 213920 128392 213972 128444
rect 245108 128392 245160 128444
rect 265348 128392 265400 128444
rect 169024 128324 169076 128376
rect 214012 128324 214064 128376
rect 238208 128324 238260 128376
rect 265532 128324 265584 128376
rect 265992 128324 266044 128376
rect 266176 128324 266228 128376
rect 231584 128256 231636 128308
rect 242440 128256 242492 128308
rect 231676 128188 231728 128240
rect 238484 128188 238536 128240
rect 281908 128188 281960 128240
rect 284576 128188 284628 128240
rect 231768 128120 231820 128172
rect 238116 128120 238168 128172
rect 281908 127644 281960 127696
rect 284760 127644 284812 127696
rect 247684 127100 247736 127152
rect 264152 127100 264204 127152
rect 192484 127032 192536 127084
rect 213920 127032 213972 127084
rect 245016 127032 245068 127084
rect 265532 127032 265584 127084
rect 167828 126964 167880 127016
rect 214012 126964 214064 127016
rect 239404 126964 239456 127016
rect 266176 126964 266228 127016
rect 231584 126896 231636 126948
rect 254676 126896 254728 126948
rect 454684 126896 454736 126948
rect 580172 126896 580224 126948
rect 231768 126828 231820 126880
rect 249156 126828 249208 126880
rect 231676 126760 231728 126812
rect 240968 126760 241020 126812
rect 282828 126692 282880 126744
rect 288624 126692 288676 126744
rect 230848 126216 230900 126268
rect 263232 126216 263284 126268
rect 249432 125740 249484 125792
rect 266176 125740 266228 125792
rect 168012 125672 168064 125724
rect 213920 125672 213972 125724
rect 254768 125672 254820 125724
rect 265532 125672 265584 125724
rect 167920 125604 167972 125656
rect 214012 125604 214064 125656
rect 263324 125604 263376 125656
rect 266268 125604 266320 125656
rect 231768 125536 231820 125588
rect 264428 125536 264480 125588
rect 230664 124924 230716 124976
rect 259184 124924 259236 124976
rect 230756 124856 230808 124908
rect 264704 124856 264756 124908
rect 282828 124448 282880 124500
rect 287888 124448 287940 124500
rect 259092 124312 259144 124364
rect 266176 124312 266228 124364
rect 173348 124244 173400 124296
rect 214012 124244 214064 124296
rect 261484 124244 261536 124296
rect 265348 124244 265400 124296
rect 166632 124176 166684 124228
rect 213920 124176 213972 124228
rect 247868 124176 247920 124228
rect 265164 124176 265216 124228
rect 231768 124108 231820 124160
rect 239496 124108 239548 124160
rect 231308 123496 231360 123548
rect 250996 123496 251048 123548
rect 282828 123496 282880 123548
rect 288532 123496 288584 123548
rect 231584 123428 231636 123480
rect 257712 123428 257764 123480
rect 257528 123020 257580 123072
rect 264428 123020 264480 123072
rect 256148 122952 256200 123004
rect 265164 122952 265216 123004
rect 171876 122884 171928 122936
rect 213920 122884 213972 122936
rect 242440 122884 242492 122936
rect 266176 122884 266228 122936
rect 170496 122816 170548 122868
rect 214012 122816 214064 122868
rect 240968 122816 241020 122868
rect 265440 122816 265492 122868
rect 231768 122748 231820 122800
rect 262956 122748 263008 122800
rect 231400 122680 231452 122732
rect 260564 122680 260616 122732
rect 231124 122612 231176 122664
rect 260104 122612 260156 122664
rect 231492 122068 231544 122120
rect 256424 122068 256476 122120
rect 253480 121592 253532 121644
rect 264704 121592 264756 121644
rect 181536 121524 181588 121576
rect 213920 121524 213972 121576
rect 176108 121456 176160 121508
rect 214012 121456 214064 121508
rect 260288 121456 260340 121508
rect 265532 121456 265584 121508
rect 231768 121388 231820 121440
rect 264612 121388 264664 121440
rect 231400 121320 231452 121372
rect 250628 121320 250680 121372
rect 231032 120708 231084 120760
rect 261760 120708 261812 120760
rect 258908 120232 258960 120284
rect 265532 120232 265584 120284
rect 174728 120164 174780 120216
rect 213920 120164 213972 120216
rect 250720 120164 250772 120216
rect 266176 120164 266228 120216
rect 166724 120096 166776 120148
rect 214012 120096 214064 120148
rect 249156 120096 249208 120148
rect 265440 120096 265492 120148
rect 231768 120028 231820 120080
rect 242256 120028 242308 120080
rect 230572 119960 230624 120012
rect 235540 119960 235592 120012
rect 231492 119348 231544 119400
rect 253664 119348 253716 119400
rect 170588 118804 170640 118856
rect 213920 118804 213972 118856
rect 252100 118804 252152 118856
rect 266176 118804 266228 118856
rect 180248 118736 180300 118788
rect 214012 118736 214064 118788
rect 241152 118736 241204 118788
rect 265440 118736 265492 118788
rect 238024 118668 238076 118720
rect 265532 118668 265584 118720
rect 282828 118600 282880 118652
rect 290096 118600 290148 118652
rect 282736 118532 282788 118584
rect 286140 118532 286192 118584
rect 230572 118396 230624 118448
rect 235356 118396 235408 118448
rect 231768 118260 231820 118312
rect 235448 118260 235500 118312
rect 231676 117988 231728 118040
rect 254952 117988 255004 118040
rect 265440 117988 265492 118040
rect 265900 117988 265952 118040
rect 235540 117920 235592 117972
rect 266084 117920 266136 117972
rect 265348 117512 265400 117564
rect 265808 117512 265860 117564
rect 254676 117444 254728 117496
rect 265532 117444 265584 117496
rect 244924 117376 244976 117428
rect 265900 117376 265952 117428
rect 178868 117308 178920 117360
rect 213920 117308 213972 117360
rect 229744 117308 229796 117360
rect 265808 117308 265860 117360
rect 231768 117240 231820 117292
rect 252284 117240 252336 117292
rect 282828 117240 282880 117292
rect 289084 117240 289136 117292
rect 231124 116628 231176 116680
rect 245200 116628 245252 116680
rect 234252 116560 234304 116612
rect 265440 116560 265492 116612
rect 282828 116424 282880 116476
rect 287796 116424 287848 116476
rect 238300 116152 238352 116204
rect 265900 116152 265952 116204
rect 260104 116084 260156 116136
rect 265808 116084 265860 116136
rect 173440 116016 173492 116068
rect 213920 116016 213972 116068
rect 251824 116016 251876 116068
rect 264612 116016 264664 116068
rect 166816 115948 166868 116000
rect 214012 115948 214064 116000
rect 262956 115948 263008 116000
rect 266084 115948 266136 116000
rect 231768 115880 231820 115932
rect 240876 115880 240928 115932
rect 230940 115812 230992 115864
rect 234068 115812 234120 115864
rect 234160 115200 234212 115252
rect 265348 115200 265400 115252
rect 282828 114792 282880 114844
rect 287336 114792 287388 114844
rect 174820 114588 174872 114640
rect 214012 114588 214064 114640
rect 243728 114588 243780 114640
rect 265808 114588 265860 114640
rect 170772 114520 170824 114572
rect 213920 114520 213972 114572
rect 239496 114520 239548 114572
rect 265900 114520 265952 114572
rect 231492 114452 231544 114504
rect 260472 114452 260524 114504
rect 231768 114384 231820 114436
rect 245292 114384 245344 114436
rect 282736 114316 282788 114368
rect 286048 114316 286100 114368
rect 282828 113432 282880 113484
rect 287612 113432 287664 113484
rect 246396 113296 246448 113348
rect 265808 113296 265860 113348
rect 172060 113228 172112 113280
rect 214012 113228 214064 113280
rect 245200 113228 245252 113280
rect 265900 113228 265952 113280
rect 169484 113160 169536 113212
rect 213920 113160 213972 113212
rect 235356 113160 235408 113212
rect 265808 113160 265860 113212
rect 231768 113092 231820 113144
rect 249064 113092 249116 113144
rect 231676 113024 231728 113076
rect 242348 113024 242400 113076
rect 282828 112684 282880 112736
rect 286508 112684 286560 112736
rect 168104 112412 168156 112464
rect 215116 112412 215168 112464
rect 231584 112412 231636 112464
rect 251916 112412 251968 112464
rect 252284 111936 252336 111988
rect 265808 111936 265860 111988
rect 171968 111868 172020 111920
rect 213920 111868 213972 111920
rect 250996 111868 251048 111920
rect 265532 111868 265584 111920
rect 170864 111800 170916 111852
rect 214012 111800 214064 111852
rect 242256 111800 242308 111852
rect 265900 111800 265952 111852
rect 3424 111732 3476 111784
rect 25504 111732 25556 111784
rect 168288 111732 168340 111784
rect 170680 111732 170732 111784
rect 231492 111732 231544 111784
rect 257344 111732 257396 111784
rect 231768 111664 231820 111716
rect 255964 111664 256016 111716
rect 282828 111120 282880 111172
rect 287704 111120 287756 111172
rect 282000 111052 282052 111104
rect 287244 111052 287296 111104
rect 260472 110576 260524 110628
rect 265164 110576 265216 110628
rect 256424 110508 256476 110560
rect 265808 110508 265860 110560
rect 173532 110440 173584 110492
rect 213920 110440 213972 110492
rect 240876 110440 240928 110492
rect 265900 110440 265952 110492
rect 167552 110372 167604 110424
rect 173164 110372 173216 110424
rect 231768 110372 231820 110424
rect 243636 110372 243688 110424
rect 230940 110168 230992 110220
rect 236736 110168 236788 110220
rect 282828 110032 282880 110084
rect 287060 110032 287112 110084
rect 282276 109896 282328 109948
rect 287152 109896 287204 109948
rect 231768 109420 231820 109472
rect 236828 109420 236880 109472
rect 253388 109148 253440 109200
rect 265808 109148 265860 109200
rect 177488 109080 177540 109132
rect 213920 109080 213972 109132
rect 246304 109080 246356 109132
rect 265900 109080 265952 109132
rect 174912 109012 174964 109064
rect 214012 109012 214064 109064
rect 242348 109012 242400 109064
rect 265348 109012 265400 109064
rect 167552 108944 167604 108996
rect 176016 108944 176068 108996
rect 231768 108944 231820 108996
rect 261668 108944 261720 108996
rect 282368 108944 282420 108996
rect 288992 108944 289044 108996
rect 231676 108876 231728 108928
rect 236644 108876 236696 108928
rect 281540 108604 281592 108656
rect 283380 108604 283432 108656
rect 231032 108536 231084 108588
rect 235264 108536 235316 108588
rect 249064 107856 249116 107908
rect 265808 107856 265860 107908
rect 257712 107788 257764 107840
rect 265532 107788 265584 107840
rect 255964 107720 256016 107772
rect 265808 107720 265860 107772
rect 182916 107652 182968 107704
rect 213920 107652 213972 107704
rect 231768 107584 231820 107636
rect 262864 107584 262916 107636
rect 281724 107584 281776 107636
rect 289820 107584 289872 107636
rect 231216 107516 231268 107568
rect 233884 107516 233936 107568
rect 231492 107176 231544 107228
rect 233976 107176 234028 107228
rect 230940 106904 230992 106956
rect 258724 106904 258776 106956
rect 251916 106428 251968 106480
rect 265808 106428 265860 106480
rect 176016 106360 176068 106412
rect 214012 106360 214064 106412
rect 259276 106360 259328 106412
rect 265440 106360 265492 106412
rect 173164 106292 173216 106344
rect 213920 106292 213972 106344
rect 263232 106292 263284 106344
rect 265900 106292 265952 106344
rect 231768 106156 231820 106208
rect 241244 106156 241296 106208
rect 231676 106088 231728 106140
rect 254860 106088 254912 106140
rect 230756 106020 230808 106072
rect 232688 106020 232740 106072
rect 230572 105544 230624 105596
rect 256332 105544 256384 105596
rect 282828 105068 282880 105120
rect 288900 105068 288952 105120
rect 170680 105000 170732 105052
rect 213920 105000 213972 105052
rect 250628 105000 250680 105052
rect 265808 105000 265860 105052
rect 168196 104932 168248 104984
rect 214012 104932 214064 104984
rect 166908 104864 166960 104916
rect 214104 104864 214156 104916
rect 260564 104864 260616 104916
rect 265440 104864 265492 104916
rect 231768 104796 231820 104848
rect 250904 104796 250956 104848
rect 281540 104796 281592 104848
rect 283748 104796 283800 104848
rect 230756 104660 230808 104712
rect 232504 104660 232556 104712
rect 281540 104524 281592 104576
rect 283288 104524 283340 104576
rect 230664 104116 230716 104168
rect 263140 104116 263192 104168
rect 258724 103708 258776 103760
rect 265164 103708 265216 103760
rect 263416 103572 263468 103624
rect 265808 103572 265860 103624
rect 168288 103504 168340 103556
rect 213920 103504 213972 103556
rect 235264 103504 235316 103556
rect 265348 103504 265400 103556
rect 231492 103436 231544 103488
rect 252192 103436 252244 103488
rect 282828 103436 282880 103488
rect 290004 103436 290056 103488
rect 231768 103368 231820 103420
rect 242624 103368 242676 103420
rect 282000 103232 282052 103284
rect 289268 103232 289320 103284
rect 65708 102416 65760 102468
rect 65984 102416 66036 102468
rect 246580 102348 246632 102400
rect 265440 102348 265492 102400
rect 169760 102212 169812 102264
rect 214012 102212 214064 102264
rect 257344 102212 257396 102264
rect 265808 102212 265860 102264
rect 168380 102144 168432 102196
rect 213920 102144 213972 102196
rect 231768 102076 231820 102128
rect 259000 102076 259052 102128
rect 214288 101056 214340 101108
rect 214932 101056 214984 101108
rect 259184 100852 259236 100904
rect 265532 100852 265584 100904
rect 65800 100784 65852 100836
rect 66168 100784 66220 100836
rect 263140 100784 263192 100836
rect 265900 100784 265952 100836
rect 249524 100716 249576 100768
rect 265808 100716 265860 100768
rect 565084 100648 565136 100700
rect 580172 100648 580224 100700
rect 231676 100580 231728 100632
rect 234252 100580 234304 100632
rect 282276 100240 282328 100292
rect 285956 100240 286008 100292
rect 230848 100104 230900 100156
rect 235540 100104 235592 100156
rect 231768 99900 231820 99952
rect 238392 99900 238444 99952
rect 230756 99832 230808 99884
rect 232596 99832 232648 99884
rect 254860 99492 254912 99544
rect 265808 99492 265860 99544
rect 238116 99424 238168 99476
rect 265532 99424 265584 99476
rect 233976 99356 234028 99408
rect 265900 99356 265952 99408
rect 231032 99288 231084 99340
rect 249248 99288 249300 99340
rect 166080 98812 166132 98864
rect 166632 98812 166684 98864
rect 166632 98676 166684 98728
rect 166908 98676 166960 98728
rect 233884 98608 233936 98660
rect 266084 98608 266136 98660
rect 262864 98064 262916 98116
rect 265716 98064 265768 98116
rect 169576 97996 169628 98048
rect 213920 97996 213972 98048
rect 231124 97996 231176 98048
rect 265808 97996 265860 98048
rect 3424 97588 3476 97640
rect 7564 97588 7616 97640
rect 231584 97588 231636 97640
rect 234160 97588 234212 97640
rect 231768 97316 231820 97368
rect 248420 97316 248472 97368
rect 267556 97316 267608 97368
rect 231308 97248 231360 97300
rect 237288 97248 237340 97300
rect 267280 97248 267332 97300
rect 256332 96772 256384 96824
rect 265532 96772 265584 96824
rect 236644 96704 236696 96756
rect 265624 96704 265676 96756
rect 165528 96636 165580 96688
rect 213920 96636 213972 96688
rect 232596 96636 232648 96688
rect 265900 96636 265952 96688
rect 247776 96364 247828 96416
rect 279424 96364 279476 96416
rect 250536 96296 250588 96348
rect 279332 96296 279384 96348
rect 265716 96228 265768 96280
rect 279240 96228 279292 96280
rect 166172 96092 166224 96144
rect 214104 96092 214156 96144
rect 267096 96092 267148 96144
rect 279516 96092 279568 96144
rect 165344 96024 165396 96076
rect 214012 96024 214064 96076
rect 165068 95956 165120 96008
rect 214656 95956 214708 96008
rect 165436 95888 165488 95940
rect 214196 95888 214248 95940
rect 230572 95276 230624 95328
rect 232504 95276 232556 95328
rect 165988 95208 166040 95260
rect 213920 95208 213972 95260
rect 228364 95208 228416 95260
rect 265716 95208 265768 95260
rect 267280 95140 267332 95192
rect 270960 95140 271012 95192
rect 265440 95072 265492 95124
rect 281540 95072 281592 95124
rect 65892 95004 65944 95056
rect 169760 95004 169812 95056
rect 194508 95004 194560 95056
rect 281632 95004 281684 95056
rect 66076 94936 66128 94988
rect 170680 94936 170732 94988
rect 65616 94868 65668 94920
rect 168380 94868 168432 94920
rect 65708 94800 65760 94852
rect 168288 94800 168340 94852
rect 65800 94732 65852 94784
rect 168196 94732 168248 94784
rect 128728 94528 128780 94580
rect 214380 94528 214432 94580
rect 110328 94460 110380 94512
rect 215024 94460 215076 94512
rect 151728 94120 151780 94172
rect 166448 94120 166500 94172
rect 124128 94052 124180 94104
rect 173348 94120 173400 94172
rect 117136 93984 117188 94036
rect 166724 93984 166776 94036
rect 122104 93916 122156 93968
rect 177396 93916 177448 93968
rect 118240 93848 118292 93900
rect 181536 93848 181588 93900
rect 151544 93780 151596 93832
rect 166356 93780 166408 93832
rect 166448 93780 166500 93832
rect 214564 93780 214616 93832
rect 267556 93780 267608 93832
rect 276940 93780 276992 93832
rect 119712 93712 119764 93764
rect 176108 93712 176160 93764
rect 109224 93644 109276 93696
rect 166816 93644 166868 93696
rect 107752 93576 107804 93628
rect 173440 93576 173492 93628
rect 105544 93508 105596 93560
rect 170772 93508 170824 93560
rect 102968 93440 103020 93492
rect 169484 93440 169536 93492
rect 106464 93372 106516 93424
rect 174820 93372 174872 93424
rect 104256 93304 104308 93356
rect 172060 93304 172112 93356
rect 101864 93236 101916 93288
rect 170864 93236 170916 93288
rect 90272 93168 90324 93220
rect 166632 93168 166684 93220
rect 111800 93100 111852 93152
rect 214932 93100 214984 93152
rect 125416 93032 125468 93084
rect 168012 93032 168064 93084
rect 135720 92964 135772 93016
rect 166540 92964 166592 93016
rect 151636 92896 151688 92948
rect 166264 92896 166316 92948
rect 118056 92420 118108 92472
rect 126060 92420 126112 92472
rect 84384 92352 84436 92404
rect 128728 92352 128780 92404
rect 153108 92352 153160 92404
rect 166448 92352 166500 92404
rect 88064 92284 88116 92336
rect 166172 92284 166224 92336
rect 100024 92216 100076 92268
rect 110328 92216 110380 92268
rect 114376 92216 114428 92268
rect 191104 92216 191156 92268
rect 89076 92148 89128 92200
rect 165436 92148 165488 92200
rect 105728 92080 105780 92132
rect 169392 92080 169444 92132
rect 111984 92012 112036 92064
rect 174636 92012 174688 92064
rect 108120 91944 108172 91996
rect 169300 91944 169352 91996
rect 125784 91876 125836 91928
rect 186964 91876 187016 91928
rect 109960 91808 110012 91860
rect 168104 91808 168156 91860
rect 129464 91740 129516 91792
rect 165068 91740 165120 91792
rect 169024 91740 169076 91792
rect 266084 91740 266136 91792
rect 120264 91672 120316 91724
rect 178776 91672 178828 91724
rect 134432 91604 134484 91656
rect 177304 91604 177356 91656
rect 86684 91536 86736 91588
rect 165344 91536 165396 91588
rect 94964 91468 95016 91520
rect 214288 91468 214340 91520
rect 112352 90992 112404 91044
rect 213184 90992 213236 91044
rect 91468 90924 91520 90976
rect 173164 90924 173216 90976
rect 110144 90856 110196 90908
rect 178868 90856 178920 90908
rect 113364 90788 113416 90840
rect 180248 90788 180300 90840
rect 115848 90720 115900 90772
rect 174728 90720 174780 90772
rect 110972 90652 111024 90704
rect 167736 90652 167788 90704
rect 115204 90584 115256 90636
rect 170588 90584 170640 90636
rect 132408 90516 132460 90568
rect 184204 90516 184256 90568
rect 121184 90448 121236 90500
rect 171876 90448 171928 90500
rect 115940 90380 115992 90432
rect 259092 90380 259144 90432
rect 7564 90312 7616 90364
rect 230664 90312 230716 90364
rect 121920 90244 121972 90296
rect 170496 90244 170548 90296
rect 122840 90176 122892 90228
rect 166080 90176 166132 90228
rect 126612 90108 126664 90160
rect 167920 90108 167972 90160
rect 97816 89632 97868 89684
rect 192484 89632 192536 89684
rect 75736 89564 75788 89616
rect 165988 89564 166040 89616
rect 95056 89496 95108 89548
rect 182916 89496 182968 89548
rect 93216 89428 93268 89480
rect 176016 89428 176068 89480
rect 96344 89360 96396 89412
rect 177488 89360 177540 89412
rect 97540 89292 97592 89344
rect 174912 89292 174964 89344
rect 99288 89224 99340 89276
rect 173532 89224 173584 89276
rect 100576 89156 100628 89208
rect 171968 89156 172020 89208
rect 115480 89088 115532 89140
rect 170404 89088 170456 89140
rect 122840 89020 122892 89072
rect 263324 89020 263376 89072
rect 51080 88952 51132 89004
rect 263416 88952 263468 89004
rect 113180 88884 113232 88936
rect 167644 88884 167696 88936
rect 125324 88816 125376 88868
rect 175924 88816 175976 88868
rect 86776 88272 86828 88324
rect 169576 88272 169628 88324
rect 99104 88204 99156 88256
rect 173256 88204 173308 88256
rect 128176 88136 128228 88188
rect 202144 88136 202196 88188
rect 104624 88068 104676 88120
rect 169116 88068 169168 88120
rect 123576 88000 123628 88052
rect 182824 88000 182876 88052
rect 126704 87932 126756 87984
rect 181444 87932 181496 87984
rect 133328 87864 133380 87916
rect 178684 87864 178736 87916
rect 130752 87796 130804 87848
rect 174544 87796 174596 87848
rect 60740 87660 60792 87712
rect 264796 87660 264848 87712
rect 49700 87592 49752 87644
rect 256240 87592 256292 87644
rect 195704 86912 195756 86964
rect 580172 86912 580224 86964
rect 63500 86300 63552 86352
rect 257620 86300 257672 86352
rect 64880 86232 64932 86284
rect 260564 86232 260616 86284
rect 3148 85484 3200 85536
rect 47584 85484 47636 85536
rect 67640 84872 67692 84924
rect 261576 84872 261628 84924
rect 46940 84804 46992 84856
rect 264704 84804 264756 84856
rect 70400 83512 70452 83564
rect 242532 83512 242584 83564
rect 71780 83444 71832 83496
rect 263232 83444 263284 83496
rect 78680 82152 78732 82204
rect 259276 82152 259328 82204
rect 56600 82084 56652 82136
rect 250812 82084 250864 82136
rect 89720 80724 89772 80776
rect 257712 80724 257764 80776
rect 9680 80656 9732 80708
rect 249432 80656 249484 80708
rect 93860 79364 93912 79416
rect 264612 79364 264664 79416
rect 52460 79296 52512 79348
rect 253572 79296 253624 79348
rect 107660 78004 107712 78056
rect 256424 78004 256476 78056
rect 44180 77936 44232 77988
rect 238300 77936 238352 77988
rect 110420 76576 110472 76628
rect 260472 76576 260524 76628
rect 34520 76508 34572 76560
rect 239496 76508 239548 76560
rect 85580 75216 85632 75268
rect 263048 75216 263100 75268
rect 16580 75148 16632 75200
rect 254860 75148 254912 75200
rect 118700 73856 118752 73908
rect 252284 73856 252336 73908
rect 27620 73788 27672 73840
rect 243728 73788 243780 73840
rect 253296 73108 253348 73160
rect 579988 73108 580040 73160
rect 121460 72496 121512 72548
rect 250996 72496 251048 72548
rect 22100 72428 22152 72480
rect 245200 72428 245252 72480
rect 3424 71680 3476 71732
rect 195244 71680 195296 71732
rect 118792 71000 118844 71052
rect 254768 71000 254820 71052
rect 88340 69708 88392 69760
rect 260380 69708 260432 69760
rect 26240 69640 26292 69692
rect 249524 69640 249576 69692
rect 106280 68348 106332 68400
rect 229928 68348 229980 68400
rect 29000 68280 29052 68332
rect 259184 68280 259236 68332
rect 110512 66920 110564 66972
rect 252008 66920 252060 66972
rect 33140 66852 33192 66904
rect 263140 66852 263192 66904
rect 120080 65560 120132 65612
rect 243544 65560 243596 65612
rect 40040 65492 40092 65544
rect 261668 65492 261720 65544
rect 124220 64200 124272 64252
rect 246488 64200 246540 64252
rect 2780 64132 2832 64184
rect 256332 64132 256384 64184
rect 99380 62840 99432 62892
rect 249340 62840 249392 62892
rect 62120 62772 62172 62824
rect 241152 62772 241204 62824
rect 69020 61412 69072 61464
rect 252100 61412 252152 61464
rect 42800 61344 42852 61396
rect 241060 61344 241112 61396
rect 209780 60664 209832 60716
rect 580172 60664 580224 60716
rect 111800 60052 111852 60104
rect 247868 60052 247920 60104
rect 24860 59984 24912 60036
rect 265900 59984 265952 60036
rect 3056 59304 3108 59356
rect 188344 59304 188396 59356
rect 60832 58624 60884 58676
rect 264520 58624 264572 58676
rect 80060 57264 80112 57316
rect 258908 57264 258960 57316
rect 38660 57196 38712 57248
rect 238208 57196 238260 57248
rect 93952 55904 94004 55956
rect 256148 55904 256200 55956
rect 31760 55836 31812 55888
rect 257436 55836 257488 55888
rect 98000 54544 98052 54596
rect 257528 54544 257580 54596
rect 35900 54476 35952 54528
rect 245108 54476 245160 54528
rect 104900 53116 104952 53168
rect 242440 53116 242492 53168
rect 74540 53048 74592 53100
rect 258816 53048 258868 53100
rect 81440 51756 81492 51808
rect 229836 51756 229888 51808
rect 109040 51688 109092 51740
rect 261484 51688 261536 51740
rect 102140 50396 102192 50448
rect 240968 50396 241020 50448
rect 13820 50328 13872 50380
rect 245016 50328 245068 50380
rect 91100 49036 91152 49088
rect 264428 49036 264480 49088
rect 11060 48968 11112 49020
rect 236644 48968 236696 49020
rect 86960 47608 87012 47660
rect 253480 47608 253532 47660
rect 15200 47540 15252 47592
rect 232596 47540 232648 47592
rect 84200 46180 84252 46232
rect 260288 46180 260340 46232
rect 3424 45500 3476 45552
rect 209044 45500 209096 45552
rect 92480 44820 92532 44872
rect 256056 44820 256108 44872
rect 12440 43392 12492 43444
rect 235356 43392 235408 43444
rect 77300 42032 77352 42084
rect 250720 42032 250772 42084
rect 44272 40672 44324 40724
rect 246580 40672 246632 40724
rect 96620 39380 96672 39432
rect 242348 39380 242400 39432
rect 45560 39312 45612 39364
rect 264336 39312 264388 39364
rect 73160 37884 73212 37936
rect 249156 37884 249208 37936
rect 66260 36524 66312 36576
rect 238024 36524 238076 36576
rect 59360 35164 59412 35216
rect 254676 35164 254728 35216
rect 20720 33736 20772 33788
rect 233976 33736 234028 33788
rect 3516 33056 3568 33108
rect 15844 33056 15896 33108
rect 206284 33056 206336 33108
rect 580172 33056 580224 33108
rect 17960 32376 18012 32428
rect 246396 32376 246448 32428
rect 55220 31016 55272 31068
rect 244924 31016 244976 31068
rect 48320 29588 48372 29640
rect 262956 29588 263008 29640
rect 35992 28228 36044 28280
rect 257344 28228 257396 28280
rect 8300 26868 8352 26920
rect 242256 26868 242308 26920
rect 114560 25576 114612 25628
rect 240876 25576 240928 25628
rect 41420 25508 41472 25560
rect 251824 25508 251876 25560
rect 103520 24148 103572 24200
rect 246304 24148 246356 24200
rect 19340 24080 19392 24132
rect 247684 24080 247736 24132
rect 100760 22788 100812 22840
rect 253388 22788 253440 22840
rect 23480 22720 23532 22772
rect 239404 22720 239456 22772
rect 11152 21360 11204 21412
rect 238116 21360 238168 21412
rect 3424 20612 3476 20664
rect 196624 20612 196676 20664
rect 260196 20612 260248 20664
rect 579988 20612 580040 20664
rect 77392 19932 77444 19984
rect 254584 19932 254636 19984
rect 75920 18572 75972 18624
rect 251916 18572 251968 18624
rect 85672 17280 85724 17332
rect 249064 17280 249116 17332
rect 4160 17212 4212 17264
rect 228364 17212 228416 17264
rect 83280 15920 83332 15972
rect 255964 15920 256016 15972
rect 20168 15852 20220 15904
rect 231124 15852 231176 15904
rect 54944 14424 54996 14476
rect 258724 14424 258776 14476
rect 69112 13064 69164 13116
rect 250628 13064 250680 13116
rect 103336 11772 103388 11824
rect 250444 11772 250496 11824
rect 58440 11704 58492 11756
rect 235264 11704 235316 11756
rect 117320 10344 117372 10396
rect 242164 10344 242216 10396
rect 7472 10276 7524 10328
rect 262864 10276 262916 10328
rect 114008 8984 114060 9036
rect 253204 8984 253256 9036
rect 2872 8916 2924 8968
rect 264244 8916 264296 8968
rect 96252 7624 96304 7676
rect 240784 7624 240836 7676
rect 3976 7556 4028 7608
rect 230756 7556 230808 7608
rect 3424 6808 3476 6860
rect 58624 6808 58676 6860
rect 267004 6808 267056 6860
rect 580172 6808 580224 6860
rect 38384 6128 38436 6180
rect 260104 6128 260156 6180
rect 6460 4768 6512 4820
rect 265808 4768 265860 4820
rect 572 4088 624 4140
rect 7564 4088 7616 4140
rect 125876 3612 125928 3664
rect 180064 3612 180116 3664
rect 28908 3544 28960 3596
rect 169024 3544 169076 3596
rect 44180 3476 44232 3528
rect 45100 3476 45152 3528
rect 52552 3476 52604 3528
rect 229744 3476 229796 3528
rect 232504 3476 232556 3528
rect 235816 3476 235868 3528
rect 31300 3408 31352 3460
rect 233884 3408 233936 3460
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 69020 3340 69072 3392
rect 69940 3340 69992 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 1676 3000 1728 3052
rect 3976 3000 4028 3052
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501022 3372 501735
rect 3332 501016 3384 501022
rect 3332 500958 3384 500964
rect 3054 475688 3110 475697
rect 3054 475623 3110 475632
rect 3068 474774 3096 475623
rect 3056 474768 3108 474774
rect 3056 474710 3108 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3344 448594 3372 449511
rect 3332 448588 3384 448594
rect 3332 448530 3384 448536
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3160 422346 3188 423535
rect 3148 422340 3200 422346
rect 3148 422282 3200 422288
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3054 306232 3110 306241
rect 3054 306167 3110 306176
rect 3068 298790 3096 306167
rect 3056 298784 3108 298790
rect 3056 298726 3108 298732
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3344 292602 3372 293111
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 3436 269074 3464 566879
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 3424 269068 3476 269074
rect 3424 269010 3476 269016
rect 3330 267200 3386 267209
rect 3330 267135 3386 267144
rect 3344 266626 3372 267135
rect 3332 266620 3384 266626
rect 3332 266562 3384 266568
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 253230 3464 254079
rect 3424 253224 3476 253230
rect 3424 253166 3476 253172
rect 3054 241088 3110 241097
rect 3054 241023 3110 241032
rect 3068 240174 3096 241023
rect 3056 240168 3108 240174
rect 3056 240110 3108 240116
rect 3528 239426 3556 514791
rect 3606 410544 3662 410553
rect 3606 410479 3662 410488
rect 3620 247042 3648 410479
rect 3700 286068 3752 286074
rect 3700 286010 3752 286016
rect 3608 247036 3660 247042
rect 3608 246978 3660 246984
rect 3516 239420 3568 239426
rect 3516 239362 3568 239368
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3712 149841 3740 286010
rect 6932 269006 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 699718 24348 703520
rect 40512 700330 40540 703520
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40500 700324 40552 700330
rect 40500 700266 40552 700272
rect 50344 700324 50396 700330
rect 50344 700266 50396 700272
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 26884 699712 26936 699718
rect 26884 699654 26936 699660
rect 25504 553444 25556 553450
rect 25504 553386 25556 553392
rect 10324 527196 10376 527202
rect 10324 527138 10376 527144
rect 6920 269000 6972 269006
rect 6920 268942 6972 268948
rect 7564 266620 7616 266626
rect 7564 266562 7616 266568
rect 7576 240106 7604 266562
rect 10336 262206 10364 527138
rect 15844 422340 15896 422346
rect 15844 422282 15896 422288
rect 11704 292596 11756 292602
rect 11704 292538 11756 292544
rect 10324 262200 10376 262206
rect 10324 262142 10376 262148
rect 11716 244254 11744 292538
rect 15856 291854 15884 422282
rect 15844 291848 15896 291854
rect 15844 291790 15896 291796
rect 18604 284368 18656 284374
rect 18604 284310 18656 284316
rect 15844 269136 15896 269142
rect 15844 269078 15896 269084
rect 11704 244248 11756 244254
rect 11704 244190 11756 244196
rect 7564 240100 7616 240106
rect 7564 240042 7616 240048
rect 7564 233912 7616 233918
rect 7564 233854 7616 233860
rect 3698 149832 3754 149841
rect 3698 149767 3754 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 7576 97646 7604 233854
rect 3424 97640 3476 97646
rect 3422 97608 3424 97617
rect 7564 97640 7616 97646
rect 3476 97608 3478 97617
rect 7564 97582 7616 97588
rect 3422 97543 3478 97552
rect 7564 90364 7616 90370
rect 7564 90306 7616 90312
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 2780 64184 2832 64190
rect 2780 64126 2832 64132
rect 2792 16574 2820 64126
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 4172 16574 4200 17206
rect 2792 16546 3648 16574
rect 4172 16546 5304 16574
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 584 480 612 4082
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1688 480 1716 2994
rect 2884 480 2912 8910
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 3976 7608 4028 7614
rect 3976 7550 4028 7556
rect 3988 3058 4016 7550
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 5276 480 5304 16546
rect 7472 10328 7524 10334
rect 7472 10270 7524 10276
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6472 480 6500 4762
rect 7484 3482 7512 10270
rect 7576 4146 7604 90306
rect 9680 80708 9732 80714
rect 9680 80650 9732 80656
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 8312 16574 8340 26862
rect 8312 16546 8800 16574
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8772 480 8800 16546
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 80650
rect 13820 50380 13872 50386
rect 13820 50322 13872 50328
rect 11060 49020 11112 49026
rect 11060 48962 11112 48968
rect 11072 6914 11100 48962
rect 12440 43444 12492 43450
rect 12440 43386 12492 43392
rect 11152 21412 11204 21418
rect 11152 21354 11204 21360
rect 11164 16574 11192 21354
rect 12452 16574 12480 43386
rect 13832 16574 13860 50322
rect 15200 47592 15252 47598
rect 15200 47534 15252 47540
rect 15212 16574 15240 47534
rect 15856 33114 15884 269078
rect 17224 264988 17276 264994
rect 17224 264930 17276 264936
rect 17236 215286 17264 264930
rect 17224 215280 17276 215286
rect 17224 215222 17276 215228
rect 18616 164218 18644 284310
rect 25516 264926 25544 553386
rect 26896 287706 26924 699654
rect 28264 632120 28316 632126
rect 28264 632062 28316 632068
rect 26884 287700 26936 287706
rect 26884 287642 26936 287648
rect 28276 267714 28304 632062
rect 29644 618316 29696 618322
rect 29644 618258 29696 618264
rect 29656 276010 29684 618258
rect 29644 276004 29696 276010
rect 29644 275946 29696 275952
rect 28264 267708 28316 267714
rect 28264 267650 28316 267656
rect 25504 264920 25556 264926
rect 25504 264862 25556 264868
rect 26884 258120 26936 258126
rect 26884 258062 26936 258068
rect 25504 236700 25556 236706
rect 25504 236642 25556 236648
rect 18604 164212 18656 164218
rect 18604 164154 18656 164160
rect 25516 111790 25544 236642
rect 26896 137970 26924 258062
rect 47584 253972 47636 253978
rect 47584 253914 47636 253920
rect 26884 137964 26936 137970
rect 26884 137906 26936 137912
rect 25504 111784 25556 111790
rect 25504 111726 25556 111732
rect 47596 85542 47624 253914
rect 50356 238746 50384 700266
rect 71792 294642 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 86224 474768 86276 474774
rect 86224 474710 86276 474716
rect 71780 294636 71832 294642
rect 71780 294578 71832 294584
rect 86236 287774 86264 474710
rect 88352 297430 88380 702406
rect 105464 699786 105492 703520
rect 105452 699780 105504 699786
rect 105452 699722 105504 699728
rect 108304 699780 108356 699786
rect 108304 699722 108356 699728
rect 88340 297424 88392 297430
rect 88340 297366 88392 297372
rect 86224 287768 86276 287774
rect 86224 287710 86276 287716
rect 58624 281580 58676 281586
rect 58624 281522 58676 281528
rect 50344 238740 50396 238746
rect 50344 238682 50396 238688
rect 51080 89004 51132 89010
rect 51080 88946 51132 88952
rect 49700 87644 49752 87650
rect 49700 87586 49752 87592
rect 47584 85536 47636 85542
rect 47584 85478 47636 85484
rect 46940 84856 46992 84862
rect 46940 84798 46992 84804
rect 44180 77988 44232 77994
rect 44180 77930 44232 77936
rect 34520 76560 34572 76566
rect 34520 76502 34572 76508
rect 16580 75200 16632 75206
rect 16580 75142 16632 75148
rect 15844 33108 15896 33114
rect 15844 33050 15896 33056
rect 16592 16574 16620 75142
rect 27620 73840 27672 73846
rect 27620 73782 27672 73788
rect 22100 72480 22152 72486
rect 22100 72422 22152 72428
rect 20720 33788 20772 33794
rect 20720 33730 20772 33736
rect 17960 32428 18012 32434
rect 17960 32370 18012 32376
rect 11164 16546 11928 16574
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 11072 6886 11192 6914
rect 11164 480 11192 6886
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13556 480 13584 16546
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 32370
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19352 16574 19380 24074
rect 20732 16574 20760 33730
rect 22112 16574 22140 72422
rect 26240 69692 26292 69698
rect 26240 69634 26292 69640
rect 24860 60036 24912 60042
rect 24860 59978 24912 59984
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23492 16574 23520 22714
rect 24872 16574 24900 59978
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 19444 480 19472 16546
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 15846
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 69634
rect 27632 16574 27660 73782
rect 29000 68332 29052 68338
rect 29000 68274 29052 68280
rect 29012 16574 29040 68274
rect 33140 66904 33192 66910
rect 33140 66846 33192 66852
rect 31760 55888 31812 55894
rect 31760 55830 31812 55836
rect 31772 16574 31800 55830
rect 33152 16574 33180 66846
rect 27632 16546 27752 16574
rect 29012 16546 30144 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 27724 480 27752 16546
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28920 480 28948 3538
rect 30116 480 30144 16546
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 31312 480 31340 3402
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 76502
rect 40040 65544 40092 65550
rect 40040 65486 40092 65492
rect 38660 57248 38712 57254
rect 38660 57190 38712 57196
rect 35900 54528 35952 54534
rect 35900 54470 35952 54476
rect 35912 6914 35940 54470
rect 35992 28280 36044 28286
rect 35992 28222 36044 28228
rect 36004 16574 36032 28222
rect 38672 16574 38700 57190
rect 40052 16574 40080 65486
rect 42800 61396 42852 61402
rect 42800 61338 42852 61344
rect 41420 25560 41472 25566
rect 41420 25502 41472 25508
rect 41432 16574 41460 25502
rect 36004 16546 36768 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 35912 6886 36032 6914
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 6180 38436 6186
rect 38384 6122 38436 6128
rect 38396 480 38424 6122
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 61338
rect 44192 3534 44220 77930
rect 44272 40724 44324 40730
rect 44272 40666 44324 40672
rect 44180 3528 44232 3534
rect 44180 3470 44232 3476
rect 44284 480 44312 40666
rect 45560 39364 45612 39370
rect 45560 39306 45612 39312
rect 45572 16574 45600 39306
rect 46952 16574 46980 84798
rect 48320 29640 48372 29646
rect 48320 29582 48372 29588
rect 48332 16574 48360 29582
rect 49712 16574 49740 87586
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 45100 3528 45152 3534
rect 45100 3470 45152 3476
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45112 354 45140 3470
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 88946
rect 56600 82136 56652 82142
rect 56600 82078 56652 82084
rect 52460 79348 52512 79354
rect 52460 79290 52512 79296
rect 52472 16574 52500 79290
rect 55220 31068 55272 31074
rect 55220 31010 55272 31016
rect 55232 16574 55260 31010
rect 56612 16574 56640 82078
rect 52472 16546 53328 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 52552 3528 52604 3534
rect 52552 3470 52604 3476
rect 52564 480 52592 3470
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54944 14476 54996 14482
rect 54944 14418 54996 14424
rect 54956 480 54984 14418
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58440 11756 58492 11762
rect 58440 11698 58492 11704
rect 58452 480 58480 11698
rect 58636 6866 58664 281522
rect 108316 238678 108344 699722
rect 136652 251190 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234724 703582 235028 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700126 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 169772 702406 170352 702434
rect 154120 700120 154172 700126
rect 154120 700062 154172 700068
rect 155224 700120 155276 700126
rect 155224 700062 155276 700068
rect 155236 286346 155264 700062
rect 156604 670744 156656 670750
rect 156604 670686 156656 670692
rect 156616 286414 156644 670686
rect 156604 286408 156656 286414
rect 156604 286350 156656 286356
rect 155224 286340 155276 286346
rect 155224 286282 155276 286288
rect 169772 273222 169800 702406
rect 195796 700664 195848 700670
rect 195796 700606 195848 700612
rect 175924 462392 175976 462398
rect 175924 462334 175976 462340
rect 169760 273216 169812 273222
rect 169760 273158 169812 273164
rect 136640 251184 136692 251190
rect 136640 251126 136692 251132
rect 175936 240038 175964 462334
rect 195336 397520 195388 397526
rect 195336 397462 195388 397468
rect 194416 285932 194468 285938
rect 194416 285874 194468 285880
rect 192484 284708 192536 284714
rect 192484 284650 192536 284656
rect 188344 284436 188396 284442
rect 188344 284378 188396 284384
rect 175924 240032 175976 240038
rect 175924 239974 175976 239980
rect 108304 238672 108356 238678
rect 108304 238614 108356 238620
rect 180064 229764 180116 229770
rect 180064 229706 180116 229712
rect 114008 178492 114060 178498
rect 114008 178434 114060 178440
rect 169300 178492 169352 178498
rect 169300 178434 169352 178440
rect 110696 178356 110748 178362
rect 110696 178298 110748 178304
rect 97816 178152 97868 178158
rect 97816 178094 97868 178100
rect 97828 176769 97856 178094
rect 110052 178084 110104 178090
rect 110052 178026 110104 178032
rect 103336 177404 103388 177410
rect 103336 177346 103388 177352
rect 103348 176769 103376 177346
rect 107016 176928 107068 176934
rect 107016 176870 107068 176876
rect 107028 176769 107056 176870
rect 108120 176860 108172 176866
rect 108120 176802 108172 176808
rect 108132 176769 108160 176802
rect 110064 176769 110092 178026
rect 110708 176769 110736 178298
rect 112628 178288 112680 178294
rect 112628 178230 112680 178236
rect 112640 176769 112668 178230
rect 114020 176769 114048 178434
rect 114376 178424 114428 178430
rect 114376 178366 114428 178372
rect 114388 176769 114416 178366
rect 169208 178356 169260 178362
rect 169208 178298 169260 178304
rect 148232 178220 148284 178226
rect 148232 178162 148284 178168
rect 134524 177540 134576 177546
rect 134524 177482 134576 177488
rect 133144 177472 133196 177478
rect 133144 177414 133196 177420
rect 129740 177404 129792 177410
rect 129740 177346 129792 177352
rect 130936 177404 130988 177410
rect 130936 177346 130988 177352
rect 127992 177336 128044 177342
rect 127992 177278 128044 177284
rect 124496 177200 124548 177206
rect 124496 177142 124548 177148
rect 122288 177132 122340 177138
rect 122288 177074 122340 177080
rect 120816 177064 120868 177070
rect 120816 177006 120868 177012
rect 118424 176996 118476 177002
rect 118424 176938 118476 176944
rect 116952 176792 117004 176798
rect 97814 176760 97870 176769
rect 97814 176695 97870 176704
rect 103334 176760 103390 176769
rect 103334 176695 103390 176704
rect 107014 176760 107070 176769
rect 107014 176695 107070 176704
rect 108118 176760 108174 176769
rect 108118 176695 108174 176704
rect 110050 176760 110106 176769
rect 110050 176695 110106 176704
rect 110694 176760 110750 176769
rect 110694 176695 110750 176704
rect 112626 176760 112682 176769
rect 112626 176695 112682 176704
rect 114006 176760 114062 176769
rect 114006 176695 114062 176704
rect 114374 176760 114430 176769
rect 114374 176695 114430 176704
rect 115846 176760 115902 176769
rect 115846 176695 115848 176704
rect 115900 176695 115902 176704
rect 116950 176760 116952 176769
rect 118436 176769 118464 176938
rect 120828 176769 120856 177006
rect 122300 176769 122328 177074
rect 124508 176769 124536 177142
rect 128004 176769 128032 177278
rect 129464 177268 129516 177274
rect 129464 177210 129516 177216
rect 129476 176769 129504 177210
rect 117004 176760 117006 176769
rect 116950 176695 117006 176704
rect 118422 176760 118478 176769
rect 118422 176695 118478 176704
rect 120814 176760 120870 176769
rect 120814 176695 120870 176704
rect 122286 176760 122342 176769
rect 122286 176695 122342 176704
rect 124494 176760 124550 176769
rect 124494 176695 124550 176704
rect 127990 176760 128046 176769
rect 127990 176695 128046 176704
rect 129462 176760 129518 176769
rect 129462 176695 129518 176704
rect 115848 176666 115900 176672
rect 125692 176656 125744 176662
rect 125692 176598 125744 176604
rect 123116 176520 123168 176526
rect 123116 176462 123168 176468
rect 119436 176452 119488 176458
rect 119436 176394 119488 176400
rect 104624 176384 104676 176390
rect 104624 176326 104676 176332
rect 98368 176316 98420 176322
rect 98368 176258 98420 176264
rect 98380 175409 98408 176258
rect 100760 176248 100812 176254
rect 100760 176190 100812 176196
rect 99472 176180 99524 176186
rect 99472 176122 99524 176128
rect 99484 175409 99512 176122
rect 100772 175409 100800 176190
rect 102048 175976 102100 175982
rect 102048 175918 102100 175924
rect 102060 175409 102088 175918
rect 104636 175409 104664 176326
rect 105728 176112 105780 176118
rect 105728 176054 105780 176060
rect 105740 175409 105768 176054
rect 98366 175400 98422 175409
rect 98366 175335 98422 175344
rect 99470 175400 99526 175409
rect 99470 175335 99526 175344
rect 100758 175400 100814 175409
rect 100758 175335 100814 175344
rect 102046 175400 102102 175409
rect 102046 175335 102102 175344
rect 104622 175400 104678 175409
rect 104622 175335 104678 175344
rect 105726 175400 105782 175409
rect 105726 175335 105782 175344
rect 119448 175001 119476 176394
rect 123128 175001 123156 176462
rect 125704 175001 125732 176598
rect 129752 176050 129780 177346
rect 130948 176769 130976 177346
rect 133156 176769 133184 177414
rect 134536 176769 134564 177482
rect 148244 176769 148272 178162
rect 165160 177540 165212 177546
rect 165160 177482 165212 177488
rect 130934 176760 130990 176769
rect 130934 176695 130990 176704
rect 133142 176760 133198 176769
rect 133142 176695 133198 176704
rect 134522 176760 134578 176769
rect 134522 176695 134578 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 135720 176588 135772 176594
rect 135720 176530 135772 176536
rect 129740 176044 129792 176050
rect 129740 175986 129792 175992
rect 128176 175908 128228 175914
rect 128176 175850 128228 175856
rect 128188 175409 128216 175850
rect 132040 175840 132092 175846
rect 132040 175782 132092 175788
rect 132052 175409 132080 175782
rect 135732 175545 135760 176530
rect 158904 175772 158956 175778
rect 158904 175714 158956 175720
rect 135718 175536 135774 175545
rect 135718 175471 135774 175480
rect 158916 175409 158944 175714
rect 128174 175400 128230 175409
rect 128174 175335 128230 175344
rect 132038 175400 132094 175409
rect 132038 175335 132094 175344
rect 158902 175400 158958 175409
rect 158902 175335 158958 175344
rect 165172 175234 165200 177482
rect 165252 177472 165304 177478
rect 165252 177414 165304 177420
rect 165160 175228 165212 175234
rect 165160 175170 165212 175176
rect 165264 175166 165292 177414
rect 165712 177404 165764 177410
rect 165712 177346 165764 177352
rect 165344 177336 165396 177342
rect 165344 177278 165396 177284
rect 165252 175160 165304 175166
rect 165252 175102 165304 175108
rect 119434 174992 119490 175001
rect 119434 174927 119490 174936
rect 123114 174992 123170 175001
rect 123114 174927 123170 174936
rect 125690 174992 125746 175001
rect 125690 174927 125746 174936
rect 165356 174554 165384 177278
rect 165436 175908 165488 175914
rect 165436 175850 165488 175856
rect 165344 174548 165396 174554
rect 165344 174490 165396 174496
rect 165448 172514 165476 175850
rect 165528 175840 165580 175846
rect 165528 175782 165580 175788
rect 165540 173874 165568 175782
rect 165528 173868 165580 173874
rect 165528 173810 165580 173816
rect 165724 173806 165752 177346
rect 165804 177268 165856 177274
rect 165804 177210 165856 177216
rect 165712 173800 165764 173806
rect 165712 173742 165764 173748
rect 165436 172508 165488 172514
rect 165436 172450 165488 172456
rect 165816 172446 165844 177210
rect 166356 177200 166408 177206
rect 166356 177142 166408 177148
rect 166264 176316 166316 176322
rect 166264 176258 166316 176264
rect 165804 172440 165856 172446
rect 165804 172382 165856 172388
rect 166276 155922 166304 176258
rect 166368 169658 166396 177142
rect 167828 176928 167880 176934
rect 167828 176870 167880 176876
rect 166540 176656 166592 176662
rect 166540 176598 166592 176604
rect 166448 176520 166500 176526
rect 166448 176462 166500 176468
rect 166460 169726 166488 176462
rect 166552 171086 166580 176598
rect 167736 176452 167788 176458
rect 167736 176394 167788 176400
rect 167644 176384 167696 176390
rect 167644 176326 167696 176332
rect 166632 175772 166684 175778
rect 166632 175714 166684 175720
rect 166540 171080 166592 171086
rect 166540 171022 166592 171028
rect 166448 169720 166500 169726
rect 166448 169662 166500 169668
rect 166356 169652 166408 169658
rect 166356 169594 166408 169600
rect 166264 155916 166316 155922
rect 166264 155858 166316 155864
rect 166448 153332 166500 153338
rect 166448 153274 166500 153280
rect 166264 153264 166316 153270
rect 166264 153206 166316 153212
rect 66166 129296 66222 129305
rect 66166 129231 66222 129240
rect 66074 128072 66130 128081
rect 66074 128007 66130 128016
rect 65982 126304 66038 126313
rect 65982 126239 66038 126248
rect 65890 123584 65946 123593
rect 65890 123519 65946 123528
rect 65798 122632 65854 122641
rect 65798 122567 65854 122576
rect 65812 103514 65840 122567
rect 65628 103486 65840 103514
rect 65628 94926 65656 103486
rect 65708 102468 65760 102474
rect 65708 102410 65760 102416
rect 65616 94920 65668 94926
rect 65616 94862 65668 94868
rect 65720 94858 65748 102410
rect 65800 100836 65852 100842
rect 65800 100778 65852 100784
rect 65708 94852 65760 94858
rect 65708 94794 65760 94800
rect 65812 94790 65840 100778
rect 65904 95062 65932 123519
rect 65996 102474 66024 126239
rect 65984 102468 66036 102474
rect 65984 102410 66036 102416
rect 65982 102368 66038 102377
rect 65982 102303 66038 102312
rect 65892 95056 65944 95062
rect 65892 94998 65944 95004
rect 65800 94784 65852 94790
rect 65800 94726 65852 94732
rect 65996 94489 66024 102303
rect 66088 94994 66116 128007
rect 66180 100842 66208 129231
rect 67638 125216 67694 125225
rect 67638 125151 67694 125160
rect 66168 100836 66220 100842
rect 66168 100778 66220 100784
rect 66166 100736 66222 100745
rect 66166 100671 66222 100680
rect 66076 94988 66128 94994
rect 66076 94930 66128 94936
rect 66180 94625 66208 100671
rect 67652 94761 67680 125151
rect 67822 120864 67878 120873
rect 67822 120799 67878 120808
rect 67836 94897 67864 120799
rect 166080 98864 166132 98870
rect 166080 98806 166132 98812
rect 165528 96688 165580 96694
rect 165528 96630 165580 96636
rect 165344 96076 165396 96082
rect 165344 96018 165396 96024
rect 165068 96008 165120 96014
rect 165068 95950 165120 95956
rect 67822 94888 67878 94897
rect 67822 94823 67878 94832
rect 67638 94752 67694 94761
rect 67638 94687 67694 94696
rect 66166 94616 66222 94625
rect 66166 94551 66222 94560
rect 128728 94580 128780 94586
rect 128728 94522 128780 94528
rect 110328 94512 110380 94518
rect 65982 94480 66038 94489
rect 110328 94454 110380 94460
rect 65982 94415 66038 94424
rect 109224 93696 109276 93702
rect 102966 93664 103022 93673
rect 102966 93599 103022 93608
rect 104254 93664 104310 93673
rect 104254 93599 104310 93608
rect 105542 93664 105598 93673
rect 105542 93599 105598 93608
rect 106462 93664 106518 93673
rect 106462 93599 106518 93608
rect 107750 93664 107806 93673
rect 107750 93599 107752 93608
rect 90270 93528 90326 93537
rect 90270 93463 90326 93472
rect 101862 93528 101918 93537
rect 102980 93498 103008 93599
rect 101862 93463 101918 93472
rect 102968 93492 103020 93498
rect 90284 93226 90312 93463
rect 101876 93294 101904 93463
rect 102968 93434 103020 93440
rect 104268 93362 104296 93599
rect 105556 93566 105584 93599
rect 105544 93560 105596 93566
rect 105544 93502 105596 93508
rect 106476 93430 106504 93599
rect 107804 93599 107806 93608
rect 109222 93664 109224 93673
rect 109276 93664 109278 93673
rect 109222 93599 109278 93608
rect 107752 93570 107804 93576
rect 106464 93424 106516 93430
rect 106464 93366 106516 93372
rect 104256 93356 104308 93362
rect 104256 93298 104308 93304
rect 101864 93288 101916 93294
rect 101864 93230 101916 93236
rect 110142 93256 110198 93265
rect 90272 93220 90324 93226
rect 110142 93191 110198 93200
rect 90272 93162 90324 93168
rect 84382 92440 84438 92449
rect 84382 92375 84384 92384
rect 84436 92375 84438 92384
rect 86682 92440 86738 92449
rect 86682 92375 86738 92384
rect 88062 92440 88118 92449
rect 88062 92375 88118 92384
rect 89074 92440 89130 92449
rect 89074 92375 89130 92384
rect 91466 92440 91522 92449
rect 91466 92375 91522 92384
rect 94962 92440 95018 92449
rect 94962 92375 95018 92384
rect 100022 92440 100078 92449
rect 100022 92375 100078 92384
rect 105726 92440 105782 92449
rect 105726 92375 105782 92384
rect 108118 92440 108174 92449
rect 108118 92375 108174 92384
rect 109958 92440 110014 92449
rect 109958 92375 110014 92384
rect 84384 92346 84436 92352
rect 75734 91760 75790 91769
rect 75734 91695 75790 91704
rect 75748 89622 75776 91695
rect 86696 91594 86724 92375
rect 88076 92342 88104 92375
rect 88064 92336 88116 92342
rect 88064 92278 88116 92284
rect 89088 92206 89116 92375
rect 89076 92200 89128 92206
rect 89076 92142 89128 92148
rect 86684 91588 86736 91594
rect 86684 91530 86736 91536
rect 86774 91216 86830 91225
rect 86774 91151 86830 91160
rect 75736 89616 75788 89622
rect 75736 89558 75788 89564
rect 86788 88330 86816 91151
rect 91480 90982 91508 92375
rect 93214 91624 93270 91633
rect 93214 91559 93270 91568
rect 91468 90976 91520 90982
rect 91468 90918 91520 90924
rect 93228 89486 93256 91559
rect 94976 91526 95004 92375
rect 100036 92274 100064 92375
rect 100024 92268 100076 92274
rect 100024 92210 100076 92216
rect 105740 92138 105768 92375
rect 105728 92132 105780 92138
rect 105728 92074 105780 92080
rect 108132 92002 108160 92375
rect 108120 91996 108172 92002
rect 108120 91938 108172 91944
rect 109972 91866 110000 92375
rect 109960 91860 110012 91866
rect 109960 91802 110012 91808
rect 95054 91760 95110 91769
rect 95054 91695 95110 91704
rect 97814 91760 97870 91769
rect 97814 91695 97870 91704
rect 100574 91760 100630 91769
rect 100574 91695 100630 91704
rect 94964 91520 95016 91526
rect 94964 91462 95016 91468
rect 95068 89554 95096 91695
rect 96342 91624 96398 91633
rect 96342 91559 96398 91568
rect 97538 91624 97594 91633
rect 97538 91559 97594 91568
rect 95056 89548 95108 89554
rect 95056 89490 95108 89496
rect 93216 89480 93268 89486
rect 93216 89422 93268 89428
rect 96356 89418 96384 91559
rect 96344 89412 96396 89418
rect 96344 89354 96396 89360
rect 97552 89350 97580 91559
rect 97828 89690 97856 91695
rect 99286 91624 99342 91633
rect 99286 91559 99342 91568
rect 99102 91216 99158 91225
rect 99102 91151 99158 91160
rect 97816 89684 97868 89690
rect 97816 89626 97868 89632
rect 97540 89344 97592 89350
rect 97540 89286 97592 89292
rect 86776 88324 86828 88330
rect 86776 88266 86828 88272
rect 99116 88262 99144 91151
rect 99300 89282 99328 91559
rect 99288 89276 99340 89282
rect 99288 89218 99340 89224
rect 100588 89214 100616 91695
rect 104622 91216 104678 91225
rect 104622 91151 104678 91160
rect 100576 89208 100628 89214
rect 100576 89150 100628 89156
rect 99104 88256 99156 88262
rect 99104 88198 99156 88204
rect 104636 88126 104664 91151
rect 110156 90914 110184 93191
rect 110340 92274 110368 94454
rect 124126 94208 124182 94217
rect 124126 94143 124182 94152
rect 124140 94110 124168 94143
rect 124128 94104 124180 94110
rect 117134 94072 117190 94081
rect 117134 94007 117136 94016
rect 117188 94007 117190 94016
rect 122102 94072 122158 94081
rect 124128 94046 124180 94052
rect 122102 94007 122158 94016
rect 117136 93978 117188 93984
rect 122116 93974 122144 94007
rect 122104 93968 122156 93974
rect 118238 93936 118294 93945
rect 122104 93910 122156 93916
rect 118238 93871 118240 93880
rect 118292 93871 118294 93880
rect 118240 93842 118292 93848
rect 119712 93764 119764 93770
rect 119712 93706 119764 93712
rect 119724 93673 119752 93706
rect 119710 93664 119766 93673
rect 119710 93599 119766 93608
rect 111798 93528 111854 93537
rect 111798 93463 111854 93472
rect 125414 93528 125470 93537
rect 125414 93463 125470 93472
rect 111812 93158 111840 93463
rect 111800 93152 111852 93158
rect 111800 93094 111852 93100
rect 125428 93090 125456 93463
rect 128174 93256 128230 93265
rect 128174 93191 128230 93200
rect 126058 93120 126114 93129
rect 125416 93084 125468 93090
rect 126058 93055 126114 93064
rect 125416 93026 125468 93032
rect 113178 92576 113234 92585
rect 113178 92511 113234 92520
rect 110970 92440 111026 92449
rect 110970 92375 111026 92384
rect 111982 92440 112038 92449
rect 111982 92375 112038 92384
rect 112350 92440 112406 92449
rect 112350 92375 112406 92384
rect 110328 92268 110380 92274
rect 110328 92210 110380 92216
rect 110144 90908 110196 90914
rect 110144 90850 110196 90856
rect 110984 90710 111012 92375
rect 111996 92070 112024 92375
rect 111984 92064 112036 92070
rect 111984 92006 112036 92012
rect 112364 91050 112392 92375
rect 112352 91044 112404 91050
rect 112352 90986 112404 90992
rect 110972 90704 111024 90710
rect 110972 90646 111024 90652
rect 113192 88942 113220 92511
rect 126072 92478 126100 93055
rect 118056 92472 118108 92478
rect 113362 92440 113418 92449
rect 113362 92375 113418 92384
rect 114374 92440 114430 92449
rect 114374 92375 114430 92384
rect 115202 92440 115258 92449
rect 115202 92375 115258 92384
rect 115846 92440 115902 92449
rect 115846 92375 115902 92384
rect 118054 92440 118056 92449
rect 126060 92472 126112 92478
rect 118108 92440 118110 92449
rect 118054 92375 118110 92384
rect 120262 92440 120318 92449
rect 120262 92375 120318 92384
rect 121182 92440 121238 92449
rect 121182 92375 121238 92384
rect 125782 92440 125838 92449
rect 126060 92414 126112 92420
rect 125782 92375 125838 92384
rect 113376 90846 113404 92375
rect 114388 92274 114416 92375
rect 114376 92268 114428 92274
rect 114376 92210 114428 92216
rect 113364 90840 113416 90846
rect 113364 90782 113416 90788
rect 115216 90642 115244 92375
rect 115478 91488 115534 91497
rect 115478 91423 115534 91432
rect 115204 90636 115256 90642
rect 115204 90578 115256 90584
rect 115492 89146 115520 91423
rect 115860 90778 115888 92375
rect 120276 91730 120304 92375
rect 120264 91724 120316 91730
rect 120264 91666 120316 91672
rect 115848 90772 115900 90778
rect 115848 90714 115900 90720
rect 121196 90506 121224 92375
rect 125796 91934 125824 92375
rect 125784 91928 125836 91934
rect 121918 91896 121974 91905
rect 125784 91870 125836 91876
rect 126610 91896 126666 91905
rect 121918 91831 121974 91840
rect 126610 91831 126666 91840
rect 121184 90500 121236 90506
rect 121184 90442 121236 90448
rect 115940 90432 115992 90438
rect 115940 90374 115992 90380
rect 115480 89140 115532 89146
rect 115480 89082 115532 89088
rect 113180 88936 113232 88942
rect 113180 88878 113232 88884
rect 104624 88120 104676 88126
rect 104624 88062 104676 88068
rect 60740 87712 60792 87718
rect 60740 87654 60792 87660
rect 59360 35216 59412 35222
rect 59360 35158 59412 35164
rect 58624 6860 58676 6866
rect 58624 6802 58676 6808
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 35158
rect 60752 3398 60780 87654
rect 63500 86352 63552 86358
rect 63500 86294 63552 86300
rect 62120 62824 62172 62830
rect 62120 62766 62172 62772
rect 60832 58676 60884 58682
rect 60832 58618 60884 58624
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 58618
rect 62132 16574 62160 62766
rect 63512 16574 63540 86294
rect 64880 86284 64932 86290
rect 64880 86226 64932 86232
rect 64892 16574 64920 86226
rect 67640 84924 67692 84930
rect 67640 84866 67692 84872
rect 66260 36576 66312 36582
rect 66260 36518 66312 36524
rect 66272 16574 66300 36518
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 84866
rect 70400 83564 70452 83570
rect 70400 83506 70452 83512
rect 69020 61464 69072 61470
rect 69020 61406 69072 61412
rect 69032 3398 69060 61406
rect 70412 16574 70440 83506
rect 71780 83496 71832 83502
rect 71780 83438 71832 83444
rect 71792 16574 71820 83438
rect 78680 82204 78732 82210
rect 78680 82146 78732 82152
rect 74540 53100 74592 53106
rect 74540 53042 74592 53048
rect 73160 37936 73212 37942
rect 73160 37878 73212 37884
rect 73172 16574 73200 37878
rect 74552 16574 74580 53042
rect 77300 42084 77352 42090
rect 77300 42026 77352 42032
rect 75920 18624 75972 18630
rect 75920 18566 75972 18572
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69112 13116 69164 13122
rect 69112 13058 69164 13064
rect 69020 3392 69072 3398
rect 69020 3334 69072 3340
rect 69124 480 69152 13058
rect 69940 3392 69992 3398
rect 69940 3334 69992 3340
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3334
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 18566
rect 77312 6914 77340 42026
rect 77392 19984 77444 19990
rect 77392 19926 77444 19932
rect 77404 16574 77432 19926
rect 78692 16574 78720 82146
rect 89720 80776 89772 80782
rect 89720 80718 89772 80724
rect 85580 75268 85632 75274
rect 85580 75210 85632 75216
rect 80060 57316 80112 57322
rect 80060 57258 80112 57264
rect 80072 16574 80100 57258
rect 81440 51808 81492 51814
rect 81440 51750 81492 51756
rect 81452 16574 81480 51750
rect 84200 46232 84252 46238
rect 84200 46174 84252 46180
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83280 15972 83332 15978
rect 83280 15914 83332 15920
rect 83292 480 83320 15914
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 46174
rect 85592 6914 85620 75210
rect 88340 69760 88392 69766
rect 88340 69702 88392 69708
rect 86960 47660 87012 47666
rect 86960 47602 87012 47608
rect 85672 17332 85724 17338
rect 85672 17274 85724 17280
rect 85684 16574 85712 17274
rect 86972 16574 87000 47602
rect 88352 16574 88380 69702
rect 89732 16574 89760 80718
rect 93860 79416 93912 79422
rect 93860 79358 93912 79364
rect 91100 49088 91152 49094
rect 91100 49030 91152 49036
rect 91112 16574 91140 49030
rect 92480 44872 92532 44878
rect 92480 44814 92532 44820
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 44814
rect 93872 6914 93900 79358
rect 107660 78056 107712 78062
rect 107660 77998 107712 78004
rect 106280 68400 106332 68406
rect 106280 68342 106332 68348
rect 99380 62892 99432 62898
rect 99380 62834 99432 62840
rect 93952 55956 94004 55962
rect 93952 55898 94004 55904
rect 93964 16574 93992 55898
rect 98000 54596 98052 54602
rect 98000 54538 98052 54544
rect 96620 39432 96672 39438
rect 96620 39374 96672 39380
rect 96632 16574 96660 39374
rect 98012 16574 98040 54538
rect 99392 16574 99420 62834
rect 104900 53168 104952 53174
rect 104900 53110 104952 53116
rect 102140 50448 102192 50454
rect 102140 50390 102192 50396
rect 100760 22840 100812 22846
rect 100760 22782 100812 22788
rect 93964 16546 94728 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 96252 7676 96304 7682
rect 96252 7618 96304 7624
rect 96264 480 96292 7618
rect 97460 480 97488 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 22782
rect 102152 16574 102180 50390
rect 103520 24200 103572 24206
rect 103520 24142 103572 24148
rect 103532 16574 103560 24142
rect 104912 16574 104940 53110
rect 106292 16574 106320 68342
rect 107672 16574 107700 77998
rect 110420 76628 110472 76634
rect 110420 76570 110472 76576
rect 109040 51740 109092 51746
rect 109040 51682 109092 51688
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102244 480 102272 16546
rect 103336 11824 103388 11830
rect 103336 11766 103388 11772
rect 103348 480 103376 11766
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 51682
rect 110432 3398 110460 76570
rect 110512 66972 110564 66978
rect 110512 66914 110564 66920
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 66914
rect 111800 60104 111852 60110
rect 111800 60046 111852 60052
rect 111812 16574 111840 60046
rect 114560 25628 114612 25634
rect 114560 25570 114612 25576
rect 114572 16574 114600 25570
rect 115952 16574 115980 90374
rect 121932 90302 121960 91831
rect 122838 91488 122894 91497
rect 122838 91423 122894 91432
rect 125322 91488 125378 91497
rect 125322 91423 125378 91432
rect 121920 90296 121972 90302
rect 121920 90238 121972 90244
rect 122852 90234 122880 91423
rect 123574 91216 123630 91225
rect 123574 91151 123630 91160
rect 122840 90228 122892 90234
rect 122840 90170 122892 90176
rect 122840 89072 122892 89078
rect 122840 89014 122892 89020
rect 118700 73908 118752 73914
rect 118700 73850 118752 73856
rect 111812 16546 112392 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114008 9036 114060 9042
rect 114008 8978 114060 8984
rect 114020 480 114048 8978
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 117320 10396 117372 10402
rect 117320 10338 117372 10344
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 10338
rect 118712 6914 118740 73850
rect 121460 72548 121512 72554
rect 121460 72490 121512 72496
rect 118792 71052 118844 71058
rect 118792 70994 118844 71000
rect 118804 16574 118832 70994
rect 120080 65612 120132 65618
rect 120080 65554 120132 65560
rect 120092 16574 120120 65554
rect 121472 16574 121500 72490
rect 122852 16574 122880 89014
rect 123588 88058 123616 91151
rect 125336 88874 125364 91423
rect 126624 90166 126652 91831
rect 126702 91216 126758 91225
rect 126702 91151 126758 91160
rect 126612 90160 126664 90166
rect 126612 90102 126664 90108
rect 125324 88868 125376 88874
rect 125324 88810 125376 88816
rect 123576 88052 123628 88058
rect 123576 87994 123628 88000
rect 126716 87990 126744 91151
rect 128188 88194 128216 93191
rect 128740 92410 128768 94522
rect 151634 94344 151690 94353
rect 151634 94279 151690 94288
rect 151542 93936 151598 93945
rect 151542 93871 151598 93880
rect 151556 93838 151584 93871
rect 151544 93832 151596 93838
rect 151544 93774 151596 93780
rect 135718 93392 135774 93401
rect 135718 93327 135774 93336
rect 135732 93022 135760 93327
rect 135720 93016 135772 93022
rect 135720 92958 135772 92964
rect 151648 92954 151676 94279
rect 151728 94172 151780 94178
rect 151728 94114 151780 94120
rect 151740 94081 151768 94114
rect 151726 94072 151782 94081
rect 151726 94007 151782 94016
rect 151636 92948 151688 92954
rect 151636 92890 151688 92896
rect 129462 92440 129518 92449
rect 128728 92404 128780 92410
rect 129462 92375 129518 92384
rect 132406 92440 132462 92449
rect 132406 92375 132462 92384
rect 134430 92440 134486 92449
rect 134430 92375 134486 92384
rect 153106 92440 153162 92449
rect 153106 92375 153108 92384
rect 128728 92346 128780 92352
rect 129476 91798 129504 92375
rect 129464 91792 129516 91798
rect 129464 91734 129516 91740
rect 130750 91216 130806 91225
rect 130750 91151 130806 91160
rect 128176 88188 128228 88194
rect 128176 88130 128228 88136
rect 126704 87984 126756 87990
rect 126704 87926 126756 87932
rect 130764 87854 130792 91151
rect 132420 90574 132448 92375
rect 134444 91662 134472 92375
rect 153160 92375 153162 92384
rect 153108 92346 153160 92352
rect 165080 91798 165108 95950
rect 165068 91792 165120 91798
rect 165068 91734 165120 91740
rect 134432 91656 134484 91662
rect 134432 91598 134484 91604
rect 165356 91594 165384 96018
rect 165436 95940 165488 95946
rect 165436 95882 165488 95888
rect 165448 92206 165476 95882
rect 165540 94489 165568 96630
rect 165988 95260 166040 95266
rect 165988 95202 166040 95208
rect 165526 94480 165582 94489
rect 165526 94415 165582 94424
rect 165436 92200 165488 92206
rect 165436 92142 165488 92148
rect 165344 91588 165396 91594
rect 165344 91530 165396 91536
rect 133326 91216 133382 91225
rect 133326 91151 133382 91160
rect 132408 90568 132460 90574
rect 132408 90510 132460 90516
rect 133340 87922 133368 91151
rect 166000 89622 166028 95202
rect 166092 90234 166120 98806
rect 166172 96144 166224 96150
rect 166172 96086 166224 96092
rect 166184 92342 166212 96086
rect 166276 92954 166304 153206
rect 166356 151836 166408 151842
rect 166356 151778 166408 151784
rect 166368 93838 166396 151778
rect 166460 94178 166488 153274
rect 166644 149054 166672 175714
rect 167656 160070 167684 176326
rect 167748 167006 167776 176394
rect 167840 170406 167868 176870
rect 169116 176180 169168 176186
rect 169116 176122 169168 176128
rect 169022 171592 169078 171601
rect 169022 171527 169078 171536
rect 167828 170400 167880 170406
rect 167828 170342 167880 170348
rect 167736 167000 167788 167006
rect 167736 166942 167788 166948
rect 167644 160064 167696 160070
rect 167644 160006 167696 160012
rect 169036 150414 169064 171527
rect 169128 157350 169156 176122
rect 169220 162858 169248 178298
rect 169312 164218 169340 178434
rect 170588 178424 170640 178430
rect 170588 178366 170640 178372
rect 170404 178152 170456 178158
rect 170404 178094 170456 178100
rect 169392 177132 169444 177138
rect 169392 177074 169444 177080
rect 169404 168366 169432 177074
rect 169392 168360 169444 168366
rect 169392 168302 169444 168308
rect 169300 164212 169352 164218
rect 169300 164154 169352 164160
rect 169208 162852 169260 162858
rect 169208 162794 169260 162800
rect 169116 157344 169168 157350
rect 169116 157286 169168 157292
rect 170416 155854 170444 178094
rect 170496 176248 170548 176254
rect 170496 176190 170548 176196
rect 170508 157282 170536 176190
rect 170600 165578 170628 178366
rect 173256 178288 173308 178294
rect 173256 178230 173308 178236
rect 170680 177064 170732 177070
rect 170680 177006 170732 177012
rect 170692 168298 170720 177006
rect 173164 175976 173216 175982
rect 173164 175918 173216 175924
rect 170680 168292 170732 168298
rect 170680 168234 170732 168240
rect 170588 165572 170640 165578
rect 170588 165514 170640 165520
rect 173176 158710 173204 175918
rect 173268 164150 173296 178230
rect 174636 176996 174688 177002
rect 174636 176938 174688 176944
rect 174544 176860 174596 176866
rect 174544 176802 174596 176808
rect 173256 164144 173308 164150
rect 173256 164086 173308 164092
rect 174556 161430 174584 176802
rect 174648 166938 174676 176938
rect 175924 176112 175976 176118
rect 175924 176054 175976 176060
rect 174636 166932 174688 166938
rect 174636 166874 174688 166880
rect 174544 161424 174596 161430
rect 174544 161366 174596 161372
rect 175936 160002 175964 176054
rect 175924 159996 175976 160002
rect 175924 159938 175976 159944
rect 173164 158704 173216 158710
rect 173164 158646 173216 158652
rect 170496 157276 170548 157282
rect 170496 157218 170548 157224
rect 170404 155848 170456 155854
rect 170404 155790 170456 155796
rect 176016 151088 176068 151094
rect 176016 151030 176068 151036
rect 173164 150476 173216 150482
rect 173164 150418 173216 150424
rect 169024 150408 169076 150414
rect 169024 150350 169076 150356
rect 166632 149048 166684 149054
rect 166632 148990 166684 148996
rect 166540 147688 166592 147694
rect 166540 147630 166592 147636
rect 166448 94172 166500 94178
rect 166448 94114 166500 94120
rect 166356 93832 166408 93838
rect 166356 93774 166408 93780
rect 166448 93832 166500 93838
rect 166448 93774 166500 93780
rect 166264 92948 166316 92954
rect 166264 92890 166316 92896
rect 166460 92410 166488 93774
rect 166552 93022 166580 147630
rect 170680 137284 170732 137290
rect 170680 137226 170732 137232
rect 170404 136672 170456 136678
rect 170404 136614 170456 136620
rect 167644 135312 167696 135318
rect 167644 135254 167696 135260
rect 166632 124228 166684 124234
rect 166632 124170 166684 124176
rect 166644 98870 166672 124170
rect 166724 120148 166776 120154
rect 166724 120090 166776 120096
rect 166632 98864 166684 98870
rect 166632 98806 166684 98812
rect 166632 98728 166684 98734
rect 166632 98670 166684 98676
rect 166644 93226 166672 98670
rect 166736 94042 166764 120090
rect 166816 116000 166868 116006
rect 166816 115942 166868 115948
rect 166724 94036 166776 94042
rect 166724 93978 166776 93984
rect 166828 93702 166856 115942
rect 167552 110424 167604 110430
rect 167552 110366 167604 110372
rect 167564 110129 167592 110366
rect 167550 110120 167606 110129
rect 167550 110055 167606 110064
rect 167552 108996 167604 109002
rect 167552 108938 167604 108944
rect 167564 108769 167592 108938
rect 167550 108760 167606 108769
rect 167550 108695 167606 108704
rect 166908 104916 166960 104922
rect 166908 104858 166960 104864
rect 166920 98734 166948 104858
rect 166908 98728 166960 98734
rect 166908 98670 166960 98676
rect 166816 93696 166868 93702
rect 166816 93638 166868 93644
rect 166632 93220 166684 93226
rect 166632 93162 166684 93168
rect 166540 93016 166592 93022
rect 166540 92958 166592 92964
rect 166448 92404 166500 92410
rect 166448 92346 166500 92352
rect 166172 92336 166224 92342
rect 166172 92278 166224 92284
rect 166080 90228 166132 90234
rect 166080 90170 166132 90176
rect 165988 89616 166040 89622
rect 165988 89558 166040 89564
rect 167656 88942 167684 135254
rect 167736 133952 167788 133958
rect 167736 133894 167788 133900
rect 167748 90710 167776 133894
rect 169208 132592 169260 132598
rect 169208 132534 169260 132540
rect 169116 131164 169168 131170
rect 169116 131106 169168 131112
rect 169024 128376 169076 128382
rect 169024 128318 169076 128324
rect 167828 127016 167880 127022
rect 167828 126958 167880 126964
rect 167840 92313 167868 126958
rect 168012 125724 168064 125730
rect 168012 125666 168064 125672
rect 167920 125656 167972 125662
rect 167920 125598 167972 125604
rect 167826 92304 167882 92313
rect 167826 92239 167882 92248
rect 167736 90704 167788 90710
rect 167736 90646 167788 90652
rect 167932 90166 167960 125598
rect 168024 93090 168052 125666
rect 168104 112464 168156 112470
rect 168104 112406 168156 112412
rect 168012 93084 168064 93090
rect 168012 93026 168064 93032
rect 168116 91866 168144 112406
rect 168288 111784 168340 111790
rect 168286 111752 168288 111761
rect 168340 111752 168342 111761
rect 168286 111687 168342 111696
rect 168196 104984 168248 104990
rect 168196 104926 168248 104932
rect 168208 94790 168236 104926
rect 168288 103556 168340 103562
rect 168288 103498 168340 103504
rect 168300 94858 168328 103498
rect 168380 102196 168432 102202
rect 168380 102138 168432 102144
rect 168392 94926 168420 102138
rect 168380 94920 168432 94926
rect 168380 94862 168432 94868
rect 168288 94852 168340 94858
rect 168288 94794 168340 94800
rect 168196 94784 168248 94790
rect 168196 94726 168248 94732
rect 169036 93809 169064 128318
rect 169022 93800 169078 93809
rect 169022 93735 169078 93744
rect 168104 91860 168156 91866
rect 168104 91802 168156 91808
rect 169024 91792 169076 91798
rect 169024 91734 169076 91740
rect 167920 90160 167972 90166
rect 167920 90102 167972 90108
rect 167644 88936 167696 88942
rect 167644 88878 167696 88884
rect 133328 87916 133380 87922
rect 133328 87858 133380 87864
rect 130752 87848 130804 87854
rect 130752 87790 130804 87796
rect 124220 64252 124272 64258
rect 124220 64194 124272 64200
rect 124232 16574 124260 64194
rect 118804 16546 119936 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 118712 6886 118832 6914
rect 118804 480 118832 6886
rect 119908 480 119936 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 125876 3664 125928 3670
rect 125876 3606 125928 3612
rect 125888 480 125916 3606
rect 169036 3602 169064 91734
rect 169128 88126 169156 131106
rect 169220 92041 169248 132534
rect 169300 132524 169352 132530
rect 169300 132466 169352 132472
rect 169206 92032 169262 92041
rect 169312 92002 169340 132466
rect 169392 131232 169444 131238
rect 169392 131174 169444 131180
rect 169404 92138 169432 131174
rect 169484 113212 169536 113218
rect 169484 113154 169536 113160
rect 169496 93498 169524 113154
rect 169760 102264 169812 102270
rect 169760 102206 169812 102212
rect 169576 98048 169628 98054
rect 169576 97990 169628 97996
rect 169484 93492 169536 93498
rect 169484 93434 169536 93440
rect 169392 92132 169444 92138
rect 169392 92074 169444 92080
rect 169206 91967 169262 91976
rect 169300 91996 169352 92002
rect 169300 91938 169352 91944
rect 169588 88330 169616 97990
rect 169772 95062 169800 102206
rect 169760 95056 169812 95062
rect 169760 94998 169812 95004
rect 170416 89146 170444 136614
rect 170496 122868 170548 122874
rect 170496 122810 170548 122816
rect 170508 90302 170536 122810
rect 170588 118856 170640 118862
rect 170588 118798 170640 118804
rect 170600 90642 170628 118798
rect 170692 111790 170720 137226
rect 171784 129804 171836 129810
rect 171784 129746 171836 129752
rect 170772 114572 170824 114578
rect 170772 114514 170824 114520
rect 170680 111784 170732 111790
rect 170680 111726 170732 111732
rect 170680 105052 170732 105058
rect 170680 104994 170732 105000
rect 170692 94994 170720 104994
rect 170680 94988 170732 94994
rect 170680 94930 170732 94936
rect 170784 93566 170812 114514
rect 170864 111852 170916 111858
rect 170864 111794 170916 111800
rect 170772 93560 170824 93566
rect 170772 93502 170824 93508
rect 170876 93294 170904 111794
rect 170864 93288 170916 93294
rect 170864 93230 170916 93236
rect 171796 92177 171824 129746
rect 171876 122936 171928 122942
rect 171876 122878 171928 122884
rect 171782 92168 171838 92177
rect 171782 92103 171838 92112
rect 170588 90636 170640 90642
rect 170588 90578 170640 90584
rect 171888 90506 171916 122878
rect 172060 113280 172112 113286
rect 172060 113222 172112 113228
rect 171968 111920 172020 111926
rect 171968 111862 172020 111868
rect 171876 90500 171928 90506
rect 171876 90442 171928 90448
rect 170496 90296 170548 90302
rect 170496 90238 170548 90244
rect 171980 89214 172008 111862
rect 172072 93362 172100 113222
rect 173176 110430 173204 150418
rect 174544 144968 174596 144974
rect 174544 144910 174596 144916
rect 173256 128444 173308 128450
rect 173256 128386 173308 128392
rect 173164 110424 173216 110430
rect 173164 110366 173216 110372
rect 173164 106344 173216 106350
rect 173164 106286 173216 106292
rect 172060 93356 172112 93362
rect 172060 93298 172112 93304
rect 173176 90982 173204 106286
rect 173164 90976 173216 90982
rect 173164 90918 173216 90924
rect 171968 89208 172020 89214
rect 171968 89150 172020 89156
rect 170404 89140 170456 89146
rect 170404 89082 170456 89088
rect 169576 88324 169628 88330
rect 169576 88266 169628 88272
rect 173268 88262 173296 128386
rect 173348 124296 173400 124302
rect 173348 124238 173400 124244
rect 173360 94178 173388 124238
rect 173440 116068 173492 116074
rect 173440 116010 173492 116016
rect 173348 94172 173400 94178
rect 173348 94114 173400 94120
rect 173452 93634 173480 116010
rect 173532 110492 173584 110498
rect 173532 110434 173584 110440
rect 173440 93628 173492 93634
rect 173440 93570 173492 93576
rect 173544 89282 173572 110434
rect 173532 89276 173584 89282
rect 173532 89218 173584 89224
rect 173256 88256 173308 88262
rect 173256 88198 173308 88204
rect 169116 88120 169168 88126
rect 169116 88062 169168 88068
rect 174556 87854 174584 144910
rect 175924 140820 175976 140826
rect 175924 140762 175976 140768
rect 174636 135380 174688 135386
rect 174636 135322 174688 135328
rect 174648 92070 174676 135322
rect 174728 120216 174780 120222
rect 174728 120158 174780 120164
rect 174636 92064 174688 92070
rect 174636 92006 174688 92012
rect 174740 90778 174768 120158
rect 174820 114640 174872 114646
rect 174820 114582 174872 114588
rect 174832 93430 174860 114582
rect 174912 109064 174964 109070
rect 174912 109006 174964 109012
rect 174820 93424 174872 93430
rect 174820 93366 174872 93372
rect 174728 90772 174780 90778
rect 174728 90714 174780 90720
rect 174924 89350 174952 109006
rect 174912 89344 174964 89350
rect 174912 89286 174964 89292
rect 175936 88874 175964 140762
rect 176028 109002 176056 151030
rect 178684 146396 178736 146402
rect 178684 146338 178736 146344
rect 177304 146328 177356 146334
rect 177304 146270 177356 146276
rect 176108 121508 176160 121514
rect 176108 121450 176160 121456
rect 176016 108996 176068 109002
rect 176016 108938 176068 108944
rect 176016 106412 176068 106418
rect 176016 106354 176068 106360
rect 176028 89486 176056 106354
rect 176120 93770 176148 121450
rect 176108 93764 176160 93770
rect 176108 93706 176160 93712
rect 177316 91662 177344 146270
rect 177396 139460 177448 139466
rect 177396 139402 177448 139408
rect 177408 93974 177436 139402
rect 177488 109132 177540 109138
rect 177488 109074 177540 109080
rect 177396 93968 177448 93974
rect 177396 93910 177448 93916
rect 177304 91656 177356 91662
rect 177304 91598 177356 91604
rect 176016 89480 176068 89486
rect 176016 89422 176068 89428
rect 177500 89418 177528 109074
rect 177488 89412 177540 89418
rect 177488 89354 177540 89360
rect 175924 88868 175976 88874
rect 175924 88810 175976 88816
rect 178696 87922 178724 146338
rect 178776 139528 178828 139534
rect 178776 139470 178828 139476
rect 178788 91730 178816 139470
rect 178868 117360 178920 117366
rect 178868 117302 178920 117308
rect 178776 91724 178828 91730
rect 178776 91666 178828 91672
rect 178880 90914 178908 117302
rect 178868 90908 178920 90914
rect 178868 90850 178920 90856
rect 178684 87916 178736 87922
rect 178684 87858 178736 87864
rect 174544 87848 174596 87854
rect 174544 87790 174596 87796
rect 180076 3670 180104 229706
rect 184204 145036 184256 145042
rect 184204 144978 184256 144984
rect 181444 142180 181496 142186
rect 181444 142122 181496 142128
rect 180156 129872 180208 129878
rect 180156 129814 180208 129820
rect 180168 91361 180196 129814
rect 180248 118788 180300 118794
rect 180248 118730 180300 118736
rect 180154 91352 180210 91361
rect 180154 91287 180210 91296
rect 180260 90846 180288 118730
rect 180248 90840 180300 90846
rect 180248 90782 180300 90788
rect 181456 87990 181484 142122
rect 182824 140888 182876 140894
rect 182824 140830 182876 140836
rect 181536 121576 181588 121582
rect 181536 121518 181588 121524
rect 181548 93906 181576 121518
rect 181536 93900 181588 93906
rect 181536 93842 181588 93848
rect 182836 88058 182864 140830
rect 182916 107704 182968 107710
rect 182916 107646 182968 107652
rect 182928 89554 182956 107646
rect 184216 90574 184244 144978
rect 186964 142248 187016 142254
rect 186964 142190 187016 142196
rect 186976 91934 187004 142190
rect 186964 91928 187016 91934
rect 186964 91870 187016 91876
rect 184204 90568 184256 90574
rect 184204 90510 184256 90516
rect 182916 89548 182968 89554
rect 182916 89490 182968 89496
rect 182824 88052 182876 88058
rect 182824 87994 182876 88000
rect 181444 87984 181496 87990
rect 181444 87926 181496 87932
rect 188356 59362 188384 284378
rect 191104 253224 191156 253230
rect 191104 253166 191156 253172
rect 191116 238474 191144 253166
rect 191104 238468 191156 238474
rect 191104 238410 191156 238416
rect 192496 189038 192524 284650
rect 193128 280220 193180 280226
rect 193128 280162 193180 280168
rect 193036 278792 193088 278798
rect 193036 278734 193088 278740
rect 192944 266416 192996 266422
rect 192944 266358 192996 266364
rect 192852 265056 192904 265062
rect 192852 264998 192904 265004
rect 192484 189032 192536 189038
rect 192484 188974 192536 188980
rect 192864 180033 192892 264998
rect 192850 180024 192906 180033
rect 192850 179959 192906 179968
rect 192484 178084 192536 178090
rect 192484 178026 192536 178032
rect 191104 176792 191156 176798
rect 191104 176734 191156 176740
rect 191116 166870 191144 176734
rect 191104 166864 191156 166870
rect 191104 166806 191156 166812
rect 192496 162790 192524 178026
rect 192956 177342 192984 266358
rect 193048 180402 193076 278734
rect 193036 180396 193088 180402
rect 193036 180338 193088 180344
rect 192944 177336 192996 177342
rect 192944 177278 192996 177284
rect 193140 176662 193168 280162
rect 194324 276072 194376 276078
rect 194324 276014 194376 276020
rect 194232 256760 194284 256766
rect 194232 256702 194284 256708
rect 194140 252612 194192 252618
rect 194140 252554 194192 252560
rect 194152 182850 194180 252554
rect 194140 182844 194192 182850
rect 194140 182786 194192 182792
rect 194244 180169 194272 256702
rect 194230 180160 194286 180169
rect 194230 180095 194286 180104
rect 193128 176656 193180 176662
rect 193128 176598 193180 176604
rect 194336 175982 194364 276014
rect 194428 180606 194456 285874
rect 195244 284640 195296 284646
rect 195244 284582 195296 284588
rect 194508 271924 194560 271930
rect 194508 271866 194560 271872
rect 194416 180600 194468 180606
rect 194416 180542 194468 180548
rect 194324 175976 194376 175982
rect 194324 175918 194376 175924
rect 192484 162784 192536 162790
rect 192484 162726 192536 162732
rect 191104 135448 191156 135454
rect 191104 135390 191156 135396
rect 191116 92274 191144 135390
rect 192484 127084 192536 127090
rect 192484 127026 192536 127032
rect 191104 92268 191156 92274
rect 191104 92210 191156 92216
rect 192496 89690 192524 127026
rect 194520 95062 194548 271866
rect 195152 258664 195204 258670
rect 195152 258606 195204 258612
rect 195164 177585 195192 258606
rect 195150 177576 195206 177585
rect 195150 177511 195206 177520
rect 194508 95056 194560 95062
rect 194508 94998 194560 95004
rect 192484 89684 192536 89690
rect 192484 89626 192536 89632
rect 195256 71738 195284 284582
rect 195348 238406 195376 397462
rect 195428 286204 195480 286210
rect 195428 286146 195480 286152
rect 195336 238400 195388 238406
rect 195336 238342 195388 238348
rect 195440 180538 195468 286146
rect 195612 286136 195664 286142
rect 195612 286078 195664 286084
rect 195520 285728 195572 285734
rect 195520 285670 195572 285676
rect 195428 180532 195480 180538
rect 195428 180474 195480 180480
rect 195532 180470 195560 285670
rect 195520 180464 195572 180470
rect 195520 180406 195572 180412
rect 195624 177750 195652 286078
rect 195704 254040 195756 254046
rect 195704 253982 195756 253988
rect 195612 177744 195664 177750
rect 195612 177686 195664 177692
rect 195716 86970 195744 253982
rect 195808 244186 195836 700606
rect 198648 700596 198700 700602
rect 198648 700538 198700 700544
rect 197268 700460 197320 700466
rect 197268 700402 197320 700408
rect 195888 700324 195940 700330
rect 195888 700266 195940 700272
rect 195796 244180 195848 244186
rect 195796 244122 195848 244128
rect 195796 241528 195848 241534
rect 195796 241470 195848 241476
rect 195808 177818 195836 241470
rect 195900 238338 195928 700266
rect 197176 456816 197228 456822
rect 197176 456758 197228 456764
rect 196716 371272 196768 371278
rect 196716 371214 196768 371220
rect 196624 285252 196676 285258
rect 196624 285194 196676 285200
rect 196440 263628 196492 263634
rect 196440 263570 196492 263576
rect 196348 248532 196400 248538
rect 196348 248474 196400 248480
rect 195888 238332 195940 238338
rect 195888 238274 195940 238280
rect 196360 177954 196388 248474
rect 196452 178022 196480 263570
rect 196532 247104 196584 247110
rect 196532 247046 196584 247052
rect 196440 178016 196492 178022
rect 196440 177958 196492 177964
rect 196348 177948 196400 177954
rect 196348 177890 196400 177896
rect 195796 177812 195848 177818
rect 195796 177754 195848 177760
rect 196544 177682 196572 247046
rect 196532 177676 196584 177682
rect 196532 177618 196584 177624
rect 195704 86964 195756 86970
rect 195704 86906 195756 86912
rect 195244 71732 195296 71738
rect 195244 71674 195296 71680
rect 188344 59356 188396 59362
rect 188344 59298 188396 59304
rect 196636 20670 196664 285194
rect 196728 239834 196756 371214
rect 197084 286000 197136 286006
rect 197084 285942 197136 285948
rect 196992 285864 197044 285870
rect 196992 285806 197044 285812
rect 196900 285796 196952 285802
rect 196900 285738 196952 285744
rect 196806 257408 196862 257417
rect 196806 257343 196862 257352
rect 196716 239828 196768 239834
rect 196716 239770 196768 239776
rect 196820 180674 196848 257343
rect 196912 180742 196940 285738
rect 196900 180736 196952 180742
rect 196900 180678 196952 180684
rect 196808 180668 196860 180674
rect 196808 180610 196860 180616
rect 197004 177886 197032 285806
rect 196992 177880 197044 177886
rect 196992 177822 197044 177828
rect 197096 176526 197124 285942
rect 197188 241641 197216 456758
rect 197280 247353 197308 700402
rect 198556 510672 198608 510678
rect 198556 510614 198608 510620
rect 198372 289128 198424 289134
rect 198372 289070 198424 289076
rect 198278 282976 198334 282985
rect 198278 282911 198334 282920
rect 197358 281616 197414 281625
rect 197358 281551 197360 281560
rect 197412 281551 197414 281560
rect 197360 281522 197412 281528
rect 197358 280256 197414 280265
rect 197358 280191 197360 280200
rect 197412 280191 197414 280200
rect 197360 280162 197412 280168
rect 197358 279440 197414 279449
rect 197358 279375 197414 279384
rect 197372 278798 197400 279375
rect 197360 278792 197412 278798
rect 197360 278734 197412 278740
rect 197450 277264 197506 277273
rect 197450 277199 197506 277208
rect 197464 276078 197492 277199
rect 197452 276072 197504 276078
rect 197452 276014 197504 276020
rect 197360 276004 197412 276010
rect 197360 275946 197412 275952
rect 197372 275913 197400 275946
rect 197358 275904 197414 275913
rect 197358 275839 197414 275848
rect 198186 274544 198242 274553
rect 198186 274479 198242 274488
rect 197360 273216 197412 273222
rect 197360 273158 197412 273164
rect 197372 272377 197400 273158
rect 197450 272912 197506 272921
rect 197450 272847 197506 272856
rect 197358 272368 197414 272377
rect 197358 272303 197414 272312
rect 197464 271930 197492 272847
rect 197452 271924 197504 271930
rect 197452 271866 197504 271872
rect 197358 269376 197414 269385
rect 197358 269311 197414 269320
rect 197372 269142 197400 269311
rect 197360 269136 197412 269142
rect 197360 269078 197412 269084
rect 197452 269068 197504 269074
rect 197452 269010 197504 269016
rect 197360 269000 197412 269006
rect 197360 268942 197412 268948
rect 197372 268025 197400 268942
rect 197464 268841 197492 269010
rect 197450 268832 197506 268841
rect 197450 268767 197506 268776
rect 197358 268016 197414 268025
rect 197358 267951 197414 267960
rect 197360 267708 197412 267714
rect 197360 267650 197412 267656
rect 197372 266665 197400 267650
rect 197450 267200 197506 267209
rect 197450 267135 197506 267144
rect 197358 266656 197414 266665
rect 197358 266591 197414 266600
rect 197464 266422 197492 267135
rect 197452 266416 197504 266422
rect 197452 266358 197504 266364
rect 197450 265840 197506 265849
rect 197450 265775 197506 265784
rect 197358 265296 197414 265305
rect 197358 265231 197414 265240
rect 197372 265062 197400 265231
rect 197360 265056 197412 265062
rect 197360 264998 197412 265004
rect 197464 264994 197492 265775
rect 197452 264988 197504 264994
rect 197452 264930 197504 264936
rect 197360 264920 197412 264926
rect 197360 264862 197412 264868
rect 197372 264489 197400 264862
rect 197358 264480 197414 264489
rect 197358 264415 197414 264424
rect 197358 263664 197414 263673
rect 197358 263599 197360 263608
rect 197412 263599 197414 263608
rect 197360 263570 197412 263576
rect 197360 262200 197412 262206
rect 197360 262142 197412 262148
rect 197372 261497 197400 262142
rect 197358 261488 197414 261497
rect 197358 261423 197414 261432
rect 197450 259312 197506 259321
rect 197450 259247 197506 259256
rect 197358 258768 197414 258777
rect 197358 258703 197414 258712
rect 197372 258126 197400 258703
rect 197464 258670 197492 259247
rect 197452 258664 197504 258670
rect 197452 258606 197504 258612
rect 197360 258120 197412 258126
rect 197360 258062 197412 258068
rect 197358 257952 197414 257961
rect 197358 257887 197414 257896
rect 197372 256766 197400 257887
rect 197360 256760 197412 256766
rect 197360 256702 197412 256708
rect 198094 256592 198150 256601
rect 198094 256527 198150 256536
rect 197450 255232 197506 255241
rect 197450 255167 197506 255176
rect 197358 254416 197414 254425
rect 197358 254351 197414 254360
rect 197372 253978 197400 254351
rect 197464 254046 197492 255167
rect 197452 254040 197504 254046
rect 197452 253982 197504 253988
rect 197360 253972 197412 253978
rect 197360 253914 197412 253920
rect 197726 253600 197782 253609
rect 197726 253535 197782 253544
rect 197358 253056 197414 253065
rect 197358 252991 197414 253000
rect 197372 252618 197400 252991
rect 197360 252612 197412 252618
rect 197360 252554 197412 252560
rect 197360 251184 197412 251190
rect 197360 251126 197412 251132
rect 197372 250073 197400 251126
rect 197358 250064 197414 250073
rect 197358 249999 197414 250008
rect 197634 249520 197690 249529
rect 197634 249455 197690 249464
rect 197542 248704 197598 248713
rect 197542 248639 197598 248648
rect 197556 248538 197584 248639
rect 197544 248532 197596 248538
rect 197544 248474 197596 248480
rect 197266 247344 197322 247353
rect 197266 247279 197322 247288
rect 197360 247036 197412 247042
rect 197360 246978 197412 246984
rect 197372 245993 197400 246978
rect 197358 245984 197414 245993
rect 197358 245919 197414 245928
rect 197360 244248 197412 244254
rect 197360 244190 197412 244196
rect 197372 243817 197400 244190
rect 197452 244180 197504 244186
rect 197452 244122 197504 244128
rect 197358 243808 197414 243817
rect 197358 243743 197414 243752
rect 197464 243001 197492 244122
rect 197450 242992 197506 243001
rect 197450 242927 197506 242936
rect 197174 241632 197230 241641
rect 197174 241567 197230 241576
rect 197648 237182 197676 249455
rect 197636 237176 197688 237182
rect 197636 237118 197688 237124
rect 197740 235278 197768 253535
rect 197910 251696 197966 251705
rect 197910 251631 197966 251640
rect 197728 235272 197780 235278
rect 197728 235214 197780 235220
rect 197924 233889 197952 251631
rect 198002 247888 198058 247897
rect 198002 247823 198058 247832
rect 198016 247110 198044 247823
rect 198004 247104 198056 247110
rect 198004 247046 198056 247052
rect 198002 242176 198058 242185
rect 198002 242111 198058 242120
rect 198016 241534 198044 242111
rect 198004 241528 198056 241534
rect 198004 241470 198056 241476
rect 197910 233880 197966 233889
rect 197910 233815 197966 233824
rect 198108 232529 198136 256527
rect 198200 239562 198228 274479
rect 198188 239556 198240 239562
rect 198188 239498 198240 239504
rect 198292 232665 198320 282911
rect 198384 255785 198412 289070
rect 198568 280809 198596 510614
rect 198660 283801 198688 700538
rect 200120 404388 200172 404394
rect 200120 404330 200172 404336
rect 200132 284118 200160 404330
rect 201512 293282 201540 702986
rect 218992 700330 219020 703520
rect 234620 700392 234672 700398
rect 234620 700334 234672 700340
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 212908 696992 212960 696998
rect 212908 696934 212960 696940
rect 204904 448588 204956 448594
rect 204904 448530 204956 448536
rect 201500 293276 201552 293282
rect 201500 293218 201552 293224
rect 204916 288386 204944 448530
rect 209964 351960 210016 351966
rect 209964 351902 210016 351908
rect 209044 291848 209096 291854
rect 209044 291790 209096 291796
rect 204904 288380 204956 288386
rect 204904 288322 204956 288328
rect 208124 288380 208176 288386
rect 208124 288322 208176 288328
rect 201316 287972 201368 287978
rect 201316 287914 201368 287920
rect 200762 285832 200818 285841
rect 200762 285767 200818 285776
rect 200132 284090 200422 284118
rect 200776 284104 200804 285767
rect 201328 284104 201356 287914
rect 202236 287904 202288 287910
rect 202236 287846 202288 287852
rect 201684 285116 201736 285122
rect 201684 285058 201736 285064
rect 201696 284104 201724 285058
rect 202248 284104 202276 287846
rect 202788 286408 202840 286414
rect 202788 286350 202840 286356
rect 207572 286408 207624 286414
rect 207572 286350 207624 286356
rect 202800 284104 202828 286350
rect 204260 286340 204312 286346
rect 204260 286282 204312 286288
rect 203708 286136 203760 286142
rect 203708 286078 203760 286084
rect 203156 285864 203208 285870
rect 203156 285806 203208 285812
rect 203168 284104 203196 285806
rect 203720 284104 203748 286078
rect 204272 284104 204300 286282
rect 207020 286204 207072 286210
rect 207020 286146 207072 286152
rect 205180 286136 205232 286142
rect 205180 286078 205232 286084
rect 204628 285932 204680 285938
rect 204628 285874 204680 285880
rect 204640 284104 204668 285874
rect 205192 284104 205220 286078
rect 206100 286068 206152 286074
rect 206100 286010 206152 286016
rect 205548 285728 205600 285734
rect 205548 285670 205600 285676
rect 205560 284104 205588 285670
rect 206112 284104 206140 286010
rect 206650 284744 206706 284753
rect 206650 284679 206706 284688
rect 206664 284104 206692 284679
rect 207032 284104 207060 286146
rect 207584 284104 207612 286350
rect 208136 284104 208164 288322
rect 208492 286476 208544 286482
rect 208492 286418 208544 286424
rect 208504 284104 208532 286418
rect 209056 284104 209084 291790
rect 209412 286612 209464 286618
rect 209412 286554 209464 286560
rect 209424 284104 209452 286554
rect 209976 284104 210004 351902
rect 211988 287224 212040 287230
rect 211988 287166 212040 287172
rect 210884 286272 210936 286278
rect 210884 286214 210936 286220
rect 210516 285796 210568 285802
rect 210516 285738 210568 285744
rect 210528 284104 210556 285738
rect 210896 284104 210924 286214
rect 211436 285932 211488 285938
rect 211436 285874 211488 285880
rect 211448 284104 211476 285874
rect 212000 284104 212028 287166
rect 212356 284776 212408 284782
rect 212356 284718 212408 284724
rect 212368 284104 212396 284718
rect 212920 284104 212948 696934
rect 223028 670744 223080 670750
rect 223028 670686 223080 670692
rect 213460 418192 213512 418198
rect 213460 418134 213512 418140
rect 213472 284104 213500 418134
rect 214564 318844 214616 318850
rect 214564 318786 214616 318792
rect 214576 291854 214604 318786
rect 218612 295996 218664 296002
rect 218612 295938 218664 295944
rect 214564 291848 214616 291854
rect 214564 291790 214616 291796
rect 216220 288652 216272 288658
rect 216220 288594 216272 288600
rect 214380 288516 214432 288522
rect 214380 288458 214432 288464
rect 213828 284368 213880 284374
rect 213828 284310 213880 284316
rect 213840 284104 213868 284310
rect 214392 284104 214420 288458
rect 215300 286340 215352 286346
rect 215300 286282 215352 286288
rect 214748 285048 214800 285054
rect 214748 284990 214800 284996
rect 214760 284104 214788 284990
rect 215312 284104 215340 286282
rect 215850 285696 215906 285705
rect 215850 285631 215906 285640
rect 215864 284104 215892 285631
rect 216232 284104 216260 288594
rect 218244 287700 218296 287706
rect 218244 287642 218296 287648
rect 217324 287564 217376 287570
rect 217324 287506 217376 287512
rect 216772 287496 216824 287502
rect 216772 287438 216824 287444
rect 216784 284104 216812 287438
rect 217336 284104 217364 287506
rect 217692 286000 217744 286006
rect 217692 285942 217744 285948
rect 217704 284104 217732 285942
rect 218256 284104 218284 287642
rect 218624 284104 218652 295938
rect 222476 288720 222528 288726
rect 222476 288662 222528 288668
rect 220084 288584 220136 288590
rect 220084 288526 220136 288532
rect 219164 286544 219216 286550
rect 219164 286486 219216 286492
rect 219176 284104 219204 286486
rect 219714 284472 219770 284481
rect 219714 284407 219770 284416
rect 219728 284104 219756 284407
rect 220096 284104 220124 288526
rect 220636 287836 220688 287842
rect 220636 287778 220688 287784
rect 220648 284104 220676 287778
rect 222108 287292 222160 287298
rect 222108 287234 222160 287240
rect 221554 286104 221610 286113
rect 221554 286039 221610 286048
rect 221186 285968 221242 285977
rect 221186 285903 221242 285912
rect 221200 284104 221228 285903
rect 221568 284104 221596 286039
rect 222120 284104 222148 287234
rect 222488 284104 222516 288662
rect 223040 284104 223068 670686
rect 233884 656940 233936 656946
rect 233884 656882 233936 656888
rect 224224 605872 224276 605878
rect 224224 605814 224276 605820
rect 224236 288386 224264 605814
rect 225972 563100 226024 563106
rect 225972 563042 226024 563048
rect 224500 288788 224552 288794
rect 224500 288730 224552 288736
rect 224224 288380 224276 288386
rect 224224 288322 224276 288328
rect 223580 284912 223632 284918
rect 223580 284854 223632 284860
rect 223592 284104 223620 284854
rect 223948 284708 224000 284714
rect 223948 284650 224000 284656
rect 223960 284104 223988 284650
rect 224512 284104 224540 288730
rect 225420 288380 225472 288386
rect 225420 288322 225472 288328
rect 225052 284844 225104 284850
rect 225052 284786 225104 284792
rect 225064 284104 225092 284786
rect 225432 284104 225460 288322
rect 225984 284104 226012 563042
rect 226984 357468 227036 357474
rect 226984 357410 227036 357416
rect 226996 288386 227024 357410
rect 232504 345092 232556 345098
rect 232504 345034 232556 345040
rect 226984 288380 227036 288386
rect 226984 288322 227036 288328
rect 228364 288380 228416 288386
rect 228364 288322 228416 288328
rect 226890 286240 226946 286249
rect 226890 286175 226946 286184
rect 226524 285728 226576 285734
rect 226524 285670 226576 285676
rect 226536 284104 226564 285670
rect 226904 284104 226932 286175
rect 227812 285796 227864 285802
rect 227812 285738 227864 285744
rect 227444 284436 227496 284442
rect 227444 284378 227496 284384
rect 227456 284104 227484 284378
rect 227824 284104 227852 285738
rect 228376 284104 228404 288322
rect 232516 287706 232544 345034
rect 232780 297424 232832 297430
rect 232780 297366 232832 297372
rect 232504 287700 232556 287706
rect 232504 287642 232556 287648
rect 231308 287632 231360 287638
rect 231308 287574 231360 287580
rect 230756 287156 230808 287162
rect 230756 287098 230808 287104
rect 229284 287088 229336 287094
rect 229284 287030 229336 287036
rect 228916 286000 228968 286006
rect 228916 285942 228968 285948
rect 228928 284104 228956 285942
rect 229296 284104 229324 287030
rect 229836 285184 229888 285190
rect 229836 285126 229888 285132
rect 229848 284104 229876 285126
rect 230388 284640 230440 284646
rect 230388 284582 230440 284588
rect 230400 284104 230428 284582
rect 230768 284104 230796 287098
rect 231320 284104 231348 287574
rect 232228 287360 232280 287366
rect 232228 287302 232280 287308
rect 231676 284980 231728 284986
rect 231676 284922 231728 284928
rect 231688 284104 231716 284922
rect 232240 284104 232268 287302
rect 232792 284104 232820 297366
rect 233896 289202 233924 656882
rect 233884 289196 233936 289202
rect 233884 289138 233936 289144
rect 234252 285864 234304 285870
rect 234252 285806 234304 285812
rect 233698 284608 233754 284617
rect 233698 284543 233754 284552
rect 233148 284436 233200 284442
rect 233148 284378 233200 284384
rect 233160 284104 233188 284378
rect 233712 284104 233740 284543
rect 234264 284104 234292 285806
rect 234632 284104 234660 700334
rect 234724 312594 234752 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700738 267688 703520
rect 251824 700732 251876 700738
rect 251824 700674 251876 700680
rect 267648 700732 267700 700738
rect 267648 700674 267700 700680
rect 235540 700528 235592 700534
rect 235540 700470 235592 700476
rect 234712 312588 234764 312594
rect 234712 312530 234764 312536
rect 235172 288448 235224 288454
rect 235172 288390 235224 288396
rect 235184 284104 235212 288390
rect 235552 284104 235580 700470
rect 247684 700324 247736 700330
rect 247684 700266 247736 700272
rect 246212 683188 246264 683194
rect 246212 683130 246264 683136
rect 240784 579692 240836 579698
rect 240784 579634 240836 579640
rect 240508 294636 240560 294642
rect 240508 294578 240560 294584
rect 239588 287428 239640 287434
rect 239588 287370 239640 287376
rect 236092 286204 236144 286210
rect 236092 286146 236144 286152
rect 236104 284104 236132 286146
rect 237564 286068 237616 286074
rect 237564 286010 237616 286016
rect 236644 284572 236696 284578
rect 236644 284514 236696 284520
rect 236656 284104 236684 284514
rect 237576 284104 237604 286010
rect 238116 284708 238168 284714
rect 238116 284650 238168 284656
rect 238128 284104 238156 284650
rect 239034 284336 239090 284345
rect 239034 284271 239090 284280
rect 239048 284104 239076 284271
rect 239600 284104 239628 287370
rect 239956 284504 240008 284510
rect 239956 284446 240008 284452
rect 239968 284104 239996 284446
rect 240520 284104 240548 294578
rect 240796 284889 240824 579634
rect 244924 501016 244976 501022
rect 244924 500958 244976 500964
rect 244372 298784 244424 298790
rect 244372 298726 244424 298732
rect 244280 293276 244332 293282
rect 244280 293218 244332 293224
rect 241428 291848 241480 291854
rect 241428 291790 241480 291796
rect 240782 284880 240838 284889
rect 240782 284815 240838 284824
rect 240876 284368 240928 284374
rect 240876 284310 240928 284316
rect 240888 284104 240916 284310
rect 241440 284104 241468 291790
rect 243636 287700 243688 287706
rect 243636 287642 243688 287648
rect 242900 285252 242952 285258
rect 242900 285194 242952 285200
rect 241980 284640 242032 284646
rect 241980 284582 242032 284588
rect 241992 284104 242020 284582
rect 242912 284104 242940 285194
rect 242624 284096 242676 284102
rect 238518 284034 238616 284050
rect 242382 284044 242624 284050
rect 242382 284038 242676 284044
rect 243358 284064 243414 284073
rect 238518 284028 238628 284034
rect 238518 284022 238576 284028
rect 242382 284022 242664 284038
rect 243648 284050 243676 287642
rect 244096 285864 244148 285870
rect 244096 285806 244148 285812
rect 243912 285796 243964 285802
rect 243912 285738 243964 285744
rect 243414 284022 243478 284050
rect 243648 284022 243846 284050
rect 243358 283999 243414 284008
rect 238576 283970 238628 283976
rect 237288 283960 237340 283966
rect 237046 283908 237288 283914
rect 237046 283902 237340 283908
rect 237046 283886 237328 283902
rect 243924 283898 243952 285738
rect 244004 284776 244056 284782
rect 244004 284718 244056 284724
rect 243912 283892 243964 283898
rect 243912 283834 243964 283840
rect 198646 283792 198702 283801
rect 198646 283727 198702 283736
rect 199566 282432 199622 282441
rect 199566 282367 199622 282376
rect 198554 280800 198610 280809
rect 198554 280735 198610 280744
rect 199474 278624 199530 278633
rect 199474 278559 199530 278568
rect 198646 278080 198702 278089
rect 198646 278015 198702 278024
rect 198554 271008 198610 271017
rect 198554 270943 198610 270952
rect 198462 263120 198518 263129
rect 198462 263055 198518 263064
rect 198370 255776 198426 255785
rect 198370 255711 198426 255720
rect 198370 252240 198426 252249
rect 198370 252175 198426 252184
rect 198278 232656 198334 232665
rect 198278 232591 198334 232600
rect 198094 232520 198150 232529
rect 198094 232455 198150 232464
rect 198384 177313 198412 252175
rect 198476 182889 198504 263055
rect 198568 186969 198596 270943
rect 198554 186960 198610 186969
rect 198554 186895 198610 186904
rect 198462 182880 198518 182889
rect 198462 182815 198518 182824
rect 198660 181393 198688 278015
rect 199290 262304 199346 262313
rect 199290 262239 199346 262248
rect 199198 245168 199254 245177
rect 199198 245103 199254 245112
rect 198646 181384 198702 181393
rect 198646 181319 198702 181328
rect 199212 180810 199240 245103
rect 199304 239494 199332 262239
rect 199382 260128 199438 260137
rect 199382 260063 199438 260072
rect 199292 239488 199344 239494
rect 199292 239430 199344 239436
rect 199396 233986 199424 260063
rect 199488 235346 199516 278559
rect 199580 236842 199608 282367
rect 199658 276720 199714 276729
rect 199658 276655 199714 276664
rect 199672 236910 199700 276655
rect 199750 275088 199806 275097
rect 199750 275023 199806 275032
rect 199660 236904 199712 236910
rect 199660 236846 199712 236852
rect 199568 236836 199620 236842
rect 199568 236778 199620 236784
rect 199476 235340 199528 235346
rect 199476 235282 199528 235288
rect 199384 233980 199436 233986
rect 199384 233922 199436 233928
rect 199764 183025 199792 275023
rect 200026 273728 200082 273737
rect 200026 273663 200082 273672
rect 199934 271552 199990 271561
rect 199934 271487 199990 271496
rect 199842 270192 199898 270201
rect 199842 270127 199898 270136
rect 199750 183016 199806 183025
rect 199750 182951 199806 182960
rect 199200 180804 199252 180810
rect 199200 180746 199252 180752
rect 199856 177614 199884 270127
rect 199948 178838 199976 271487
rect 199936 178832 199988 178838
rect 199936 178774 199988 178780
rect 200040 178770 200068 273663
rect 244016 267734 244044 284718
rect 244108 283626 244136 285806
rect 244096 283620 244148 283626
rect 244096 283562 244148 283568
rect 244292 278905 244320 293218
rect 244278 278896 244334 278905
rect 244278 278831 244334 278840
rect 244384 278089 244412 298726
rect 244464 283960 244516 283966
rect 244464 283902 244516 283908
rect 244370 278080 244426 278089
rect 244370 278015 244426 278024
rect 244370 271552 244426 271561
rect 244370 271487 244426 271496
rect 244016 267706 244136 267734
rect 244108 259418 244136 267706
rect 244096 259412 244148 259418
rect 244096 259354 244148 259360
rect 244094 250608 244150 250617
rect 244094 250543 244150 250552
rect 244002 244352 244058 244361
rect 244002 244287 244058 244296
rect 243910 240544 243966 240553
rect 243910 240479 243966 240488
rect 243924 240310 243952 240479
rect 243912 240304 243964 240310
rect 243912 240246 243964 240252
rect 200118 240136 200174 240145
rect 200118 240071 200174 240080
rect 200132 180305 200160 240071
rect 200118 180296 200174 180305
rect 200118 180231 200174 180240
rect 200224 180130 200252 240244
rect 200592 238066 200620 240219
rect 200580 238060 200632 238066
rect 200580 238002 200632 238008
rect 200212 180124 200264 180130
rect 200212 180066 200264 180072
rect 201144 180062 201172 240219
rect 201408 240168 201460 240174
rect 201408 240110 201460 240116
rect 201420 239970 201448 240110
rect 201408 239964 201460 239970
rect 201408 239906 201460 239912
rect 201512 182918 201540 240219
rect 202064 238610 202092 240219
rect 202052 238604 202104 238610
rect 202052 238546 202104 238552
rect 201500 182912 201552 182918
rect 201500 182854 201552 182860
rect 201132 180056 201184 180062
rect 201132 179998 201184 180004
rect 200028 178764 200080 178770
rect 200028 178706 200080 178712
rect 199844 177608 199896 177614
rect 199844 177550 199896 177556
rect 202616 177410 202644 240219
rect 202984 178702 203012 240219
rect 203536 182986 203564 240219
rect 204088 187134 204116 240219
rect 204456 238542 204484 240219
rect 204444 238536 204496 238542
rect 204444 238478 204496 238484
rect 205008 236026 205036 240219
rect 204996 236020 205048 236026
rect 204996 235962 205048 235968
rect 204076 187128 204128 187134
rect 204076 187070 204128 187076
rect 203524 182980 203576 182986
rect 203524 182922 203576 182928
rect 205376 180198 205404 240219
rect 205928 186998 205956 240219
rect 206284 236020 206336 236026
rect 206284 235962 206336 235968
rect 205916 186992 205968 186998
rect 205916 186934 205968 186940
rect 205364 180192 205416 180198
rect 205364 180134 205416 180140
rect 202972 178696 203024 178702
rect 202972 178638 203024 178644
rect 202604 177404 202656 177410
rect 202604 177346 202656 177352
rect 198370 177304 198426 177313
rect 198370 177239 198426 177248
rect 202144 176724 202196 176730
rect 202144 176666 202196 176672
rect 197084 176520 197136 176526
rect 197084 176462 197136 176468
rect 202156 165510 202184 176666
rect 202144 165504 202196 165510
rect 202144 165446 202196 165452
rect 202144 143608 202196 143614
rect 202144 143550 202196 143556
rect 202156 88194 202184 143550
rect 202144 88188 202196 88194
rect 202144 88130 202196 88136
rect 206296 33114 206324 235962
rect 206480 188426 206508 240219
rect 206468 188420 206520 188426
rect 206468 188362 206520 188368
rect 206848 177274 206876 240219
rect 207400 238134 207428 240219
rect 207388 238128 207440 238134
rect 207388 238070 207440 238076
rect 207952 237969 207980 240219
rect 207938 237960 207994 237969
rect 207938 237895 207994 237904
rect 208320 198014 208348 240219
rect 208872 238338 208900 240219
rect 209240 238406 209268 240219
rect 209228 238400 209280 238406
rect 209228 238342 209280 238348
rect 208860 238332 208912 238338
rect 208860 238274 208912 238280
rect 209044 237040 209096 237046
rect 209044 236982 209096 236988
rect 208308 198008 208360 198014
rect 208308 197950 208360 197956
rect 206836 177268 206888 177274
rect 206836 177210 206888 177216
rect 209056 45558 209084 236982
rect 209792 60722 209820 240219
rect 210344 233918 210372 240219
rect 210332 233912 210384 233918
rect 210332 233854 210384 233860
rect 210712 180441 210740 240219
rect 211264 184210 211292 240219
rect 211252 184204 211304 184210
rect 211252 184146 211304 184152
rect 211816 181694 211844 240219
rect 212184 236774 212212 240219
rect 212736 240106 212764 240219
rect 212724 240100 212776 240106
rect 212724 240042 212776 240048
rect 213104 238202 213132 240219
rect 213092 238196 213144 238202
rect 213092 238138 213144 238144
rect 212172 236768 212224 236774
rect 212172 236710 212224 236716
rect 213656 183054 213684 240219
rect 214208 191146 214236 240219
rect 214576 238678 214604 240219
rect 214564 238672 214616 238678
rect 214564 238614 214616 238620
rect 215128 238338 215156 240219
rect 215680 238406 215708 240219
rect 215668 238400 215720 238406
rect 215668 238342 215720 238348
rect 215116 238332 215168 238338
rect 215116 238274 215168 238280
rect 216048 237386 216076 240219
rect 216600 239902 216628 240219
rect 216588 239896 216640 239902
rect 216588 239838 216640 239844
rect 216036 237380 216088 237386
rect 216036 237322 216088 237328
rect 214196 191140 214248 191146
rect 214196 191082 214248 191088
rect 213644 183048 213696 183054
rect 213644 182990 213696 182996
rect 211804 181688 211856 181694
rect 211804 181630 211856 181636
rect 210698 180432 210754 180441
rect 210698 180367 210754 180376
rect 213184 178220 213236 178226
rect 213184 178162 213236 178168
rect 213196 150249 213224 178162
rect 217152 177206 217180 240219
rect 217520 181490 217548 240219
rect 218072 184414 218100 240219
rect 218060 184408 218112 184414
rect 218060 184350 218112 184356
rect 218440 181558 218468 240219
rect 218992 238270 219020 240219
rect 219544 238746 219572 240219
rect 219532 238740 219584 238746
rect 219532 238682 219584 238688
rect 218980 238264 219032 238270
rect 218980 238206 219032 238212
rect 218428 181552 218480 181558
rect 218428 181494 218480 181500
rect 217508 181484 217560 181490
rect 217508 181426 217560 181432
rect 219912 177478 219940 240219
rect 220464 178906 220492 240219
rect 221016 180266 221044 240219
rect 221384 239698 221412 240219
rect 221936 239834 221964 240219
rect 221924 239828 221976 239834
rect 221924 239770 221976 239776
rect 221372 239692 221424 239698
rect 221372 239634 221424 239640
rect 222304 187066 222332 240219
rect 222292 187060 222344 187066
rect 222292 187002 222344 187008
rect 221004 180260 221056 180266
rect 221004 180202 221056 180208
rect 222856 179518 222884 240219
rect 223408 179994 223436 240219
rect 223396 179988 223448 179994
rect 223396 179930 223448 179936
rect 222844 179512 222896 179518
rect 222844 179454 222896 179460
rect 223776 178974 223804 240219
rect 224328 184346 224356 240219
rect 224316 184340 224368 184346
rect 224316 184282 224368 184288
rect 223764 178968 223816 178974
rect 223764 178910 223816 178916
rect 220452 178900 220504 178906
rect 220452 178842 220504 178848
rect 224880 177614 224908 240219
rect 225248 239970 225276 240219
rect 225236 239964 225288 239970
rect 225236 239906 225288 239912
rect 225800 180577 225828 240219
rect 226168 181626 226196 240219
rect 226720 184278 226748 240219
rect 226708 184272 226760 184278
rect 226708 184214 226760 184220
rect 226156 181620 226208 181626
rect 226156 181562 226208 181568
rect 225786 180568 225842 180577
rect 225786 180503 225842 180512
rect 224868 177608 224920 177614
rect 224868 177550 224920 177556
rect 219900 177472 219952 177478
rect 219900 177414 219952 177420
rect 217140 177200 217192 177206
rect 217140 177142 217192 177148
rect 227272 177138 227300 240219
rect 227640 239834 227668 240219
rect 227628 239828 227680 239834
rect 227628 239770 227680 239776
rect 228192 239358 228220 240219
rect 228180 239352 228232 239358
rect 228180 239294 228232 239300
rect 228744 180334 228772 240219
rect 229112 188358 229140 240219
rect 229560 237176 229612 237182
rect 229560 237118 229612 237124
rect 229572 229094 229600 237118
rect 229664 237046 229692 240219
rect 229744 238400 229796 238406
rect 229744 238342 229796 238348
rect 229652 237040 229704 237046
rect 229652 236982 229704 236988
rect 229572 229066 229692 229094
rect 229468 188420 229520 188426
rect 229468 188362 229520 188368
rect 229100 188352 229152 188358
rect 229100 188294 229152 188300
rect 229284 183048 229336 183054
rect 229284 182990 229336 182996
rect 228732 180328 228784 180334
rect 228732 180270 228784 180276
rect 229100 179512 229152 179518
rect 229100 179454 229152 179460
rect 227260 177132 227312 177138
rect 227260 177074 227312 177080
rect 213920 176588 213972 176594
rect 213920 176530 213972 176536
rect 213932 176225 213960 176530
rect 227720 176520 227772 176526
rect 227720 176462 227772 176468
rect 227732 176225 227760 176462
rect 213918 176216 213974 176225
rect 213918 176151 213974 176160
rect 227718 176216 227774 176225
rect 227718 176151 227774 176160
rect 214564 176044 214616 176050
rect 214564 175986 214616 175992
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175137 213960 175170
rect 214012 175160 214064 175166
rect 213918 175128 213974 175137
rect 214012 175102 214064 175108
rect 213918 175063 213974 175072
rect 214024 174729 214052 175102
rect 214010 174720 214066 174729
rect 214010 174655 214066 174664
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173777 213960 173810
rect 214012 173800 214064 173806
rect 213918 173768 213974 173777
rect 214012 173742 214064 173748
rect 213918 173703 213974 173712
rect 214024 173369 214052 173742
rect 214010 173360 214066 173369
rect 214010 173295 214066 173304
rect 214012 172508 214064 172514
rect 214012 172450 214064 172456
rect 213920 172440 213972 172446
rect 213918 172408 213920 172417
rect 213972 172408 213974 172417
rect 213918 172343 213974 172352
rect 214024 172009 214052 172450
rect 214010 172000 214066 172009
rect 214010 171935 214066 171944
rect 213920 171080 213972 171086
rect 213920 171022 213972 171028
rect 213932 170785 213960 171022
rect 213918 170776 213974 170785
rect 213918 170711 213974 170720
rect 214012 169720 214064 169726
rect 213918 169688 213974 169697
rect 214012 169662 214064 169668
rect 213918 169623 213920 169632
rect 213972 169623 213974 169632
rect 213920 169594 213972 169600
rect 214024 169425 214052 169662
rect 214010 169416 214066 169425
rect 214010 169351 214066 169360
rect 213920 168360 213972 168366
rect 213920 168302 213972 168308
rect 213932 168065 213960 168302
rect 214012 168292 214064 168298
rect 214012 168234 214064 168240
rect 213918 168056 213974 168065
rect 213918 167991 213974 168000
rect 214024 167929 214052 168234
rect 214010 167920 214066 167929
rect 214010 167855 214066 167864
rect 213920 167000 213972 167006
rect 213918 166968 213920 166977
rect 213972 166968 213974 166977
rect 213918 166903 213974 166912
rect 214012 166932 214064 166938
rect 214012 166874 214064 166880
rect 214024 166705 214052 166874
rect 214104 166864 214156 166870
rect 214104 166806 214156 166812
rect 214010 166696 214066 166705
rect 214010 166631 214066 166640
rect 214116 166161 214144 166806
rect 214102 166152 214158 166161
rect 214102 166087 214158 166096
rect 214012 165572 214064 165578
rect 214012 165514 214064 165520
rect 213920 165504 213972 165510
rect 213918 165472 213920 165481
rect 213972 165472 213974 165481
rect 213918 165407 213974 165416
rect 214024 164801 214052 165514
rect 214010 164792 214066 164801
rect 214010 164727 214066 164736
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163985 213960 164154
rect 214012 164144 214064 164150
rect 214012 164086 214064 164092
rect 213918 163976 213974 163985
rect 213918 163911 213974 163920
rect 214024 163441 214052 164086
rect 214010 163432 214066 163441
rect 214010 163367 214066 163376
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162625 213960 162794
rect 214012 162784 214064 162790
rect 214012 162726 214064 162732
rect 213918 162616 213974 162625
rect 213918 162551 213974 162560
rect 214024 162081 214052 162726
rect 214010 162072 214066 162081
rect 214010 162007 214066 162016
rect 214576 161474 214604 175986
rect 214656 174548 214708 174554
rect 214656 174490 214708 174496
rect 214668 171057 214696 174490
rect 214654 171048 214710 171057
rect 214654 170983 214710 170992
rect 214748 170400 214800 170406
rect 214748 170342 214800 170348
rect 214484 161446 214604 161474
rect 213920 161424 213972 161430
rect 213918 161392 213920 161401
rect 213972 161392 213974 161401
rect 213918 161327 213974 161336
rect 214012 160064 214064 160070
rect 214012 160006 214064 160012
rect 213920 159996 213972 160002
rect 213920 159938 213972 159944
rect 213932 159905 213960 159938
rect 213918 159896 213974 159905
rect 213918 159831 213974 159840
rect 214024 159497 214052 160006
rect 214010 159488 214066 159497
rect 214010 159423 214066 159432
rect 213920 158704 213972 158710
rect 214484 158681 214512 161446
rect 214760 160857 214788 170342
rect 214746 160848 214802 160857
rect 214746 160783 214802 160792
rect 213920 158646 213972 158652
rect 214470 158672 214526 158681
rect 213932 158137 213960 158646
rect 214470 158607 214526 158616
rect 213918 158128 213974 158137
rect 213918 158063 213974 158072
rect 214012 157344 214064 157350
rect 213918 157312 213974 157321
rect 214012 157286 214064 157292
rect 213918 157247 213920 157256
rect 213972 157247 213974 157256
rect 213920 157218 213972 157224
rect 214024 156913 214052 157286
rect 214010 156904 214066 156913
rect 214010 156839 214066 156848
rect 213918 155952 213974 155961
rect 213918 155887 213920 155896
rect 213972 155887 213974 155896
rect 213920 155858 213972 155864
rect 214012 155848 214064 155854
rect 214012 155790 214064 155796
rect 214024 155417 214052 155790
rect 214010 155408 214066 155417
rect 214010 155343 214066 155352
rect 214010 153912 214066 153921
rect 214010 153847 214066 153856
rect 213918 153504 213974 153513
rect 213918 153439 213974 153448
rect 213932 153270 213960 153439
rect 214024 153338 214052 153847
rect 214012 153332 214064 153338
rect 214012 153274 214064 153280
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 213918 152688 213974 152697
rect 213918 152623 213974 152632
rect 213932 151842 213960 152623
rect 214746 152144 214802 152153
rect 214746 152079 214802 152088
rect 213920 151836 213972 151842
rect 214760 151814 214788 152079
rect 214838 152008 214894 152017
rect 214838 151943 214894 151952
rect 213920 151778 213972 151784
rect 214576 151786 214788 151814
rect 214010 150920 214066 150929
rect 214010 150855 214066 150864
rect 214024 150482 214052 150855
rect 214012 150476 214064 150482
rect 214012 150418 214064 150424
rect 213920 150408 213972 150414
rect 213920 150350 213972 150356
rect 213182 150240 213238 150249
rect 213182 150175 213238 150184
rect 213932 149569 213960 150350
rect 213918 149560 213974 149569
rect 213918 149495 213974 149504
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148753 213960 148990
rect 213918 148744 213974 148753
rect 213918 148679 213974 148688
rect 213918 148064 213974 148073
rect 213918 147999 213974 148008
rect 213932 147694 213960 147999
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 214010 146704 214066 146713
rect 214010 146639 214066 146648
rect 213918 146432 213974 146441
rect 213918 146367 213920 146376
rect 213972 146367 213974 146376
rect 213920 146338 213972 146344
rect 214024 146334 214052 146639
rect 214012 146328 214064 146334
rect 214012 146270 214064 146276
rect 214010 145344 214066 145353
rect 214010 145279 214066 145288
rect 214024 145042 214052 145279
rect 214012 145036 214064 145042
rect 214012 144978 214064 144984
rect 213920 144968 213972 144974
rect 213918 144936 213920 144945
rect 213972 144936 213974 144945
rect 213918 144871 213974 144880
rect 214470 143984 214526 143993
rect 214470 143919 214526 143928
rect 213920 143608 213972 143614
rect 213918 143576 213920 143585
rect 213972 143576 213974 143585
rect 213918 143511 213974 143520
rect 214010 142760 214066 142769
rect 214010 142695 214066 142704
rect 213918 142352 213974 142361
rect 213918 142287 213974 142296
rect 213932 142254 213960 142287
rect 213920 142248 213972 142254
rect 213920 142190 213972 142196
rect 214024 142186 214052 142695
rect 214012 142180 214064 142186
rect 214012 142122 214064 142128
rect 214010 141400 214066 141409
rect 214010 141335 214066 141344
rect 213918 140992 213974 141001
rect 213918 140927 213974 140936
rect 213932 140894 213960 140927
rect 213920 140888 213972 140894
rect 213920 140830 213972 140836
rect 214024 140826 214052 141335
rect 214012 140820 214064 140826
rect 214012 140762 214064 140768
rect 214010 140040 214066 140049
rect 214010 139975 214066 139984
rect 213918 139632 213974 139641
rect 213918 139567 213974 139576
rect 213932 139534 213960 139567
rect 213920 139528 213972 139534
rect 213920 139470 213972 139476
rect 214024 139466 214052 139975
rect 214012 139460 214064 139466
rect 214012 139402 214064 139408
rect 213918 136776 213974 136785
rect 213918 136711 213974 136720
rect 213932 136678 213960 136711
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 214010 136096 214066 136105
rect 214010 136031 214066 136040
rect 214024 135454 214052 136031
rect 214102 135688 214158 135697
rect 214102 135623 214158 135632
rect 214012 135448 214064 135454
rect 213918 135416 213974 135425
rect 214012 135390 214064 135396
rect 213918 135351 213920 135360
rect 213972 135351 213974 135360
rect 213920 135322 213972 135328
rect 214116 135318 214144 135623
rect 214104 135312 214156 135318
rect 214104 135254 214156 135260
rect 213918 134328 213974 134337
rect 213918 134263 213974 134272
rect 213932 133958 213960 134263
rect 214484 133958 214512 143919
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 214472 133952 214524 133958
rect 214472 133894 214524 133900
rect 214576 133346 214604 151786
rect 214852 151094 214880 151943
rect 214840 151088 214892 151094
rect 214840 151030 214892 151036
rect 214746 150784 214802 150793
rect 214746 150719 214802 150728
rect 214760 137290 214788 150719
rect 229112 150657 229140 179454
rect 229192 177608 229244 177614
rect 229192 177550 229244 177556
rect 229204 169561 229232 177550
rect 229190 169552 229246 169561
rect 229190 169487 229246 169496
rect 229296 154329 229324 182990
rect 229376 180532 229428 180538
rect 229376 180474 229428 180480
rect 229388 174321 229416 180474
rect 229374 174312 229430 174321
rect 229374 174247 229430 174256
rect 229376 174208 229428 174214
rect 229376 174150 229428 174156
rect 229282 154320 229338 154329
rect 229282 154255 229338 154264
rect 229388 153377 229416 174150
rect 229480 161537 229508 188362
rect 229560 178900 229612 178906
rect 229560 178842 229612 178848
rect 229572 169017 229600 178842
rect 229558 169008 229614 169017
rect 229558 168943 229614 168952
rect 229466 161528 229522 161537
rect 229466 161463 229522 161472
rect 229374 153368 229430 153377
rect 229374 153303 229430 153312
rect 229098 150648 229154 150657
rect 229098 150583 229154 150592
rect 214838 138136 214894 138145
rect 214838 138071 214894 138080
rect 214748 137284 214800 137290
rect 214748 137226 214800 137232
rect 214656 133952 214708 133958
rect 214656 133894 214708 133900
rect 214564 133340 214616 133346
rect 214564 133282 214616 133288
rect 214564 133136 214616 133142
rect 214564 133078 214616 133084
rect 214010 132832 214066 132841
rect 214010 132767 214066 132776
rect 213920 132592 213972 132598
rect 213918 132560 213920 132569
rect 213972 132560 213974 132569
rect 214024 132530 214052 132767
rect 213918 132495 213974 132504
rect 214012 132524 214064 132530
rect 214012 132466 214064 132472
rect 214010 131472 214066 131481
rect 214010 131407 214066 131416
rect 214024 131238 214052 131407
rect 214012 131232 214064 131238
rect 213918 131200 213974 131209
rect 214012 131174 214064 131180
rect 213918 131135 213920 131144
rect 213972 131135 213974 131144
rect 213920 131106 213972 131112
rect 214010 130112 214066 130121
rect 214010 130047 214066 130056
rect 213920 129872 213972 129878
rect 213918 129840 213920 129849
rect 213972 129840 213974 129849
rect 214024 129810 214052 130047
rect 213918 129775 213974 129784
rect 214012 129804 214064 129810
rect 214012 129746 214064 129752
rect 214010 128888 214066 128897
rect 214010 128823 214066 128832
rect 213918 128480 213974 128489
rect 213918 128415 213920 128424
rect 213972 128415 213974 128424
rect 213920 128386 213972 128392
rect 214024 128382 214052 128823
rect 214012 128376 214064 128382
rect 214012 128318 214064 128324
rect 214010 127528 214066 127537
rect 214010 127463 214066 127472
rect 213918 127120 213974 127129
rect 213918 127055 213920 127064
rect 213972 127055 213974 127064
rect 213920 127026 213972 127032
rect 214024 127022 214052 127463
rect 214012 127016 214064 127022
rect 214012 126958 214064 126964
rect 214010 126168 214066 126177
rect 214010 126103 214066 126112
rect 213918 125760 213974 125769
rect 213918 125695 213920 125704
rect 213972 125695 213974 125704
rect 213920 125666 213972 125672
rect 214024 125662 214052 126103
rect 214012 125656 214064 125662
rect 214012 125598 214064 125604
rect 214010 124808 214066 124817
rect 214010 124743 214066 124752
rect 214024 124302 214052 124743
rect 214012 124296 214064 124302
rect 213918 124264 213974 124273
rect 214012 124238 214064 124244
rect 213918 124199 213920 124208
rect 213972 124199 213974 124208
rect 213920 124170 213972 124176
rect 214010 123584 214066 123593
rect 214010 123519 214066 123528
rect 213918 123176 213974 123185
rect 213918 123111 213974 123120
rect 213932 122942 213960 123111
rect 213920 122936 213972 122942
rect 213920 122878 213972 122884
rect 214024 122874 214052 123519
rect 214012 122868 214064 122874
rect 214012 122810 214064 122816
rect 214010 122224 214066 122233
rect 214010 122159 214066 122168
rect 213918 121816 213974 121825
rect 213918 121751 213974 121760
rect 213932 121582 213960 121751
rect 213920 121576 213972 121582
rect 213920 121518 213972 121524
rect 214024 121514 214052 122159
rect 214012 121508 214064 121514
rect 214012 121450 214064 121456
rect 214010 120864 214066 120873
rect 214010 120799 214066 120808
rect 213918 120456 213974 120465
rect 213918 120391 213974 120400
rect 213932 120222 213960 120391
rect 213920 120216 213972 120222
rect 213920 120158 213972 120164
rect 214024 120154 214052 120799
rect 214012 120148 214064 120154
rect 214012 120090 214064 120096
rect 213918 119640 213974 119649
rect 213918 119575 213974 119584
rect 213932 118862 213960 119575
rect 214010 118960 214066 118969
rect 214010 118895 214066 118904
rect 213920 118856 213972 118862
rect 213182 118824 213238 118833
rect 213920 118798 213972 118804
rect 214024 118794 214052 118895
rect 213182 118759 213238 118768
rect 214012 118788 214064 118794
rect 213196 91050 213224 118759
rect 214012 118730 214064 118736
rect 213920 117360 213972 117366
rect 213918 117328 213920 117337
rect 213972 117328 213974 117337
rect 213918 117263 213974 117272
rect 214010 116240 214066 116249
rect 214010 116175 214066 116184
rect 213920 116068 213972 116074
rect 213920 116010 213972 116016
rect 213932 115977 213960 116010
rect 214024 116006 214052 116175
rect 214012 116000 214064 116006
rect 213918 115968 213974 115977
rect 214012 115942 214064 115948
rect 213918 115903 213974 115912
rect 214010 115016 214066 115025
rect 214010 114951 214066 114960
rect 214024 114646 214052 114951
rect 214012 114640 214064 114646
rect 213918 114608 213974 114617
rect 214012 114582 214064 114588
rect 213918 114543 213920 114552
rect 213972 114543 213974 114552
rect 213920 114514 213972 114520
rect 214010 113656 214066 113665
rect 214010 113591 214066 113600
rect 214024 113286 214052 113591
rect 214012 113280 214064 113286
rect 213918 113248 213974 113257
rect 214012 113222 214064 113228
rect 213918 113183 213920 113192
rect 213972 113183 213974 113192
rect 213920 113154 213972 113160
rect 214010 112296 214066 112305
rect 214010 112231 214066 112240
rect 213920 111920 213972 111926
rect 213918 111888 213920 111897
rect 213972 111888 213974 111897
rect 214024 111858 214052 112231
rect 213918 111823 213974 111832
rect 214012 111852 214064 111858
rect 214012 111794 214064 111800
rect 213918 110528 213974 110537
rect 213918 110463 213920 110472
rect 213972 110463 213974 110472
rect 213920 110434 213972 110440
rect 214010 109712 214066 109721
rect 214010 109647 214066 109656
rect 213918 109168 213974 109177
rect 213918 109103 213920 109112
rect 213972 109103 213974 109112
rect 213920 109074 213972 109080
rect 214024 109070 214052 109647
rect 214012 109064 214064 109070
rect 214012 109006 214064 109012
rect 213918 108352 213974 108361
rect 213918 108287 213974 108296
rect 213932 107710 213960 108287
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 214010 106992 214066 107001
rect 214010 106927 214066 106936
rect 213918 106584 213974 106593
rect 213918 106519 213974 106528
rect 213932 106350 213960 106519
rect 214024 106418 214052 106927
rect 214012 106412 214064 106418
rect 214012 106354 214064 106360
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 214102 105768 214158 105777
rect 214102 105703 214158 105712
rect 214010 105360 214066 105369
rect 214010 105295 214066 105304
rect 213918 105088 213974 105097
rect 213918 105023 213920 105032
rect 213972 105023 213974 105032
rect 213920 104994 213972 105000
rect 214024 104990 214052 105295
rect 214012 104984 214064 104990
rect 214012 104926 214064 104932
rect 214116 104922 214144 105703
rect 214104 104916 214156 104922
rect 214104 104858 214156 104864
rect 213918 103728 213974 103737
rect 213918 103663 213974 103672
rect 213932 103562 213960 103663
rect 213920 103556 213972 103562
rect 213920 103498 213972 103504
rect 214010 102640 214066 102649
rect 214010 102575 214066 102584
rect 213918 102368 213974 102377
rect 213918 102303 213974 102312
rect 213932 102202 213960 102303
rect 214024 102270 214052 102575
rect 214012 102264 214064 102270
rect 214012 102206 214064 102212
rect 213920 102196 213972 102202
rect 213920 102138 213972 102144
rect 214288 101108 214340 101114
rect 214288 101050 214340 101056
rect 214194 99784 214250 99793
rect 214194 99719 214250 99728
rect 214102 99512 214158 99521
rect 214102 99447 214158 99456
rect 213918 98424 213974 98433
rect 213918 98359 213974 98368
rect 213932 98054 213960 98359
rect 213920 98048 213972 98054
rect 213920 97990 213972 97996
rect 214010 98016 214066 98025
rect 214010 97951 214066 97960
rect 213918 97064 213974 97073
rect 213918 96999 213974 97008
rect 213932 96694 213960 96999
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 214024 96082 214052 97951
rect 214116 96150 214144 99447
rect 214104 96144 214156 96150
rect 214104 96086 214156 96092
rect 214012 96076 214064 96082
rect 214012 96018 214064 96024
rect 214208 95946 214236 99719
rect 214196 95940 214248 95946
rect 214196 95882 214248 95888
rect 213918 95840 213974 95849
rect 213918 95775 213974 95784
rect 213932 95266 213960 95775
rect 213920 95260 213972 95266
rect 213920 95202 213972 95208
rect 214300 91526 214328 101050
rect 214378 100872 214434 100881
rect 214378 100807 214434 100816
rect 214392 94586 214420 100807
rect 214380 94580 214432 94586
rect 214380 94522 214432 94528
rect 214576 93838 214604 133078
rect 214668 96014 214696 133894
rect 214852 122834 214880 138071
rect 229664 136921 229692 229066
rect 229756 170134 229784 238342
rect 230216 236706 230244 240219
rect 230584 237182 230612 240219
rect 231144 239986 231172 240219
rect 231144 239958 231256 239986
rect 231228 238754 231256 239958
rect 231228 238726 231348 238754
rect 230572 237176 230624 237182
rect 230572 237118 230624 237124
rect 230756 236904 230808 236910
rect 230756 236846 230808 236852
rect 230204 236700 230256 236706
rect 230204 236642 230256 236648
rect 230664 235340 230716 235346
rect 230664 235282 230716 235288
rect 230572 233980 230624 233986
rect 230572 233922 230624 233928
rect 229836 180056 229888 180062
rect 229836 179998 229888 180004
rect 229848 174214 229876 179998
rect 230480 177540 230532 177546
rect 230480 177482 230532 177488
rect 229836 174208 229888 174214
rect 229836 174150 229888 174156
rect 229744 170128 229796 170134
rect 229744 170070 229796 170076
rect 230492 158681 230520 177482
rect 230478 158672 230534 158681
rect 230478 158607 230534 158616
rect 230584 156618 230612 233922
rect 230676 173777 230704 235282
rect 230768 176050 230796 236846
rect 231216 236836 231268 236842
rect 231216 236778 231268 236784
rect 230940 180804 230992 180810
rect 230940 180746 230992 180752
rect 230848 178832 230900 178838
rect 230848 178774 230900 178780
rect 230756 176044 230808 176050
rect 230756 175986 230808 175992
rect 230756 175092 230808 175098
rect 230756 175034 230808 175040
rect 230768 174729 230796 175034
rect 230754 174720 230810 174729
rect 230754 174655 230810 174664
rect 230662 173768 230718 173777
rect 230662 173703 230718 173712
rect 230756 170128 230808 170134
rect 230756 170070 230808 170076
rect 230664 159792 230716 159798
rect 230664 159734 230716 159740
rect 230676 159633 230704 159734
rect 230662 159624 230718 159633
rect 230662 159559 230718 159568
rect 230584 156590 230704 156618
rect 230572 155916 230624 155922
rect 230572 155858 230624 155864
rect 230480 155848 230532 155854
rect 230478 155816 230480 155825
rect 230532 155816 230534 155825
rect 230478 155751 230534 155760
rect 230480 155304 230532 155310
rect 230478 155272 230480 155281
rect 230532 155272 230534 155281
rect 230478 155207 230534 155216
rect 230584 154873 230612 155858
rect 230570 154864 230626 154873
rect 230570 154799 230626 154808
rect 230676 153762 230704 156590
rect 230768 153882 230796 170070
rect 230860 153921 230888 178774
rect 230846 153912 230902 153921
rect 230756 153876 230808 153882
rect 230846 153847 230902 153856
rect 230756 153818 230808 153824
rect 230676 153734 230888 153762
rect 230756 153672 230808 153678
rect 230756 153614 230808 153620
rect 230768 151065 230796 153614
rect 230754 151056 230810 151065
rect 230754 150991 230810 151000
rect 230756 150340 230808 150346
rect 230756 150282 230808 150288
rect 230768 149705 230796 150282
rect 230754 149696 230810 149705
rect 230754 149631 230810 149640
rect 230572 147144 230624 147150
rect 230572 147086 230624 147092
rect 230584 146849 230612 147086
rect 230570 146840 230626 146849
rect 230570 146775 230626 146784
rect 230860 145897 230888 153734
rect 230846 145888 230902 145897
rect 230846 145823 230902 145832
rect 230952 138281 230980 180746
rect 231032 178764 231084 178770
rect 231032 178706 231084 178712
rect 231044 170746 231072 178706
rect 231124 173868 231176 173874
rect 231124 173810 231176 173816
rect 231136 173369 231164 173810
rect 231122 173360 231178 173369
rect 231122 173295 231178 173304
rect 231032 170740 231084 170746
rect 231032 170682 231084 170688
rect 231228 170626 231256 236778
rect 231320 229094 231348 238726
rect 231504 238474 231532 240219
rect 231952 239556 232004 239562
rect 231952 239498 232004 239504
rect 231492 238468 231544 238474
rect 231492 238410 231544 238416
rect 231860 237176 231912 237182
rect 231860 237118 231912 237124
rect 231320 229066 231624 229094
rect 231398 177712 231454 177721
rect 231398 177647 231454 177656
rect 231308 176044 231360 176050
rect 231308 175986 231360 175992
rect 231044 170598 231256 170626
rect 231044 161945 231072 170598
rect 231124 170536 231176 170542
rect 231216 170536 231268 170542
rect 231124 170478 231176 170484
rect 231214 170504 231216 170513
rect 231268 170504 231270 170513
rect 231030 161936 231086 161945
rect 231030 161871 231086 161880
rect 231032 158364 231084 158370
rect 231032 158306 231084 158312
rect 231044 157729 231072 158306
rect 231030 157720 231086 157729
rect 231030 157655 231086 157664
rect 231136 156233 231164 170478
rect 231214 170439 231270 170448
rect 231320 169969 231348 175986
rect 231412 171358 231440 177647
rect 231492 173800 231544 173806
rect 231492 173742 231544 173748
rect 231504 172825 231532 173742
rect 231490 172816 231546 172825
rect 231490 172751 231546 172760
rect 231492 172440 231544 172446
rect 231492 172382 231544 172388
rect 231504 171873 231532 172382
rect 231490 171864 231546 171873
rect 231490 171799 231546 171808
rect 231400 171352 231452 171358
rect 231400 171294 231452 171300
rect 231306 169960 231362 169969
rect 231306 169895 231362 169904
rect 231492 168292 231544 168298
rect 231492 168234 231544 168240
rect 231400 168224 231452 168230
rect 231400 168166 231452 168172
rect 231412 167113 231440 168166
rect 231504 167657 231532 168234
rect 231490 167648 231546 167657
rect 231490 167583 231546 167592
rect 231398 167104 231454 167113
rect 231398 167039 231454 167048
rect 231308 166728 231360 166734
rect 231306 166696 231308 166705
rect 231360 166696 231362 166705
rect 231306 166631 231362 166640
rect 231400 164824 231452 164830
rect 231398 164792 231400 164801
rect 231452 164792 231454 164801
rect 231398 164727 231454 164736
rect 231492 164212 231544 164218
rect 231492 164154 231544 164160
rect 231400 163872 231452 163878
rect 231398 163840 231400 163849
rect 231452 163840 231454 163849
rect 231398 163775 231454 163784
rect 231504 162897 231532 164154
rect 231490 162888 231546 162897
rect 231490 162823 231546 162832
rect 231216 159996 231268 160002
rect 231216 159938 231268 159944
rect 231228 159089 231256 159938
rect 231214 159080 231270 159089
rect 231214 159015 231270 159024
rect 231492 157276 231544 157282
rect 231492 157218 231544 157224
rect 231504 156777 231532 157218
rect 231490 156768 231546 156777
rect 231490 156703 231546 156712
rect 231122 156224 231178 156233
rect 231122 156159 231178 156168
rect 231124 153128 231176 153134
rect 231124 153070 231176 153076
rect 231136 152561 231164 153070
rect 231308 153060 231360 153066
rect 231308 153002 231360 153008
rect 231122 152552 231178 152561
rect 231122 152487 231178 152496
rect 231320 152017 231348 153002
rect 231306 152008 231362 152017
rect 231306 151943 231362 151952
rect 231596 151609 231624 229066
rect 231766 175264 231822 175273
rect 231766 175199 231822 175208
rect 231780 175166 231808 175199
rect 231768 175160 231820 175166
rect 231768 175102 231820 175108
rect 231768 172508 231820 172514
rect 231768 172450 231820 172456
rect 231780 172417 231808 172450
rect 231766 172408 231822 172417
rect 231676 172372 231728 172378
rect 231766 172343 231822 172352
rect 231676 172314 231728 172320
rect 231688 171465 231716 172314
rect 231674 171456 231730 171465
rect 231674 171391 231730 171400
rect 231676 171352 231728 171358
rect 231676 171294 231728 171300
rect 231582 151600 231638 151609
rect 231582 151535 231638 151544
rect 231216 148776 231268 148782
rect 231214 148744 231216 148753
rect 231268 148744 231270 148753
rect 231214 148679 231270 148688
rect 231688 146305 231716 171294
rect 231768 171080 231820 171086
rect 231768 171022 231820 171028
rect 231780 170921 231808 171022
rect 231766 170912 231822 170921
rect 231766 170847 231822 170856
rect 231768 169720 231820 169726
rect 231768 169662 231820 169668
rect 231780 168609 231808 169662
rect 231766 168600 231822 168609
rect 231766 168535 231822 168544
rect 231768 168360 231820 168366
rect 231768 168302 231820 168308
rect 231780 168065 231808 168302
rect 231766 168056 231822 168065
rect 231766 167991 231822 168000
rect 231768 166660 231820 166666
rect 231768 166602 231820 166608
rect 231780 166161 231808 166602
rect 231766 166152 231822 166161
rect 231766 166087 231822 166096
rect 231768 165776 231820 165782
rect 231766 165744 231768 165753
rect 231820 165744 231822 165753
rect 231766 165679 231822 165688
rect 231768 165572 231820 165578
rect 231768 165514 231820 165520
rect 231780 165209 231808 165514
rect 231766 165200 231822 165209
rect 231766 165135 231822 165144
rect 231768 164960 231820 164966
rect 231768 164902 231820 164908
rect 231780 164393 231808 164902
rect 231766 164384 231822 164393
rect 231766 164319 231822 164328
rect 231768 163464 231820 163470
rect 231766 163432 231768 163441
rect 231820 163432 231822 163441
rect 231766 163367 231822 163376
rect 231768 161424 231820 161430
rect 231768 161366 231820 161372
rect 231780 160993 231808 161366
rect 231766 160984 231822 160993
rect 231766 160919 231822 160928
rect 231768 160608 231820 160614
rect 231766 160576 231768 160585
rect 231820 160576 231822 160585
rect 231766 160511 231822 160520
rect 231766 160032 231822 160041
rect 231766 159967 231822 159976
rect 231780 159934 231808 159967
rect 231768 159928 231820 159934
rect 231768 159870 231820 159876
rect 231768 158704 231820 158710
rect 231768 158646 231820 158652
rect 231780 158137 231808 158646
rect 231766 158128 231822 158137
rect 231766 158063 231822 158072
rect 231768 157344 231820 157350
rect 231768 157286 231820 157292
rect 231780 157185 231808 157286
rect 231766 157176 231822 157185
rect 231766 157111 231822 157120
rect 231768 153196 231820 153202
rect 231768 153138 231820 153144
rect 231780 152969 231808 153138
rect 231766 152960 231822 152969
rect 231766 152895 231822 152904
rect 231768 150408 231820 150414
rect 231768 150350 231820 150356
rect 231780 150113 231808 150350
rect 231766 150104 231822 150113
rect 231766 150039 231822 150048
rect 231768 149048 231820 149054
rect 231768 148990 231820 148996
rect 231780 148209 231808 148990
rect 231766 148200 231822 148209
rect 231766 148135 231822 148144
rect 231768 147620 231820 147626
rect 231768 147562 231820 147568
rect 231780 147257 231808 147562
rect 231766 147248 231822 147257
rect 231766 147183 231822 147192
rect 231674 146296 231730 146305
rect 231308 146260 231360 146266
rect 231674 146231 231730 146240
rect 231308 146202 231360 146208
rect 231320 145353 231348 146202
rect 231676 145648 231728 145654
rect 231676 145590 231728 145596
rect 231306 145344 231362 145353
rect 231306 145279 231362 145288
rect 231124 145036 231176 145042
rect 231124 144978 231176 144984
rect 231136 144945 231164 144978
rect 231122 144936 231178 144945
rect 231122 144871 231178 144880
rect 231308 144900 231360 144906
rect 231308 144842 231360 144848
rect 231320 144401 231348 144842
rect 231306 144392 231362 144401
rect 231306 144327 231362 144336
rect 231308 143540 231360 143546
rect 231308 143482 231360 143488
rect 231320 143041 231348 143482
rect 231306 143032 231362 143041
rect 231306 142967 231362 142976
rect 231688 142497 231716 145590
rect 231768 144832 231820 144838
rect 231768 144774 231820 144780
rect 231780 143993 231808 144774
rect 231766 143984 231822 143993
rect 231766 143919 231822 143928
rect 231768 143472 231820 143478
rect 231766 143440 231768 143449
rect 231820 143440 231822 143449
rect 231766 143375 231822 143384
rect 231674 142488 231730 142497
rect 231674 142423 231730 142432
rect 231768 142112 231820 142118
rect 231766 142080 231768 142089
rect 231820 142080 231822 142089
rect 231400 142044 231452 142050
rect 231766 142015 231822 142024
rect 231400 141986 231452 141992
rect 231412 141137 231440 141986
rect 231768 141704 231820 141710
rect 231766 141672 231768 141681
rect 231820 141672 231822 141681
rect 231766 141607 231822 141616
rect 231398 141128 231454 141137
rect 231398 141063 231454 141072
rect 231768 140752 231820 140758
rect 231768 140694 231820 140700
rect 231216 140684 231268 140690
rect 231216 140626 231268 140632
rect 231228 140185 231256 140626
rect 231214 140176 231270 140185
rect 231214 140111 231270 140120
rect 231216 140072 231268 140078
rect 231216 140014 231268 140020
rect 231124 138780 231176 138786
rect 231124 138722 231176 138728
rect 230938 138272 230994 138281
rect 230938 138207 230994 138216
rect 229650 136912 229706 136921
rect 229650 136847 229706 136856
rect 229928 136672 229980 136678
rect 229928 136614 229980 136620
rect 215114 134192 215170 134201
rect 215114 134127 215170 134136
rect 214760 122806 214880 122834
rect 214656 96008 214708 96014
rect 214656 95950 214708 95956
rect 214564 93832 214616 93838
rect 214564 93774 214616 93780
rect 214760 93129 214788 122806
rect 214838 117600 214894 117609
rect 214838 117535 214894 117544
rect 214852 100994 214880 117535
rect 215128 112470 215156 134127
rect 229836 133952 229888 133958
rect 229836 133894 229888 133900
rect 229744 117360 229796 117366
rect 229744 117302 229796 117308
rect 215116 112464 215168 112470
rect 215116 112406 215168 112412
rect 215022 110936 215078 110945
rect 215022 110871 215078 110880
rect 214930 107672 214986 107681
rect 214930 107607 214986 107616
rect 214944 101114 214972 107607
rect 214932 101108 214984 101114
rect 214932 101050 214984 101056
rect 214852 100966 214972 100994
rect 214944 93158 214972 100966
rect 215036 94518 215064 110871
rect 228364 95260 228416 95266
rect 228364 95202 228416 95208
rect 215024 94512 215076 94518
rect 215024 94454 215076 94460
rect 214932 93152 214984 93158
rect 214746 93120 214802 93129
rect 214932 93094 214984 93100
rect 214746 93055 214802 93064
rect 214288 91520 214340 91526
rect 214288 91462 214340 91468
rect 213184 91044 213236 91050
rect 213184 90986 213236 90992
rect 209780 60716 209832 60722
rect 209780 60658 209832 60664
rect 209044 45552 209096 45558
rect 209044 45494 209096 45500
rect 206284 33108 206336 33114
rect 206284 33050 206336 33056
rect 196624 20664 196676 20670
rect 196624 20606 196676 20612
rect 228376 17270 228404 95202
rect 228364 17264 228416 17270
rect 228364 17206 228416 17212
rect 180064 3664 180116 3670
rect 180064 3606 180116 3612
rect 169024 3596 169076 3602
rect 169024 3538 169076 3544
rect 229756 3534 229784 117302
rect 229848 51814 229876 133894
rect 229940 68406 229968 136614
rect 230664 133748 230716 133754
rect 230664 133690 230716 133696
rect 230676 133521 230704 133690
rect 230662 133512 230718 133521
rect 230662 133447 230718 133456
rect 230940 131096 230992 131102
rect 230940 131038 230992 131044
rect 230952 129849 230980 131038
rect 231032 130824 231084 130830
rect 231032 130766 231084 130772
rect 231044 130665 231072 130766
rect 231030 130656 231086 130665
rect 231030 130591 231086 130600
rect 230938 129840 230994 129849
rect 230938 129775 230994 129784
rect 230848 126268 230900 126274
rect 230848 126210 230900 126216
rect 230664 124976 230716 124982
rect 230664 124918 230716 124924
rect 230676 122834 230704 124918
rect 230756 124908 230808 124914
rect 230756 124850 230808 124856
rect 230768 123185 230796 124850
rect 230860 124137 230888 126210
rect 231136 124545 231164 138722
rect 231122 124536 231178 124545
rect 231122 124471 231178 124480
rect 230846 124128 230902 124137
rect 230846 124063 230902 124072
rect 230754 123176 230810 123185
rect 230754 123111 230810 123120
rect 230676 122806 230796 122834
rect 230572 120012 230624 120018
rect 230572 119954 230624 119960
rect 230584 118969 230612 119954
rect 230570 118960 230626 118969
rect 230570 118895 230626 118904
rect 230572 118448 230624 118454
rect 230570 118416 230572 118425
rect 230624 118416 230626 118425
rect 230570 118351 230626 118360
rect 230768 117473 230796 122806
rect 231124 122664 231176 122670
rect 231124 122606 231176 122612
rect 231136 122233 231164 122606
rect 231122 122224 231178 122233
rect 231122 122159 231178 122168
rect 231032 120760 231084 120766
rect 231032 120702 231084 120708
rect 230754 117464 230810 117473
rect 230754 117399 230810 117408
rect 230940 115864 230992 115870
rect 230940 115806 230992 115812
rect 230952 115161 230980 115806
rect 230938 115152 230994 115161
rect 230938 115087 230994 115096
rect 231044 114209 231072 120702
rect 231124 116680 231176 116686
rect 231124 116622 231176 116628
rect 231030 114200 231086 114209
rect 231030 114135 231086 114144
rect 230940 110220 230992 110226
rect 230940 110162 230992 110168
rect 230952 109857 230980 110162
rect 230938 109848 230994 109857
rect 230938 109783 230994 109792
rect 231032 108588 231084 108594
rect 231032 108530 231084 108536
rect 231044 107953 231072 108530
rect 231030 107944 231086 107953
rect 231030 107879 231086 107888
rect 230940 106956 230992 106962
rect 230940 106898 230992 106904
rect 230756 106072 230808 106078
rect 230756 106014 230808 106020
rect 230768 105641 230796 106014
rect 230754 105632 230810 105641
rect 230572 105596 230624 105602
rect 230754 105567 230810 105576
rect 230572 105538 230624 105544
rect 230584 102785 230612 105538
rect 230756 104712 230808 104718
rect 230754 104680 230756 104689
rect 230808 104680 230810 104689
rect 230754 104615 230810 104624
rect 230952 104281 230980 106898
rect 230938 104272 230994 104281
rect 230938 104207 230994 104216
rect 230664 104168 230716 104174
rect 230664 104110 230716 104116
rect 230570 102776 230626 102785
rect 230570 102711 230626 102720
rect 230676 101833 230704 104110
rect 230662 101824 230718 101833
rect 230662 101759 230718 101768
rect 231136 100881 231164 116622
rect 231228 113174 231256 140014
rect 231780 139777 231808 140694
rect 231766 139768 231822 139777
rect 231766 139703 231822 139712
rect 231766 139224 231822 139233
rect 231872 139210 231900 237118
rect 231964 147801 231992 239498
rect 232056 177614 232084 240219
rect 232608 239630 232636 240219
rect 232976 240038 233004 240219
rect 232964 240032 233016 240038
rect 232964 239974 233016 239980
rect 233528 239766 233556 240219
rect 233516 239760 233568 239766
rect 233516 239702 233568 239708
rect 232596 239624 232648 239630
rect 232596 239566 232648 239572
rect 233148 239420 233200 239426
rect 233148 239362 233200 239368
rect 233160 238406 233188 239362
rect 233148 238400 233200 238406
rect 233148 238342 233200 238348
rect 233424 187128 233476 187134
rect 233424 187070 233476 187076
rect 232136 181688 232188 181694
rect 232136 181630 232188 181636
rect 232044 177608 232096 177614
rect 232044 177550 232096 177556
rect 232148 155310 232176 181630
rect 232320 180600 232372 180606
rect 232320 180542 232372 180548
rect 232228 179988 232280 179994
rect 232228 179930 232280 179936
rect 232240 155854 232268 179930
rect 232332 159798 232360 180542
rect 232412 178968 232464 178974
rect 232412 178910 232464 178916
rect 232320 159792 232372 159798
rect 232320 159734 232372 159740
rect 232228 155848 232280 155854
rect 232228 155790 232280 155796
rect 232136 155304 232188 155310
rect 232136 155246 232188 155252
rect 231950 147792 232006 147801
rect 231950 147727 232006 147736
rect 232424 147150 232452 178910
rect 233240 177676 233292 177682
rect 233240 177618 233292 177624
rect 233252 170542 233280 177618
rect 233240 170536 233292 170542
rect 233240 170478 233292 170484
rect 233436 148782 233464 187070
rect 233516 184408 233568 184414
rect 233516 184350 233568 184356
rect 233528 150346 233556 184350
rect 233976 180736 234028 180742
rect 233976 180678 234028 180684
rect 233700 180668 233752 180674
rect 233700 180610 233752 180616
rect 233608 177268 233660 177274
rect 233608 177210 233660 177216
rect 233516 150340 233568 150346
rect 233516 150282 233568 150288
rect 233424 148776 233476 148782
rect 233424 148718 233476 148724
rect 232412 147144 232464 147150
rect 232412 147086 232464 147092
rect 232504 146328 232556 146334
rect 232504 146270 232556 146276
rect 231822 139182 231900 139210
rect 231766 139159 231822 139168
rect 231308 138848 231360 138854
rect 231306 138816 231308 138825
rect 231360 138816 231362 138825
rect 231306 138751 231362 138760
rect 231676 137964 231728 137970
rect 231676 137906 231728 137912
rect 231688 137329 231716 137906
rect 231768 137896 231820 137902
rect 231766 137864 231768 137873
rect 231820 137864 231822 137873
rect 231766 137799 231822 137808
rect 231674 137320 231730 137329
rect 231308 137284 231360 137290
rect 231674 137255 231730 137264
rect 231308 137226 231360 137232
rect 231320 125089 231348 137226
rect 231400 136604 231452 136610
rect 231400 136546 231452 136552
rect 231412 135969 231440 136546
rect 231768 136536 231820 136542
rect 231768 136478 231820 136484
rect 231398 135960 231454 135969
rect 231398 135895 231454 135904
rect 231780 135425 231808 136478
rect 231766 135416 231822 135425
rect 231766 135351 231822 135360
rect 231676 135244 231728 135250
rect 231676 135186 231728 135192
rect 231584 135176 231636 135182
rect 231584 135118 231636 135124
rect 231596 134065 231624 135118
rect 231688 134473 231716 135186
rect 231768 135108 231820 135114
rect 231768 135050 231820 135056
rect 231780 135017 231808 135050
rect 231766 135008 231822 135017
rect 231766 134943 231822 134952
rect 231674 134464 231730 134473
rect 231674 134399 231730 134408
rect 231582 134056 231638 134065
rect 231582 133991 231638 134000
rect 231676 133884 231728 133890
rect 231676 133826 231728 133832
rect 231688 132569 231716 133826
rect 231768 133816 231820 133822
rect 231768 133758 231820 133764
rect 231780 133113 231808 133758
rect 231766 133104 231822 133113
rect 231766 133039 231822 133048
rect 231674 132560 231730 132569
rect 231674 132495 231730 132504
rect 231768 132456 231820 132462
rect 231768 132398 231820 132404
rect 231676 132388 231728 132394
rect 231676 132330 231728 132336
rect 231584 132320 231636 132326
rect 231584 132262 231636 132268
rect 231596 131209 231624 132262
rect 231688 131617 231716 132330
rect 231780 132161 231808 132398
rect 231766 132152 231822 132161
rect 231766 132087 231822 132096
rect 231674 131608 231730 131617
rect 231674 131543 231730 131552
rect 231582 131200 231638 131209
rect 231582 131135 231638 131144
rect 231492 131028 231544 131034
rect 231492 130970 231544 130976
rect 231504 130257 231532 130970
rect 231490 130248 231546 130257
rect 231490 130183 231546 130192
rect 231768 129736 231820 129742
rect 231768 129678 231820 129684
rect 231676 129532 231728 129538
rect 231676 129474 231728 129480
rect 231688 129305 231716 129474
rect 231674 129296 231730 129305
rect 231674 129231 231730 129240
rect 231780 128897 231808 129678
rect 231766 128888 231822 128897
rect 231766 128823 231822 128832
rect 231674 128344 231730 128353
rect 231584 128308 231636 128314
rect 231674 128279 231730 128288
rect 231584 128250 231636 128256
rect 231596 127401 231624 128250
rect 231688 128246 231716 128279
rect 231676 128240 231728 128246
rect 231676 128182 231728 128188
rect 231768 128172 231820 128178
rect 231768 128114 231820 128120
rect 231780 127945 231808 128114
rect 231766 127936 231822 127945
rect 231766 127871 231822 127880
rect 231582 127392 231638 127401
rect 231582 127327 231638 127336
rect 231674 126984 231730 126993
rect 231584 126948 231636 126954
rect 231674 126919 231730 126928
rect 231584 126890 231636 126896
rect 231596 126041 231624 126890
rect 231688 126818 231716 126919
rect 231768 126880 231820 126886
rect 231768 126822 231820 126828
rect 231676 126812 231728 126818
rect 231676 126754 231728 126760
rect 231780 126449 231808 126822
rect 231766 126440 231822 126449
rect 231766 126375 231822 126384
rect 231582 126032 231638 126041
rect 231582 125967 231638 125976
rect 231768 125588 231820 125594
rect 231768 125530 231820 125536
rect 231780 125497 231808 125530
rect 231766 125488 231822 125497
rect 231766 125423 231822 125432
rect 231306 125080 231362 125089
rect 231306 125015 231362 125024
rect 231768 124160 231820 124166
rect 231768 124102 231820 124108
rect 231780 123593 231808 124102
rect 231766 123584 231822 123593
rect 231308 123548 231360 123554
rect 231766 123519 231822 123528
rect 231308 123490 231360 123496
rect 231320 114617 231348 123490
rect 231584 123480 231636 123486
rect 231584 123422 231636 123428
rect 231400 122732 231452 122738
rect 231400 122674 231452 122680
rect 231412 121689 231440 122674
rect 231492 122120 231544 122126
rect 231492 122062 231544 122068
rect 231398 121680 231454 121689
rect 231398 121615 231454 121624
rect 231400 121372 231452 121378
rect 231400 121314 231452 121320
rect 231412 120329 231440 121314
rect 231504 121281 231532 122062
rect 231490 121272 231546 121281
rect 231490 121207 231546 121216
rect 231398 120320 231454 120329
rect 231398 120255 231454 120264
rect 231492 119400 231544 119406
rect 231596 119377 231624 123422
rect 231768 122800 231820 122806
rect 231768 122742 231820 122748
rect 231780 122641 231808 122742
rect 231766 122632 231822 122641
rect 231766 122567 231822 122576
rect 231768 121440 231820 121446
rect 231768 121382 231820 121388
rect 231780 120737 231808 121382
rect 231766 120728 231822 120737
rect 231766 120663 231822 120672
rect 231768 120080 231820 120086
rect 231768 120022 231820 120028
rect 231780 119785 231808 120022
rect 231766 119776 231822 119785
rect 231766 119711 231822 119720
rect 231492 119342 231544 119348
rect 231582 119368 231638 119377
rect 231504 116521 231532 119342
rect 231582 119303 231638 119312
rect 231768 118312 231820 118318
rect 231768 118254 231820 118260
rect 231676 118040 231728 118046
rect 231780 118017 231808 118254
rect 231676 117982 231728 117988
rect 231766 118008 231822 118017
rect 231490 116512 231546 116521
rect 231490 116447 231546 116456
rect 231688 116113 231716 117982
rect 231766 117943 231822 117952
rect 231768 117292 231820 117298
rect 231768 117234 231820 117240
rect 231780 117065 231808 117234
rect 231766 117056 231822 117065
rect 231766 116991 231822 117000
rect 231674 116104 231730 116113
rect 231674 116039 231730 116048
rect 231768 115932 231820 115938
rect 231768 115874 231820 115880
rect 231780 115569 231808 115874
rect 231766 115560 231822 115569
rect 231766 115495 231822 115504
rect 231306 114608 231362 114617
rect 231306 114543 231362 114552
rect 231492 114504 231544 114510
rect 231492 114446 231544 114452
rect 231504 113665 231532 114446
rect 231768 114436 231820 114442
rect 231768 114378 231820 114384
rect 231490 113656 231546 113665
rect 231490 113591 231546 113600
rect 231780 113257 231808 114378
rect 231766 113248 231822 113257
rect 231766 113183 231822 113192
rect 231228 113146 231348 113174
rect 231216 107568 231268 107574
rect 231216 107510 231268 107516
rect 231228 106593 231256 107510
rect 231214 106584 231270 106593
rect 231214 106519 231270 106528
rect 231122 100872 231178 100881
rect 231122 100807 231178 100816
rect 230848 100156 230900 100162
rect 230848 100098 230900 100104
rect 230756 99884 230808 99890
rect 230756 99826 230808 99832
rect 230768 98025 230796 99826
rect 230860 99521 230888 100098
rect 230846 99512 230902 99521
rect 230846 99447 230902 99456
rect 231032 99340 231084 99346
rect 231032 99282 231084 99288
rect 231044 98977 231072 99282
rect 231030 98968 231086 98977
rect 231030 98903 231086 98912
rect 231320 98569 231348 113146
rect 231768 113144 231820 113150
rect 231768 113086 231820 113092
rect 231676 113076 231728 113082
rect 231676 113018 231728 113024
rect 231584 112464 231636 112470
rect 231584 112406 231636 112412
rect 231492 111784 231544 111790
rect 231492 111726 231544 111732
rect 231504 110809 231532 111726
rect 231596 111353 231624 112406
rect 231688 112305 231716 113018
rect 231780 112713 231808 113086
rect 231766 112704 231822 112713
rect 231766 112639 231822 112648
rect 231674 112296 231730 112305
rect 231674 112231 231730 112240
rect 231766 111752 231822 111761
rect 231766 111687 231768 111696
rect 231820 111687 231822 111696
rect 231768 111658 231820 111664
rect 231582 111344 231638 111353
rect 231582 111279 231638 111288
rect 231490 110800 231546 110809
rect 231490 110735 231546 110744
rect 231768 110424 231820 110430
rect 231766 110392 231768 110401
rect 231820 110392 231822 110401
rect 231766 110327 231822 110336
rect 231768 109472 231820 109478
rect 231766 109440 231768 109449
rect 231820 109440 231822 109449
rect 231766 109375 231822 109384
rect 231768 108996 231820 109002
rect 231768 108938 231820 108944
rect 231676 108928 231728 108934
rect 231674 108896 231676 108905
rect 231728 108896 231730 108905
rect 231674 108831 231730 108840
rect 231780 108497 231808 108938
rect 231766 108488 231822 108497
rect 231766 108423 231822 108432
rect 231768 107636 231820 107642
rect 231768 107578 231820 107584
rect 231780 107545 231808 107578
rect 231766 107536 231822 107545
rect 231766 107471 231822 107480
rect 231492 107228 231544 107234
rect 231492 107170 231544 107176
rect 231504 107137 231532 107170
rect 231490 107128 231546 107137
rect 231490 107063 231546 107072
rect 231768 106208 231820 106214
rect 231766 106176 231768 106185
rect 231820 106176 231822 106185
rect 231676 106140 231728 106146
rect 231766 106111 231822 106120
rect 231676 106082 231728 106088
rect 231688 105233 231716 106082
rect 231674 105224 231730 105233
rect 231674 105159 231730 105168
rect 231768 104848 231820 104854
rect 231768 104790 231820 104796
rect 231780 103737 231808 104790
rect 232516 104718 232544 146270
rect 232688 145580 232740 145586
rect 232688 145522 232740 145528
rect 232596 140820 232648 140826
rect 232596 140762 232648 140768
rect 232504 104712 232556 104718
rect 232504 104654 232556 104660
rect 231766 103728 231822 103737
rect 231766 103663 231822 103672
rect 231492 103488 231544 103494
rect 231492 103430 231544 103436
rect 231504 102377 231532 103430
rect 231768 103420 231820 103426
rect 231768 103362 231820 103368
rect 231780 103329 231808 103362
rect 231766 103320 231822 103329
rect 231766 103255 231822 103264
rect 231490 102368 231546 102377
rect 231490 102303 231546 102312
rect 231768 102128 231820 102134
rect 231768 102070 231820 102076
rect 231780 101425 231808 102070
rect 231766 101416 231822 101425
rect 231766 101351 231822 101360
rect 231676 100632 231728 100638
rect 231676 100574 231728 100580
rect 231688 100473 231716 100574
rect 231674 100464 231730 100473
rect 231674 100399 231730 100408
rect 231768 99952 231820 99958
rect 231766 99920 231768 99929
rect 231820 99920 231822 99929
rect 232608 99890 232636 140762
rect 232700 106078 232728 145522
rect 233620 145042 233648 177210
rect 233712 158370 233740 180610
rect 233792 180396 233844 180402
rect 233792 180338 233844 180344
rect 233804 164830 233832 180338
rect 233884 177540 233936 177546
rect 233884 177482 233936 177488
rect 233896 177138 233924 177482
rect 233884 177132 233936 177138
rect 233884 177074 233936 177080
rect 233792 164824 233844 164830
rect 233792 164766 233844 164772
rect 233988 163878 234016 180678
rect 234080 177682 234108 240219
rect 234160 177948 234212 177954
rect 234160 177890 234212 177896
rect 234068 177676 234120 177682
rect 234068 177618 234120 177624
rect 233976 163872 234028 163878
rect 233976 163814 234028 163820
rect 233700 158364 233752 158370
rect 233700 158306 233752 158312
rect 233976 147756 234028 147762
rect 233976 147698 234028 147704
rect 233884 147688 233936 147694
rect 233884 147630 233936 147636
rect 233608 145036 233660 145042
rect 233608 144978 233660 144984
rect 233896 107574 233924 147630
rect 233884 107568 233936 107574
rect 233884 107510 233936 107516
rect 233988 107234 234016 147698
rect 234068 140072 234120 140078
rect 234068 140014 234120 140020
rect 234080 115870 234108 140014
rect 234172 138854 234200 177890
rect 234448 160614 234476 240219
rect 234620 238332 234672 238338
rect 234620 238274 234672 238280
rect 234632 164966 234660 238274
rect 235000 237998 235028 240219
rect 234988 237992 235040 237998
rect 234988 237934 235040 237940
rect 235264 233708 235316 233714
rect 235264 233650 235316 233656
rect 234896 180464 234948 180470
rect 234896 180406 234948 180412
rect 234712 178016 234764 178022
rect 234712 177958 234764 177964
rect 234724 166666 234752 177958
rect 234804 177812 234856 177818
rect 234804 177754 234856 177760
rect 234712 166660 234764 166666
rect 234712 166602 234764 166608
rect 234620 164960 234672 164966
rect 234620 164902 234672 164908
rect 234436 160608 234488 160614
rect 234436 160550 234488 160556
rect 234816 146266 234844 177754
rect 234908 153134 234936 180406
rect 235172 177880 235224 177886
rect 235172 177822 235224 177828
rect 235080 177744 235132 177750
rect 235080 177686 235132 177692
rect 234988 177200 235040 177206
rect 234988 177142 235040 177148
rect 235000 165782 235028 177142
rect 234988 165776 235040 165782
rect 234988 165718 235040 165724
rect 235092 163470 235120 177686
rect 235080 163464 235132 163470
rect 235080 163406 235132 163412
rect 234896 153128 234948 153134
rect 234896 153070 234948 153076
rect 234804 146260 234856 146266
rect 234804 146202 234856 146208
rect 235184 141710 235212 177822
rect 235276 166734 235304 233650
rect 235368 199442 235396 240219
rect 235928 240038 235956 240219
rect 235916 240032 235968 240038
rect 235916 239974 235968 239980
rect 236472 238474 236500 240219
rect 236460 238468 236512 238474
rect 236460 238410 236512 238416
rect 236644 235408 236696 235414
rect 236644 235350 236696 235356
rect 235356 199436 235408 199442
rect 235356 199378 235408 199384
rect 235632 169788 235684 169794
rect 235632 169730 235684 169736
rect 235264 166728 235316 166734
rect 235264 166670 235316 166676
rect 235356 158840 235408 158846
rect 235356 158782 235408 158788
rect 235264 149116 235316 149122
rect 235264 149058 235316 149064
rect 235172 141704 235224 141710
rect 235172 141646 235224 141652
rect 234160 138848 234212 138854
rect 234160 138790 234212 138796
rect 234252 116612 234304 116618
rect 234252 116554 234304 116560
rect 234068 115864 234120 115870
rect 234068 115806 234120 115812
rect 234160 115252 234212 115258
rect 234160 115194 234212 115200
rect 233976 107228 234028 107234
rect 233976 107170 234028 107176
rect 232688 106072 232740 106078
rect 232688 106014 232740 106020
rect 231766 99855 231822 99864
rect 232596 99884 232648 99890
rect 232596 99826 232648 99832
rect 233976 99408 234028 99414
rect 233976 99350 234028 99356
rect 233884 98660 233936 98666
rect 233884 98602 233936 98608
rect 231306 98560 231362 98569
rect 231306 98495 231362 98504
rect 231124 98048 231176 98054
rect 230754 98016 230810 98025
rect 231124 97990 231176 97996
rect 230754 97951 230810 97960
rect 230754 97064 230810 97073
rect 230754 96999 230810 97008
rect 230662 96656 230718 96665
rect 230662 96591 230718 96600
rect 230570 95840 230626 95849
rect 230570 95775 230626 95784
rect 230584 95334 230612 95775
rect 230572 95328 230624 95334
rect 230572 95270 230624 95276
rect 230676 90370 230704 96591
rect 230664 90364 230716 90370
rect 230664 90306 230716 90312
rect 229928 68400 229980 68406
rect 229928 68342 229980 68348
rect 229836 51808 229888 51814
rect 229836 51750 229888 51756
rect 230768 7614 230796 96999
rect 231136 15910 231164 97990
rect 231584 97640 231636 97646
rect 231582 97608 231584 97617
rect 231636 97608 231638 97617
rect 231582 97543 231638 97552
rect 231768 97368 231820 97374
rect 231768 97310 231820 97316
rect 231308 97300 231360 97306
rect 231308 97242 231360 97248
rect 231320 96665 231348 97242
rect 231780 97073 231808 97310
rect 231766 97064 231822 97073
rect 231766 96999 231822 97008
rect 232596 96688 232648 96694
rect 231306 96656 231362 96665
rect 232596 96630 232648 96636
rect 231306 96591 231362 96600
rect 232504 95328 232556 95334
rect 232504 95270 232556 95276
rect 231124 15904 231176 15910
rect 231124 15846 231176 15852
rect 230756 7608 230808 7614
rect 230756 7550 230808 7556
rect 232516 3534 232544 95270
rect 232608 47598 232636 96630
rect 232596 47592 232648 47598
rect 232596 47534 232648 47540
rect 229744 3528 229796 3534
rect 229744 3470 229796 3476
rect 232504 3528 232556 3534
rect 232504 3470 232556 3476
rect 233896 3466 233924 98602
rect 233988 33794 234016 99350
rect 234172 97646 234200 115194
rect 234264 100638 234292 116554
rect 235276 108594 235304 149058
rect 235368 118454 235396 158782
rect 235540 158772 235592 158778
rect 235540 158714 235592 158720
rect 235448 158024 235500 158030
rect 235448 157966 235500 157972
rect 235356 118448 235408 118454
rect 235356 118390 235408 118396
rect 235460 118318 235488 157966
rect 235552 120018 235580 158714
rect 235644 130830 235672 169730
rect 236656 153066 236684 235350
rect 236840 181694 236868 240219
rect 237288 234660 237340 234666
rect 237288 234602 237340 234608
rect 236828 181688 236880 181694
rect 236828 181630 236880 181636
rect 236644 153060 236696 153066
rect 236644 153002 236696 153008
rect 236736 150612 236788 150618
rect 236736 150554 236788 150560
rect 236644 150476 236696 150482
rect 236644 150418 236696 150424
rect 235632 130824 235684 130830
rect 235632 130766 235684 130772
rect 235540 120012 235592 120018
rect 235540 119954 235592 119960
rect 235448 118312 235500 118318
rect 235448 118254 235500 118260
rect 235540 117972 235592 117978
rect 235540 117914 235592 117920
rect 235356 113212 235408 113218
rect 235356 113154 235408 113160
rect 235264 108588 235316 108594
rect 235264 108530 235316 108536
rect 235264 103556 235316 103562
rect 235264 103498 235316 103504
rect 234252 100632 234304 100638
rect 234252 100574 234304 100580
rect 234160 97640 234212 97646
rect 234160 97582 234212 97588
rect 233976 33788 234028 33794
rect 233976 33730 234028 33736
rect 235276 11762 235304 103498
rect 235368 43450 235396 113154
rect 235552 100162 235580 117914
rect 236656 108934 236684 150418
rect 236748 110226 236776 150554
rect 236828 150544 236880 150550
rect 236828 150486 236880 150492
rect 236736 110220 236788 110226
rect 236736 110162 236788 110168
rect 236840 109478 236868 150486
rect 236828 109472 236880 109478
rect 236828 109414 236880 109420
rect 236644 108928 236696 108934
rect 236644 108870 236696 108876
rect 235540 100156 235592 100162
rect 235540 100098 235592 100104
rect 237300 97306 237328 234602
rect 237392 184414 237420 240219
rect 237944 233714 237972 240219
rect 238024 236700 238076 236706
rect 238024 236642 238076 236648
rect 237932 233708 237984 233714
rect 237932 233650 237984 233656
rect 237380 184408 237432 184414
rect 237380 184350 237432 184356
rect 238036 143478 238064 236642
rect 238116 235476 238168 235482
rect 238116 235418 238168 235424
rect 238128 202842 238156 235418
rect 238312 234666 238340 240219
rect 238872 240106 238900 240219
rect 238860 240100 238912 240106
rect 238860 240042 238912 240048
rect 239232 239426 239260 240219
rect 239220 239420 239272 239426
rect 239220 239362 239272 239368
rect 239784 238678 239812 240219
rect 239772 238672 239824 238678
rect 239772 238614 239824 238620
rect 239404 236020 239456 236026
rect 239404 235962 239456 235968
rect 238300 234660 238352 234666
rect 238300 234602 238352 234608
rect 238116 202836 238168 202842
rect 238116 202778 238168 202784
rect 239416 172378 239444 235962
rect 240336 177818 240364 240219
rect 240704 238746 240732 240219
rect 240692 238740 240744 238746
rect 240692 238682 240744 238688
rect 240876 237448 240928 237454
rect 240876 237390 240928 237396
rect 240784 236088 240836 236094
rect 240784 236030 240836 236036
rect 240324 177812 240376 177818
rect 240324 177754 240376 177760
rect 239404 172372 239456 172378
rect 239404 172314 239456 172320
rect 238300 168428 238352 168434
rect 238300 168370 238352 168376
rect 238116 167068 238168 167074
rect 238116 167010 238168 167016
rect 238024 143472 238076 143478
rect 238024 143414 238076 143420
rect 238128 128178 238156 167010
rect 238312 129538 238340 168370
rect 239496 163124 239548 163130
rect 239496 163066 239548 163072
rect 238484 158092 238536 158098
rect 238484 158034 238536 158040
rect 238392 138712 238444 138718
rect 238392 138654 238444 138660
rect 238300 129532 238352 129538
rect 238300 129474 238352 129480
rect 238208 128376 238260 128382
rect 238208 128318 238260 128324
rect 238116 128172 238168 128178
rect 238116 128114 238168 128120
rect 238024 118720 238076 118726
rect 238024 118662 238076 118668
rect 237288 97300 237340 97306
rect 237288 97242 237340 97248
rect 236644 96756 236696 96762
rect 236644 96698 236696 96704
rect 236656 49026 236684 96698
rect 236644 49020 236696 49026
rect 236644 48962 236696 48968
rect 235356 43444 235408 43450
rect 235356 43386 235408 43392
rect 238036 36582 238064 118662
rect 238116 99476 238168 99482
rect 238116 99418 238168 99424
rect 238024 36576 238076 36582
rect 238024 36518 238076 36524
rect 238128 21418 238156 99418
rect 238220 57254 238248 128318
rect 238300 116204 238352 116210
rect 238300 116146 238352 116152
rect 238312 77994 238340 116146
rect 238404 99958 238432 138654
rect 238496 128246 238524 158034
rect 238484 128240 238536 128246
rect 238484 128182 238536 128188
rect 239404 127016 239456 127022
rect 239404 126958 239456 126964
rect 238392 99952 238444 99958
rect 238392 99894 238444 99900
rect 238300 77988 238352 77994
rect 238300 77930 238352 77936
rect 238208 57248 238260 57254
rect 238208 57190 238260 57196
rect 239416 22778 239444 126958
rect 239508 124166 239536 163066
rect 240796 160002 240824 236030
rect 240888 165578 240916 237390
rect 241256 178838 241284 240219
rect 241244 178832 241296 178838
rect 241244 178774 241296 178780
rect 241060 173936 241112 173942
rect 241060 173878 241112 173884
rect 240968 166320 241020 166326
rect 240968 166262 241020 166268
rect 240876 165572 240928 165578
rect 240876 165514 240928 165520
rect 240784 159996 240836 160002
rect 240784 159938 240836 159944
rect 240876 155984 240928 155990
rect 240876 155926 240928 155932
rect 240784 135516 240836 135522
rect 240784 135458 240836 135464
rect 239496 124160 239548 124166
rect 239496 124102 239548 124108
rect 239496 114572 239548 114578
rect 239496 114514 239548 114520
rect 239508 76566 239536 114514
rect 239496 76560 239548 76566
rect 239496 76502 239548 76508
rect 239404 22772 239456 22778
rect 239404 22714 239456 22720
rect 238116 21412 238168 21418
rect 238116 21354 238168 21360
rect 235264 11756 235316 11762
rect 235264 11698 235316 11704
rect 240796 7682 240824 135458
rect 240888 115938 240916 155926
rect 240980 126818 241008 166262
rect 241072 135114 241100 173878
rect 241152 160132 241204 160138
rect 241152 160074 241204 160080
rect 241164 144838 241192 160074
rect 241808 145654 241836 240219
rect 242176 160138 242204 240219
rect 242728 238406 242756 240219
rect 242900 240168 242952 240174
rect 242900 240110 242952 240116
rect 242716 238400 242768 238406
rect 242716 238342 242768 238348
rect 242912 175166 242940 240110
rect 243280 236026 243308 240219
rect 243544 239896 243596 239902
rect 243544 239838 243596 239844
rect 243556 239766 243584 239838
rect 243452 239760 243504 239766
rect 243452 239702 243504 239708
rect 243544 239760 243596 239766
rect 243544 239702 243596 239708
rect 243464 239562 243492 239702
rect 243452 239556 243504 239562
rect 243452 239498 243504 239504
rect 243268 236020 243320 236026
rect 243268 235962 243320 235968
rect 243648 178770 243676 240219
rect 243820 240168 243872 240174
rect 243820 240110 243872 240116
rect 243832 239986 243860 240110
rect 243740 239958 243860 239986
rect 243910 240000 243966 240009
rect 243740 238542 243768 239958
rect 243910 239935 243966 239944
rect 243820 239896 243872 239902
rect 243820 239838 243872 239844
rect 243832 238610 243860 239838
rect 243924 238746 243952 239935
rect 243912 238740 243964 238746
rect 243912 238682 243964 238688
rect 243820 238604 243872 238610
rect 243820 238546 243872 238552
rect 243728 238536 243780 238542
rect 243728 238478 243780 238484
rect 243636 178764 243688 178770
rect 243636 178706 243688 178712
rect 242900 175160 242952 175166
rect 242900 175102 242952 175108
rect 244016 168230 244044 244287
rect 244004 168224 244056 168230
rect 244004 168166 244056 168172
rect 242440 167136 242492 167142
rect 242440 167078 242492 167084
rect 242164 160132 242216 160138
rect 242164 160074 242216 160080
rect 242256 160132 242308 160138
rect 242256 160074 242308 160080
rect 241796 145648 241848 145654
rect 241796 145590 241848 145596
rect 241152 144832 241204 144838
rect 241152 144774 241204 144780
rect 241244 144220 241296 144226
rect 241244 144162 241296 144168
rect 241060 135108 241112 135114
rect 241060 135050 241112 135056
rect 241060 129940 241112 129946
rect 241060 129882 241112 129888
rect 240968 126812 241020 126818
rect 240968 126754 241020 126760
rect 240968 122868 241020 122874
rect 240968 122810 241020 122816
rect 240876 115932 240928 115938
rect 240876 115874 240928 115880
rect 240876 110492 240928 110498
rect 240876 110434 240928 110440
rect 240888 25634 240916 110434
rect 240980 50454 241008 122810
rect 241072 61402 241100 129882
rect 241152 118788 241204 118794
rect 241152 118730 241204 118736
rect 241164 62830 241192 118730
rect 241256 106214 241284 144162
rect 242164 138032 242216 138038
rect 242164 137974 242216 137980
rect 241244 106208 241296 106214
rect 241244 106150 241296 106156
rect 241152 62824 241204 62830
rect 241152 62766 241204 62772
rect 241060 61396 241112 61402
rect 241060 61338 241112 61344
rect 240968 50448 241020 50454
rect 240968 50390 241020 50396
rect 240876 25628 240928 25634
rect 240876 25570 240928 25576
rect 242176 10402 242204 137974
rect 242268 120086 242296 160074
rect 242348 153264 242400 153270
rect 242348 153206 242400 153212
rect 242256 120080 242308 120086
rect 242256 120022 242308 120028
rect 242360 113082 242388 153206
rect 242452 128314 242480 167078
rect 244108 157282 244136 250543
rect 244186 241904 244242 241913
rect 244186 241839 244242 241848
rect 244200 177750 244228 241839
rect 244280 240780 244332 240786
rect 244280 240722 244332 240728
rect 244292 239902 244320 240722
rect 244280 239896 244332 239902
rect 244280 239838 244332 239844
rect 244188 177744 244240 177750
rect 244188 177686 244240 177692
rect 244096 157276 244148 157282
rect 244096 157218 244148 157224
rect 243636 151836 243688 151842
rect 243636 151778 243688 151784
rect 242624 144968 242676 144974
rect 242624 144910 242676 144916
rect 242532 132524 242584 132530
rect 242532 132466 242584 132472
rect 242440 128308 242492 128314
rect 242440 128250 242492 128256
rect 242440 122936 242492 122942
rect 242440 122878 242492 122884
rect 242348 113076 242400 113082
rect 242348 113018 242400 113024
rect 242256 111852 242308 111858
rect 242256 111794 242308 111800
rect 242268 26926 242296 111794
rect 242348 109064 242400 109070
rect 242348 109006 242400 109012
rect 242360 39438 242388 109006
rect 242452 53174 242480 122878
rect 242544 83570 242572 132466
rect 242636 103426 242664 144910
rect 243544 139460 243596 139466
rect 243544 139402 243596 139408
rect 242624 103420 242676 103426
rect 242624 103362 242676 103368
rect 242532 83564 242584 83570
rect 242532 83506 242584 83512
rect 243556 65618 243584 139402
rect 243648 110430 243676 151778
rect 244384 142050 244412 271487
rect 244476 237454 244504 283902
rect 244646 273728 244702 273737
rect 244646 273663 244702 273672
rect 244554 273184 244610 273193
rect 244554 273119 244610 273128
rect 244464 237448 244516 237454
rect 244464 237390 244516 237396
rect 244568 159934 244596 273119
rect 244660 175098 244688 273663
rect 244738 270192 244794 270201
rect 244738 270127 244794 270136
rect 244648 175092 244700 175098
rect 244648 175034 244700 175040
rect 244752 173806 244780 270127
rect 244830 264480 244886 264489
rect 244830 264415 244886 264424
rect 244740 173800 244792 173806
rect 244740 173742 244792 173748
rect 244844 172514 244872 264415
rect 244936 260681 244964 500958
rect 245660 289196 245712 289202
rect 245660 289138 245712 289144
rect 245672 283801 245700 289138
rect 246120 287768 246172 287774
rect 246120 287710 246172 287716
rect 246026 284880 246082 284889
rect 246026 284815 246082 284824
rect 245658 283792 245714 283801
rect 245658 283727 245714 283736
rect 245198 283248 245254 283257
rect 245198 283183 245254 283192
rect 245014 262304 245070 262313
rect 245014 262239 245070 262248
rect 244922 260672 244978 260681
rect 244922 260607 244978 260616
rect 244922 255232 244978 255241
rect 244922 255167 244978 255176
rect 244832 172508 244884 172514
rect 244832 172450 244884 172456
rect 244936 164218 244964 255167
rect 245028 172446 245056 262239
rect 245106 260944 245162 260953
rect 245106 260879 245162 260888
rect 245016 172440 245068 172446
rect 245016 172382 245068 172388
rect 244924 164212 244976 164218
rect 244924 164154 244976 164160
rect 244556 159928 244608 159934
rect 244556 159870 244608 159876
rect 245120 144906 245148 260879
rect 245108 144900 245160 144906
rect 245108 144842 245160 144848
rect 245212 143546 245240 283183
rect 245936 282872 245988 282878
rect 245936 282814 245988 282820
rect 245842 282432 245898 282441
rect 245842 282367 245898 282376
rect 245658 281072 245714 281081
rect 245658 281007 245714 281016
rect 245672 280294 245700 281007
rect 245660 280288 245712 280294
rect 245660 280230 245712 280236
rect 245658 279440 245714 279449
rect 245658 279375 245714 279384
rect 245672 278798 245700 279375
rect 245660 278792 245712 278798
rect 245660 278734 245712 278740
rect 245752 275936 245804 275942
rect 245750 275904 245752 275913
rect 245804 275904 245806 275913
rect 245750 275839 245806 275848
rect 245750 274544 245806 274553
rect 245750 274479 245806 274488
rect 245764 273290 245792 274479
rect 245752 273284 245804 273290
rect 245752 273226 245804 273232
rect 245750 272368 245806 272377
rect 245750 272303 245806 272312
rect 245764 271998 245792 272303
rect 245752 271992 245804 271998
rect 245752 271934 245804 271940
rect 245750 269648 245806 269657
rect 245750 269583 245806 269592
rect 245764 269142 245792 269583
rect 245752 269136 245804 269142
rect 245752 269078 245804 269084
rect 245658 268832 245714 268841
rect 245658 268767 245714 268776
rect 245672 267850 245700 268767
rect 245750 268016 245806 268025
rect 245750 267951 245806 267960
rect 245660 267844 245712 267850
rect 245660 267786 245712 267792
rect 245764 267782 245792 267951
rect 245752 267776 245804 267782
rect 245752 267718 245804 267724
rect 245750 267472 245806 267481
rect 245750 267407 245806 267416
rect 245660 266756 245712 266762
rect 245660 266698 245712 266704
rect 245672 263945 245700 266698
rect 245764 266490 245792 267407
rect 245752 266484 245804 266490
rect 245752 266426 245804 266432
rect 245750 265840 245806 265849
rect 245750 265775 245806 265784
rect 245764 265169 245792 265775
rect 245750 265160 245806 265169
rect 245750 265095 245806 265104
rect 245658 263936 245714 263945
rect 245658 263871 245714 263880
rect 245750 263120 245806 263129
rect 245750 263055 245806 263064
rect 245658 261760 245714 261769
rect 245658 261695 245714 261704
rect 245672 252521 245700 261695
rect 245764 259162 245792 263055
rect 245856 259350 245884 282367
rect 245948 281625 245976 282814
rect 245934 281616 245990 281625
rect 245934 281551 245990 281560
rect 245934 280256 245990 280265
rect 245934 280191 245936 280200
rect 245988 280191 245990 280200
rect 245936 280162 245988 280168
rect 246040 280106 246068 284815
rect 245948 280078 246068 280106
rect 245948 266762 245976 280078
rect 246132 277394 246160 287710
rect 246040 277366 246160 277394
rect 245936 266756 245988 266762
rect 245936 266698 245988 266704
rect 245934 266656 245990 266665
rect 245934 266591 245990 266600
rect 245948 266422 245976 266591
rect 245936 266416 245988 266422
rect 245936 266358 245988 266364
rect 245934 259584 245990 259593
rect 245934 259519 245990 259528
rect 245948 259486 245976 259519
rect 245936 259480 245988 259486
rect 245936 259422 245988 259428
rect 245844 259344 245896 259350
rect 245844 259286 245896 259292
rect 245764 259134 245976 259162
rect 245844 259072 245896 259078
rect 245844 259014 245896 259020
rect 245750 258768 245806 258777
rect 245750 258703 245806 258712
rect 245764 258126 245792 258703
rect 245752 258120 245804 258126
rect 245752 258062 245804 258068
rect 245750 256592 245806 256601
rect 245750 256527 245806 256536
rect 245764 255338 245792 256527
rect 245752 255332 245804 255338
rect 245752 255274 245804 255280
rect 245658 252512 245714 252521
rect 245658 252447 245714 252456
rect 245750 248704 245806 248713
rect 245750 248639 245806 248648
rect 245660 248396 245712 248402
rect 245660 248338 245712 248344
rect 245672 247353 245700 248338
rect 245658 247344 245714 247353
rect 245658 247279 245714 247288
rect 245660 244248 245712 244254
rect 245660 244190 245712 244196
rect 245672 243001 245700 244190
rect 245658 242992 245714 243001
rect 245658 242927 245714 242936
rect 245658 241632 245714 241641
rect 245658 241567 245714 241576
rect 245292 240916 245344 240922
rect 245292 240858 245344 240864
rect 245304 240009 245332 240858
rect 245290 240000 245346 240009
rect 245290 239935 245346 239944
rect 245292 239896 245344 239902
rect 245292 239838 245344 239844
rect 245304 239426 245332 239838
rect 245292 239420 245344 239426
rect 245292 239362 245344 239368
rect 245672 235482 245700 241567
rect 245764 236706 245792 248639
rect 245752 236700 245804 236706
rect 245752 236642 245804 236648
rect 245856 236094 245884 259014
rect 245844 236088 245896 236094
rect 245844 236030 245896 236036
rect 245660 235476 245712 235482
rect 245660 235418 245712 235424
rect 245948 229770 245976 259134
rect 246040 256834 246068 277366
rect 246120 276004 246172 276010
rect 246120 275946 246172 275952
rect 246132 275369 246160 275946
rect 246118 275360 246174 275369
rect 246118 275295 246174 275304
rect 246120 266348 246172 266354
rect 246120 266290 246172 266296
rect 246132 265305 246160 266290
rect 246118 265296 246174 265305
rect 246118 265231 246174 265240
rect 246118 265160 246174 265169
rect 246118 265095 246174 265104
rect 246028 256828 246080 256834
rect 246028 256770 246080 256776
rect 246028 256692 246080 256698
rect 246028 256634 246080 256640
rect 246040 256057 246068 256634
rect 246026 256048 246082 256057
rect 246026 255983 246082 255992
rect 246026 253872 246082 253881
rect 246026 253807 246082 253816
rect 246040 252618 246068 253807
rect 246028 252612 246080 252618
rect 246028 252554 246080 252560
rect 246026 251696 246082 251705
rect 246026 251631 246082 251640
rect 246040 251258 246068 251631
rect 246028 251252 246080 251258
rect 246028 251194 246080 251200
rect 246026 250336 246082 250345
rect 246026 250271 246082 250280
rect 246040 249830 246068 250271
rect 246028 249824 246080 249830
rect 246028 249766 246080 249772
rect 246028 248192 246080 248198
rect 246026 248160 246028 248169
rect 246080 248160 246082 248169
rect 246026 248095 246082 248104
rect 246028 247036 246080 247042
rect 246028 246978 246080 246984
rect 246040 246537 246068 246978
rect 246026 246528 246082 246537
rect 246026 246463 246082 246472
rect 246026 245984 246082 245993
rect 246026 245919 246082 245928
rect 246040 245682 246068 245919
rect 246028 245676 246080 245682
rect 246028 245618 246080 245624
rect 246026 243808 246082 243817
rect 246026 243743 246082 243752
rect 246040 242962 246068 243743
rect 246028 242956 246080 242962
rect 246028 242898 246080 242904
rect 246028 241460 246080 241466
rect 246028 241402 246080 241408
rect 246040 240281 246068 241402
rect 246026 240272 246082 240281
rect 246026 240207 246082 240216
rect 246132 235414 246160 265095
rect 246224 256970 246252 683130
rect 246856 312588 246908 312594
rect 246856 312530 246908 312536
rect 246302 276720 246358 276729
rect 246302 276655 246358 276664
rect 246212 256964 246264 256970
rect 246212 256906 246264 256912
rect 246212 256828 246264 256834
rect 246212 256770 246264 256776
rect 246224 254425 246252 256770
rect 246210 254416 246266 254425
rect 246210 254351 246266 254360
rect 246120 235408 246172 235414
rect 246120 235350 246172 235356
rect 245936 229764 245988 229770
rect 245936 229706 245988 229712
rect 246316 176118 246344 276655
rect 246394 271008 246450 271017
rect 246394 270943 246450 270952
rect 246408 177585 246436 270943
rect 246486 258224 246542 258233
rect 246486 258159 246488 258168
rect 246540 258159 246542 258168
rect 246488 258130 246540 258136
rect 246670 257408 246726 257417
rect 246670 257343 246726 257352
rect 246488 256964 246540 256970
rect 246488 256906 246540 256912
rect 246500 252249 246528 256906
rect 246578 253056 246634 253065
rect 246578 252991 246634 253000
rect 246486 252240 246542 252249
rect 246486 252175 246542 252184
rect 246488 252136 246540 252142
rect 246488 252078 246540 252084
rect 246394 177576 246450 177585
rect 246394 177511 246450 177520
rect 246304 176112 246356 176118
rect 246304 176054 246356 176060
rect 246500 176050 246528 252078
rect 246592 177886 246620 252991
rect 246684 252142 246712 257343
rect 246672 252136 246724 252142
rect 246672 252078 246724 252084
rect 246868 249529 246896 312530
rect 247132 288652 247184 288658
rect 247132 288594 247184 288600
rect 247040 286272 247092 286278
rect 247040 286214 247092 286220
rect 246854 249520 246910 249529
rect 246854 249455 246910 249464
rect 246670 242448 246726 242457
rect 246670 242383 246726 242392
rect 246684 180402 246712 242383
rect 246672 180396 246724 180402
rect 246672 180338 246724 180344
rect 246580 177880 246632 177886
rect 246580 177822 246632 177828
rect 246488 176044 246540 176050
rect 246488 175986 246540 175992
rect 245292 146940 245344 146946
rect 245292 146882 245344 146888
rect 245200 143540 245252 143546
rect 245200 143482 245252 143488
rect 245200 142180 245252 142186
rect 245200 142122 245252 142128
rect 244372 142044 244424 142050
rect 244372 141986 244424 141992
rect 244280 140888 244332 140894
rect 244280 140830 244332 140836
rect 244292 140146 244320 140830
rect 244280 140140 244332 140146
rect 244280 140082 244332 140088
rect 245108 128444 245160 128450
rect 245108 128386 245160 128392
rect 245016 127084 245068 127090
rect 245016 127026 245068 127032
rect 244924 117428 244976 117434
rect 244924 117370 244976 117376
rect 243728 114640 243780 114646
rect 243728 114582 243780 114588
rect 243636 110424 243688 110430
rect 243636 110366 243688 110372
rect 243740 73846 243768 114582
rect 243728 73840 243780 73846
rect 243728 73782 243780 73788
rect 243544 65612 243596 65618
rect 243544 65554 243596 65560
rect 242440 53168 242492 53174
rect 242440 53110 242492 53116
rect 242348 39432 242400 39438
rect 242348 39374 242400 39380
rect 244936 31074 244964 117370
rect 245028 50386 245056 127026
rect 245120 54534 245148 128386
rect 245212 116686 245240 142122
rect 245200 116680 245252 116686
rect 245200 116622 245252 116628
rect 245304 114442 245332 146882
rect 246488 139528 246540 139534
rect 246488 139470 246540 139476
rect 245292 114436 245344 114442
rect 245292 114378 245344 114384
rect 246396 113348 246448 113354
rect 246396 113290 246448 113296
rect 245200 113280 245252 113286
rect 245200 113222 245252 113228
rect 245212 72486 245240 113222
rect 246304 109132 246356 109138
rect 246304 109074 246356 109080
rect 245200 72480 245252 72486
rect 245200 72422 245252 72428
rect 245108 54528 245160 54534
rect 245108 54470 245160 54476
rect 245016 50380 245068 50386
rect 245016 50322 245068 50328
rect 244924 31068 244976 31074
rect 244924 31010 244976 31016
rect 242256 26920 242308 26926
rect 242256 26862 242308 26868
rect 246316 24206 246344 109074
rect 246408 32434 246436 113290
rect 246500 64258 246528 139470
rect 247052 137902 247080 286214
rect 247144 150414 247172 288594
rect 247224 287836 247276 287842
rect 247224 287778 247276 287784
rect 247236 169726 247264 287778
rect 247316 284912 247368 284918
rect 247316 284854 247368 284860
rect 247224 169720 247276 169726
rect 247224 169662 247276 169668
rect 247328 168298 247356 284854
rect 247696 239358 247724 700266
rect 249064 643136 249116 643142
rect 249064 643078 249116 643084
rect 248604 287564 248656 287570
rect 248604 287506 248656 287512
rect 248512 286340 248564 286346
rect 248512 286282 248564 286288
rect 248418 286240 248474 286249
rect 248418 286175 248474 286184
rect 247776 286136 247828 286142
rect 247776 286078 247828 286084
rect 247684 239352 247736 239358
rect 247684 239294 247736 239300
rect 247316 168292 247368 168298
rect 247316 168234 247368 168240
rect 247132 150408 247184 150414
rect 247132 150350 247184 150356
rect 247040 137896 247092 137902
rect 247040 137838 247092 137844
rect 247684 127152 247736 127158
rect 247684 127094 247736 127100
rect 246580 102400 246632 102406
rect 246580 102342 246632 102348
rect 246488 64252 246540 64258
rect 246488 64194 246540 64200
rect 246592 40730 246620 102342
rect 246580 40724 246632 40730
rect 246580 40666 246632 40672
rect 246396 32428 246448 32434
rect 246396 32370 246448 32376
rect 246304 24200 246356 24206
rect 246304 24142 246356 24148
rect 247696 24138 247724 127094
rect 247788 96422 247816 286078
rect 247868 124228 247920 124234
rect 247868 124170 247920 124176
rect 247776 96416 247828 96422
rect 247776 96358 247828 96364
rect 247880 60110 247908 124170
rect 248432 97374 248460 286175
rect 248524 142118 248552 286282
rect 248616 161430 248644 287506
rect 248696 287496 248748 287502
rect 248696 287438 248748 287444
rect 248708 168366 248736 287438
rect 248788 286544 248840 286550
rect 248788 286486 248840 286492
rect 248800 171086 248828 286486
rect 248972 244316 249024 244322
rect 248972 244258 249024 244264
rect 248984 239902 249012 244258
rect 249076 239970 249104 643078
rect 250444 536852 250496 536858
rect 250444 536794 250496 536800
rect 250076 288720 250128 288726
rect 250076 288662 250128 288668
rect 249892 288516 249944 288522
rect 249892 288458 249944 288464
rect 249800 287088 249852 287094
rect 249800 287030 249852 287036
rect 249156 285116 249208 285122
rect 249156 285058 249208 285064
rect 249064 239964 249116 239970
rect 249064 239906 249116 239912
rect 248972 239896 249024 239902
rect 248972 239838 249024 239844
rect 249168 193186 249196 285058
rect 249248 284436 249300 284442
rect 249248 284378 249300 284384
rect 249260 206990 249288 284378
rect 249432 242208 249484 242214
rect 249432 242150 249484 242156
rect 249444 238474 249472 242150
rect 249432 238468 249484 238474
rect 249432 238410 249484 238416
rect 249248 206984 249300 206990
rect 249248 206926 249300 206932
rect 249156 193180 249208 193186
rect 249156 193122 249208 193128
rect 249248 174548 249300 174554
rect 249248 174490 249300 174496
rect 248788 171080 248840 171086
rect 248788 171022 248840 171028
rect 248696 168360 248748 168366
rect 248696 168302 248748 168308
rect 249156 165776 249208 165782
rect 249156 165718 249208 165724
rect 248604 161424 248656 161430
rect 248604 161366 248656 161372
rect 249064 153332 249116 153338
rect 249064 153274 249116 153280
rect 248512 142112 248564 142118
rect 248512 142054 248564 142060
rect 249076 113150 249104 153274
rect 249168 126886 249196 165718
rect 249156 126880 249208 126886
rect 249156 126822 249208 126828
rect 249156 120148 249208 120154
rect 249156 120090 249208 120096
rect 249064 113144 249116 113150
rect 249064 113086 249116 113092
rect 249064 107908 249116 107914
rect 249064 107850 249116 107856
rect 248420 97368 248472 97374
rect 248420 97310 248472 97316
rect 247868 60104 247920 60110
rect 247868 60046 247920 60052
rect 247684 24132 247736 24138
rect 247684 24074 247736 24080
rect 249076 17338 249104 107850
rect 249168 37942 249196 120090
rect 249260 99346 249288 174490
rect 249432 169856 249484 169862
rect 249432 169798 249484 169804
rect 249340 136740 249392 136746
rect 249340 136682 249392 136688
rect 249248 99340 249300 99346
rect 249248 99282 249300 99288
rect 249352 62898 249380 136682
rect 249444 132326 249472 169798
rect 249524 164280 249576 164286
rect 249524 164222 249576 164228
rect 249536 137290 249564 164222
rect 249812 137970 249840 287030
rect 249904 140690 249932 288458
rect 249984 287156 250036 287162
rect 249984 287098 250036 287104
rect 249996 149054 250024 287098
rect 250088 155922 250116 288662
rect 250168 285184 250220 285190
rect 250168 285126 250220 285132
rect 250180 157350 250208 285126
rect 250456 239562 250484 536794
rect 250628 324352 250680 324358
rect 250628 324294 250680 324300
rect 250536 285728 250588 285734
rect 250536 285670 250588 285676
rect 250444 239556 250496 239562
rect 250444 239498 250496 239504
rect 250168 157344 250220 157350
rect 250168 157286 250220 157292
rect 250076 155916 250128 155922
rect 250076 155858 250128 155864
rect 249984 149048 250036 149054
rect 249984 148990 250036 148996
rect 249892 140684 249944 140690
rect 249892 140626 249944 140632
rect 249800 137964 249852 137970
rect 249800 137906 249852 137912
rect 249524 137284 249576 137290
rect 249524 137226 249576 137232
rect 250444 136808 250496 136814
rect 250444 136750 250496 136756
rect 249432 132320 249484 132326
rect 249432 132262 249484 132268
rect 249432 125792 249484 125798
rect 249432 125734 249484 125740
rect 249444 80714 249472 125734
rect 249524 100768 249576 100774
rect 249524 100710 249576 100716
rect 249432 80708 249484 80714
rect 249432 80650 249484 80656
rect 249536 69698 249564 100710
rect 249524 69692 249576 69698
rect 249524 69634 249576 69640
rect 249340 62892 249392 62898
rect 249340 62834 249392 62840
rect 249156 37936 249208 37942
rect 249156 37878 249208 37884
rect 249064 17332 249116 17338
rect 249064 17274 249116 17280
rect 250456 11830 250484 136750
rect 250548 96354 250576 285670
rect 250640 248198 250668 324294
rect 250720 298172 250772 298178
rect 250720 298114 250772 298120
rect 250628 248192 250680 248198
rect 250628 248134 250680 248140
rect 250732 239766 250760 298114
rect 251364 288788 251416 288794
rect 251364 288730 251416 288736
rect 251272 288584 251324 288590
rect 251272 288526 251324 288532
rect 251180 287632 251232 287638
rect 251180 287574 251232 287580
rect 250720 239760 250772 239766
rect 250720 239702 250772 239708
rect 250812 172576 250864 172582
rect 250812 172518 250864 172524
rect 250720 171148 250772 171154
rect 250720 171090 250772 171096
rect 250628 160200 250680 160206
rect 250628 160142 250680 160148
rect 250640 121378 250668 160142
rect 250732 132394 250760 171090
rect 250824 133754 250852 172518
rect 250996 154624 251048 154630
rect 250996 154566 251048 154572
rect 250904 145036 250956 145042
rect 250904 144978 250956 144984
rect 250812 133748 250864 133754
rect 250812 133690 250864 133696
rect 250720 132388 250772 132394
rect 250720 132330 250772 132336
rect 250812 131300 250864 131306
rect 250812 131242 250864 131248
rect 250628 121372 250680 121378
rect 250628 121314 250680 121320
rect 250720 120216 250772 120222
rect 250720 120158 250772 120164
rect 250628 105052 250680 105058
rect 250628 104994 250680 105000
rect 250536 96348 250588 96354
rect 250536 96290 250588 96296
rect 250640 13122 250668 104994
rect 250732 42090 250760 120158
rect 250824 82142 250852 131242
rect 250916 104854 250944 144978
rect 251008 123554 251036 154566
rect 251192 140758 251220 287574
rect 251284 147626 251312 288526
rect 251376 158710 251404 288730
rect 251548 284844 251600 284850
rect 251548 284786 251600 284792
rect 251456 284028 251508 284034
rect 251456 283970 251508 283976
rect 251364 158704 251416 158710
rect 251364 158646 251416 158652
rect 251468 153202 251496 283970
rect 251560 173874 251588 284786
rect 251836 239834 251864 700674
rect 283852 696250 283880 703520
rect 300136 700670 300164 703520
rect 300124 700664 300176 700670
rect 300124 700606 300176 700612
rect 332520 700602 332548 703520
rect 332508 700596 332560 700602
rect 332508 700538 332560 700544
rect 348804 699718 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 347044 699712 347096 699718
rect 347044 699654 347096 699660
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 253204 696244 253256 696250
rect 253204 696186 253256 696192
rect 283840 696244 283892 696250
rect 283840 696186 283892 696192
rect 251916 430636 251968 430642
rect 251916 430578 251968 430584
rect 251928 248402 251956 430578
rect 252008 284572 252060 284578
rect 252008 284514 252060 284520
rect 251916 248396 251968 248402
rect 251916 248338 251968 248344
rect 251824 239828 251876 239834
rect 251824 239770 251876 239776
rect 252020 179382 252048 284514
rect 253216 238678 253244 696186
rect 295984 683188 296036 683194
rect 295984 683130 296036 683136
rect 260104 630692 260156 630698
rect 260104 630634 260156 630640
rect 255964 616888 256016 616894
rect 255964 616830 256016 616836
rect 253294 284336 253350 284345
rect 253294 284271 253350 284280
rect 253204 238672 253256 238678
rect 253204 238614 253256 238620
rect 252008 179376 252060 179382
rect 252008 179318 252060 179324
rect 251548 173868 251600 173874
rect 251548 173810 251600 173816
rect 252100 172644 252152 172650
rect 252100 172586 252152 172592
rect 251824 171216 251876 171222
rect 251824 171158 251876 171164
rect 251456 153196 251508 153202
rect 251456 153138 251508 153144
rect 251272 147620 251324 147626
rect 251272 147562 251324 147568
rect 251180 140752 251232 140758
rect 251180 140694 251232 140700
rect 251836 132462 251864 171158
rect 251916 151904 251968 151910
rect 251916 151846 251968 151852
rect 251824 132456 251876 132462
rect 251824 132398 251876 132404
rect 250996 123548 251048 123554
rect 250996 123490 251048 123496
rect 251824 116068 251876 116074
rect 251824 116010 251876 116016
rect 250996 111920 251048 111926
rect 250996 111862 251048 111868
rect 250904 104848 250956 104854
rect 250904 104790 250956 104796
rect 250812 82136 250864 82142
rect 250812 82078 250864 82084
rect 251008 72554 251036 111862
rect 250996 72548 251048 72554
rect 250996 72490 251048 72496
rect 250720 42084 250772 42090
rect 250720 42026 250772 42032
rect 251836 25566 251864 116010
rect 251928 112470 251956 151846
rect 252008 138100 252060 138106
rect 252008 138042 252060 138048
rect 251916 112464 251968 112470
rect 251916 112406 251968 112412
rect 251916 106480 251968 106486
rect 251916 106422 251968 106428
rect 251824 25560 251876 25566
rect 251824 25502 251876 25508
rect 251928 18630 251956 106422
rect 252020 66978 252048 138042
rect 252112 135182 252140 172586
rect 252284 156664 252336 156670
rect 252284 156606 252336 156612
rect 252192 143608 252244 143614
rect 252192 143550 252244 143556
rect 252100 135176 252152 135182
rect 252100 135118 252152 135124
rect 252100 118856 252152 118862
rect 252100 118798 252152 118804
rect 252008 66972 252060 66978
rect 252008 66914 252060 66920
rect 252112 61470 252140 118798
rect 252204 103494 252232 143550
rect 252296 117298 252324 156606
rect 253204 138168 253256 138174
rect 253204 138110 253256 138116
rect 252284 117292 252336 117298
rect 252284 117234 252336 117240
rect 252284 111988 252336 111994
rect 252284 111930 252336 111936
rect 252192 103488 252244 103494
rect 252192 103430 252244 103436
rect 252296 73914 252324 111930
rect 252284 73908 252336 73914
rect 252284 73850 252336 73856
rect 252100 61464 252152 61470
rect 252100 61406 252152 61412
rect 251916 18624 251968 18630
rect 251916 18566 251968 18572
rect 250628 13116 250680 13122
rect 250628 13058 250680 13064
rect 250444 11824 250496 11830
rect 250444 11766 250496 11772
rect 242164 10396 242216 10402
rect 242164 10338 242216 10344
rect 253216 9042 253244 138110
rect 253308 73166 253336 284271
rect 255976 247042 256004 616830
rect 258724 470620 258776 470626
rect 258724 470562 258776 470568
rect 256056 285048 256108 285054
rect 256056 284990 256108 284996
rect 255964 247036 256016 247042
rect 255964 246978 256016 246984
rect 256068 219434 256096 284990
rect 258736 275942 258764 470562
rect 258724 275936 258776 275942
rect 258724 275878 258776 275884
rect 258724 271924 258776 271930
rect 258724 271866 258776 271872
rect 258736 237386 258764 271866
rect 260116 237998 260144 630634
rect 294604 524476 294656 524482
rect 294604 524418 294656 524424
rect 286324 484424 286376 484430
rect 286324 484366 286376 484372
rect 280896 286612 280948 286618
rect 280896 286554 280948 286560
rect 278044 286204 278096 286210
rect 278044 286146 278096 286152
rect 265624 285932 265676 285938
rect 265624 285874 265676 285880
rect 260194 284608 260250 284617
rect 260194 284543 260250 284552
rect 260104 237992 260156 237998
rect 260104 237934 260156 237940
rect 258724 237380 258776 237386
rect 258724 237322 258776 237328
rect 256056 219428 256108 219434
rect 256056 219370 256108 219376
rect 258908 174072 258960 174078
rect 258908 174014 258960 174020
rect 256148 174004 256200 174010
rect 256148 173946 256200 173952
rect 253480 172712 253532 172718
rect 253480 172654 253532 172660
rect 253388 169924 253440 169930
rect 253388 169866 253440 169872
rect 253400 131034 253428 169866
rect 253492 133822 253520 172654
rect 254676 165708 254728 165714
rect 254676 165650 254728 165656
rect 254584 164348 254636 164354
rect 254584 164290 254636 164296
rect 253664 157412 253716 157418
rect 253664 157354 253716 157360
rect 253480 133816 253532 133822
rect 253480 133758 253532 133764
rect 253572 131232 253624 131238
rect 253572 131174 253624 131180
rect 253388 131028 253440 131034
rect 253388 130970 253440 130976
rect 253480 121644 253532 121650
rect 253480 121586 253532 121592
rect 253388 109200 253440 109206
rect 253388 109142 253440 109148
rect 253296 73160 253348 73166
rect 253296 73102 253348 73108
rect 253400 22846 253428 109142
rect 253492 47666 253520 121586
rect 253584 79354 253612 131174
rect 253676 119406 253704 157354
rect 254596 138786 254624 164290
rect 254584 138780 254636 138786
rect 254584 138722 254636 138728
rect 254584 134020 254636 134026
rect 254584 133962 254636 133968
rect 253664 119400 253716 119406
rect 253664 119342 253716 119348
rect 253572 79348 253624 79354
rect 253572 79290 253624 79296
rect 253480 47660 253532 47666
rect 253480 47602 253532 47608
rect 253388 22840 253440 22846
rect 253388 22782 253440 22788
rect 254596 19990 254624 133962
rect 254688 126954 254716 165650
rect 254952 156052 255004 156058
rect 254952 155994 255004 156000
rect 254860 146396 254912 146402
rect 254860 146338 254912 146344
rect 254676 126948 254728 126954
rect 254676 126890 254728 126896
rect 254768 125724 254820 125730
rect 254768 125666 254820 125672
rect 254676 117496 254728 117502
rect 254676 117438 254728 117444
rect 254688 35222 254716 117438
rect 254780 71058 254808 125666
rect 254872 106146 254900 146338
rect 254964 118046 254992 155994
rect 255964 153400 256016 153406
rect 255964 153342 256016 153348
rect 254952 118040 255004 118046
rect 254952 117982 255004 117988
rect 255976 111722 256004 153342
rect 256160 136542 256188 173946
rect 256240 171284 256292 171290
rect 256240 171226 256292 171232
rect 256148 136536 256200 136542
rect 256148 136478 256200 136484
rect 256056 135380 256108 135386
rect 256056 135322 256108 135328
rect 255964 111716 256016 111722
rect 255964 111658 256016 111664
rect 255964 107772 256016 107778
rect 255964 107714 256016 107720
rect 254860 106140 254912 106146
rect 254860 106082 254912 106088
rect 254860 99544 254912 99550
rect 254860 99486 254912 99492
rect 254872 75206 254900 99486
rect 254860 75200 254912 75206
rect 254860 75142 254912 75148
rect 254768 71052 254820 71058
rect 254768 70994 254820 71000
rect 254676 35216 254728 35222
rect 254676 35158 254728 35164
rect 254584 19984 254636 19990
rect 254584 19926 254636 19932
rect 255976 15978 256004 107714
rect 256068 44878 256096 135322
rect 256252 133890 256280 171226
rect 257528 168496 257580 168502
rect 257528 168438 257580 168444
rect 256424 161492 256476 161498
rect 256424 161434 256476 161440
rect 256332 145104 256384 145110
rect 256332 145046 256384 145052
rect 256240 133884 256292 133890
rect 256240 133826 256292 133832
rect 256240 129872 256292 129878
rect 256240 129814 256292 129820
rect 256148 123004 256200 123010
rect 256148 122946 256200 122952
rect 256160 55962 256188 122946
rect 256252 87650 256280 129814
rect 256344 105602 256372 145046
rect 256436 122126 256464 161434
rect 257344 151088 257396 151094
rect 257344 151030 257396 151036
rect 256424 122120 256476 122126
rect 256424 122062 256476 122068
rect 257356 111790 257384 151030
rect 257540 129742 257568 168438
rect 257712 160268 257764 160274
rect 257712 160210 257764 160216
rect 257620 132592 257672 132598
rect 257620 132534 257672 132540
rect 257528 129736 257580 129742
rect 257528 129678 257580 129684
rect 257436 128512 257488 128518
rect 257436 128454 257488 128460
rect 257344 111784 257396 111790
rect 257344 111726 257396 111732
rect 256424 110560 256476 110566
rect 256424 110502 256476 110508
rect 256332 105596 256384 105602
rect 256332 105538 256384 105544
rect 256332 96824 256384 96830
rect 256332 96766 256384 96772
rect 256240 87644 256292 87650
rect 256240 87586 256292 87592
rect 256344 64190 256372 96766
rect 256436 78062 256464 110502
rect 257344 102264 257396 102270
rect 257344 102206 257396 102212
rect 256424 78056 256476 78062
rect 256424 77998 256476 78004
rect 256332 64184 256384 64190
rect 256332 64126 256384 64132
rect 256148 55956 256200 55962
rect 256148 55898 256200 55904
rect 256056 44872 256108 44878
rect 256056 44814 256108 44820
rect 257356 28286 257384 102206
rect 257448 55894 257476 128454
rect 257528 123072 257580 123078
rect 257528 123014 257580 123020
rect 257436 55888 257488 55894
rect 257436 55830 257488 55836
rect 257540 54602 257568 123014
rect 257632 86358 257660 132534
rect 257724 123486 257752 160210
rect 258724 146464 258776 146470
rect 258724 146406 258776 146412
rect 257712 123480 257764 123486
rect 257712 123422 257764 123428
rect 257712 107840 257764 107846
rect 257712 107782 257764 107788
rect 257620 86352 257672 86358
rect 257620 86294 257672 86300
rect 257724 80782 257752 107782
rect 258736 106962 258764 146406
rect 258920 135250 258948 174014
rect 259092 168564 259144 168570
rect 259092 168506 259144 168512
rect 259000 139596 259052 139602
rect 259000 139538 259052 139544
rect 258908 135244 258960 135250
rect 258908 135186 258960 135192
rect 258816 134088 258868 134094
rect 258816 134030 258868 134036
rect 258724 106956 258776 106962
rect 258724 106898 258776 106904
rect 258724 103760 258776 103766
rect 258724 103702 258776 103708
rect 257712 80776 257764 80782
rect 257712 80718 257764 80724
rect 257528 54596 257580 54602
rect 257528 54538 257580 54544
rect 257344 28280 257396 28286
rect 257344 28222 257396 28228
rect 255964 15972 256016 15978
rect 255964 15914 256016 15920
rect 258736 14482 258764 103702
rect 258828 53106 258856 134030
rect 258908 120284 258960 120290
rect 258908 120226 258960 120232
rect 258920 57322 258948 120226
rect 259012 102134 259040 139538
rect 259104 131102 259132 168506
rect 260104 162988 260156 162994
rect 260104 162930 260156 162936
rect 259184 157480 259236 157486
rect 259184 157422 259236 157428
rect 259092 131096 259144 131102
rect 259092 131038 259144 131044
rect 259196 124982 259224 157422
rect 259184 124976 259236 124982
rect 259184 124918 259236 124924
rect 259092 124364 259144 124370
rect 259092 124306 259144 124312
rect 259000 102128 259052 102134
rect 259000 102070 259052 102076
rect 259104 90438 259132 124306
rect 260116 122670 260144 162930
rect 260104 122664 260156 122670
rect 260104 122606 260156 122612
rect 260104 116136 260156 116142
rect 260104 116078 260156 116084
rect 259276 106412 259328 106418
rect 259276 106354 259328 106360
rect 259184 100904 259236 100910
rect 259184 100846 259236 100852
rect 259092 90432 259144 90438
rect 259092 90374 259144 90380
rect 259196 68338 259224 100846
rect 259288 82210 259316 106354
rect 259276 82204 259328 82210
rect 259276 82146 259328 82152
rect 259184 68332 259236 68338
rect 259184 68274 259236 68280
rect 258908 57316 258960 57322
rect 258908 57258 258960 57264
rect 258816 53100 258868 53106
rect 258816 53042 258868 53048
rect 258724 14476 258776 14482
rect 258724 14418 258776 14424
rect 253204 9036 253256 9042
rect 253204 8978 253256 8984
rect 240784 7676 240836 7682
rect 240784 7618 240836 7624
rect 260116 6186 260144 116078
rect 260208 20670 260236 284543
rect 264426 174448 264482 174457
rect 264426 174383 264482 174392
rect 264440 173942 264468 174383
rect 264428 173936 264480 173942
rect 264428 173878 264480 173884
rect 263324 172916 263376 172922
rect 263324 172858 263376 172864
rect 263232 164416 263284 164422
rect 263232 164358 263284 164364
rect 260564 161764 260616 161770
rect 260564 161706 260616 161712
rect 260472 154760 260524 154766
rect 260472 154702 260524 154708
rect 260380 135448 260432 135454
rect 260380 135390 260432 135396
rect 260288 121508 260340 121514
rect 260288 121450 260340 121456
rect 260300 46238 260328 121450
rect 260392 69766 260420 135390
rect 260484 114510 260512 154702
rect 260576 122738 260604 161706
rect 262954 159896 263010 159905
rect 262954 159831 263010 159840
rect 261760 154692 261812 154698
rect 261760 154634 261812 154640
rect 261668 149252 261720 149258
rect 261668 149194 261720 149200
rect 261574 141944 261630 141953
rect 261574 141879 261630 141888
rect 261588 138718 261616 141879
rect 261576 138712 261628 138718
rect 261576 138654 261628 138660
rect 261576 132660 261628 132666
rect 261576 132602 261628 132608
rect 261484 124296 261536 124302
rect 261484 124238 261536 124244
rect 260564 122732 260616 122738
rect 260564 122674 260616 122680
rect 260472 114504 260524 114510
rect 260472 114446 260524 114452
rect 260472 110628 260524 110634
rect 260472 110570 260524 110576
rect 260484 76634 260512 110570
rect 260564 104916 260616 104922
rect 260564 104858 260616 104864
rect 260576 86290 260604 104858
rect 260564 86284 260616 86290
rect 260564 86226 260616 86232
rect 260472 76628 260524 76634
rect 260472 76570 260524 76576
rect 260380 69760 260432 69766
rect 260380 69702 260432 69708
rect 261496 51746 261524 124238
rect 261588 84930 261616 132602
rect 261680 109002 261708 149194
rect 261772 120766 261800 154634
rect 262864 149184 262916 149190
rect 262864 149126 262916 149132
rect 262586 135824 262642 135833
rect 262586 135759 262642 135768
rect 262600 135386 262628 135759
rect 262588 135380 262640 135386
rect 262588 135322 262640 135328
rect 261760 120760 261812 120766
rect 261760 120702 261812 120708
rect 261668 108996 261720 109002
rect 261668 108938 261720 108944
rect 262876 107642 262904 149126
rect 262968 122806 262996 159831
rect 263140 143676 263192 143682
rect 263140 143618 263192 143624
rect 263048 135312 263100 135318
rect 263048 135254 263100 135260
rect 262956 122800 263008 122806
rect 262956 122742 263008 122748
rect 262956 116000 263008 116006
rect 262956 115942 263008 115948
rect 262864 107636 262916 107642
rect 262864 107578 262916 107584
rect 261666 100600 261722 100609
rect 261666 100535 261722 100544
rect 261576 84924 261628 84930
rect 261576 84866 261628 84872
rect 261680 65550 261708 100535
rect 262864 98116 262916 98122
rect 262864 98058 262916 98064
rect 261668 65544 261720 65550
rect 261668 65486 261720 65492
rect 261484 51740 261536 51746
rect 261484 51682 261536 51688
rect 260288 46232 260340 46238
rect 260288 46174 260340 46180
rect 260196 20664 260248 20670
rect 260196 20606 260248 20612
rect 262876 10334 262904 98058
rect 262968 29646 262996 115942
rect 263060 75274 263088 135254
rect 263152 104174 263180 143618
rect 263244 126274 263272 164358
rect 263336 136610 263364 172858
rect 265254 172000 265310 172009
rect 265254 171935 265310 171944
rect 265268 171290 265296 171935
rect 265438 171592 265494 171601
rect 265438 171527 265494 171536
rect 265256 171284 265308 171290
rect 265256 171226 265308 171232
rect 265452 171222 265480 171527
rect 265440 171216 265492 171222
rect 265440 171158 265492 171164
rect 265530 171184 265586 171193
rect 265530 171119 265532 171128
rect 265584 171119 265586 171128
rect 265532 171090 265584 171096
rect 265530 170640 265586 170649
rect 265530 170575 265586 170584
rect 265162 170232 265218 170241
rect 265162 170167 265218 170176
rect 265176 169794 265204 170167
rect 265544 169862 265572 170575
rect 265532 169856 265584 169862
rect 265532 169798 265584 169804
rect 265164 169788 265216 169794
rect 265164 169730 265216 169736
rect 265346 167648 265402 167657
rect 265346 167583 265402 167592
rect 265162 167104 265218 167113
rect 265360 167074 265388 167583
rect 265162 167039 265218 167048
rect 265348 167068 265400 167074
rect 265176 166326 265204 167039
rect 265348 167010 265400 167016
rect 265164 166320 265216 166326
rect 265164 166262 265216 166268
rect 265438 166016 265494 166025
rect 265438 165951 265494 165960
rect 264426 165744 264482 165753
rect 265452 165714 265480 165951
rect 264426 165679 264482 165688
rect 265440 165708 265492 165714
rect 264242 140176 264298 140185
rect 264242 140111 264298 140120
rect 263324 136604 263376 136610
rect 263324 136546 263376 136552
rect 264152 127152 264204 127158
rect 264152 127094 264204 127100
rect 264164 126857 264192 127094
rect 264150 126848 264206 126857
rect 264150 126783 264206 126792
rect 263232 126268 263284 126274
rect 263232 126210 263284 126216
rect 263324 125656 263376 125662
rect 263324 125598 263376 125604
rect 263232 106344 263284 106350
rect 263232 106286 263284 106292
rect 263140 104168 263192 104174
rect 263140 104110 263192 104116
rect 263140 100836 263192 100842
rect 263140 100778 263192 100784
rect 263048 75268 263100 75274
rect 263048 75210 263100 75216
rect 263152 66910 263180 100778
rect 263244 83502 263272 106286
rect 263336 89078 263364 125598
rect 263416 103624 263468 103630
rect 263416 103566 263468 103572
rect 263324 89072 263376 89078
rect 263324 89014 263376 89020
rect 263428 89010 263456 103566
rect 263416 89004 263468 89010
rect 263416 88946 263468 88952
rect 263232 83496 263284 83502
rect 263232 83438 263284 83444
rect 263140 66904 263192 66910
rect 263140 66846 263192 66852
rect 262956 29640 263008 29646
rect 262956 29582 263008 29588
rect 262864 10328 262916 10334
rect 262864 10270 262916 10276
rect 264256 8974 264284 140111
rect 264334 130248 264390 130257
rect 264334 130183 264390 130192
rect 264348 39370 264376 130183
rect 264440 125594 264468 165679
rect 265440 165650 265492 165656
rect 265438 165064 265494 165073
rect 265438 164999 265494 165008
rect 265452 164286 265480 164999
rect 265440 164280 265492 164286
rect 265440 164222 265492 164228
rect 265162 163840 265218 163849
rect 265162 163775 265218 163784
rect 264702 163432 264758 163441
rect 264702 163367 264758 163376
rect 264612 159316 264664 159322
rect 264612 159258 264664 159264
rect 264520 153264 264572 153270
rect 264520 153206 264572 153212
rect 264532 153105 264560 153206
rect 264518 153096 264574 153105
rect 264518 153031 264574 153040
rect 264518 135960 264574 135969
rect 264518 135895 264574 135904
rect 264532 135454 264560 135895
rect 264520 135448 264572 135454
rect 264520 135390 264572 135396
rect 264520 134020 264572 134026
rect 264520 133962 264572 133968
rect 264532 133793 264560 133962
rect 264518 133784 264574 133793
rect 264518 133719 264574 133728
rect 264518 132016 264574 132025
rect 264518 131951 264574 131960
rect 264428 125588 264480 125594
rect 264428 125530 264480 125536
rect 264428 123072 264480 123078
rect 264428 123014 264480 123020
rect 264440 122641 264468 123014
rect 264426 122632 264482 122641
rect 264426 122567 264482 122576
rect 264426 122088 264482 122097
rect 264426 122023 264482 122032
rect 264440 49094 264468 122023
rect 264532 58682 264560 131951
rect 264624 121446 264652 159258
rect 264716 124914 264744 163367
rect 265176 163130 265204 163775
rect 265164 163124 265216 163130
rect 265164 163066 265216 163072
rect 265438 162072 265494 162081
rect 265438 162007 265494 162016
rect 265452 161770 265480 162007
rect 265440 161764 265492 161770
rect 265440 161706 265492 161712
rect 265532 160268 265584 160274
rect 265532 160210 265584 160216
rect 265544 160177 265572 160210
rect 265530 160168 265586 160177
rect 265530 160103 265586 160112
rect 265438 159080 265494 159089
rect 265438 159015 265494 159024
rect 265452 158846 265480 159015
rect 265440 158840 265492 158846
rect 265346 158808 265402 158817
rect 265440 158782 265492 158788
rect 265346 158743 265402 158752
rect 265360 158030 265388 158743
rect 265348 158024 265400 158030
rect 265348 157966 265400 157972
rect 265162 157856 265218 157865
rect 265162 157791 265218 157800
rect 265176 156670 265204 157791
rect 265164 156664 265216 156670
rect 265164 156606 265216 156612
rect 265438 155680 265494 155689
rect 265438 155615 265494 155624
rect 265452 154630 265480 155615
rect 265530 155272 265586 155281
rect 265530 155207 265586 155216
rect 265544 154698 265572 155207
rect 265532 154692 265584 154698
rect 265532 154634 265584 154640
rect 265440 154624 265492 154630
rect 265440 154566 265492 154572
rect 265530 153912 265586 153921
rect 265530 153847 265586 153856
rect 265544 153338 265572 153847
rect 265532 153332 265584 153338
rect 265532 153274 265584 153280
rect 265254 152688 265310 152697
rect 265254 152623 265310 152632
rect 265268 151910 265296 152623
rect 265256 151904 265308 151910
rect 265256 151846 265308 151852
rect 265346 150920 265402 150929
rect 265346 150855 265402 150864
rect 265360 150550 265388 150855
rect 265348 150544 265400 150550
rect 265070 150512 265126 150521
rect 265348 150486 265400 150492
rect 265070 150447 265072 150456
rect 265124 150447 265126 150456
rect 265072 150418 265124 150424
rect 265346 150104 265402 150113
rect 265346 150039 265402 150048
rect 265360 149258 265388 150039
rect 265530 149696 265586 149705
rect 265530 149631 265586 149640
rect 265348 149252 265400 149258
rect 265348 149194 265400 149200
rect 265544 149122 265572 149631
rect 265532 149116 265584 149122
rect 265532 149058 265584 149064
rect 265254 147928 265310 147937
rect 265254 147863 265310 147872
rect 265268 145586 265296 147863
rect 265530 147112 265586 147121
rect 265530 147047 265586 147056
rect 265544 146402 265572 147047
rect 265532 146396 265584 146402
rect 265532 146338 265584 146344
rect 265346 146160 265402 146169
rect 265346 146095 265402 146104
rect 265256 145580 265308 145586
rect 265256 145522 265308 145528
rect 265162 145344 265218 145353
rect 265162 145279 265218 145288
rect 265176 144974 265204 145279
rect 265164 144968 265216 144974
rect 265164 144910 265216 144916
rect 265360 144650 265388 146095
rect 265268 144622 265388 144650
rect 265268 144226 265296 144622
rect 265346 144528 265402 144537
rect 265346 144463 265402 144472
rect 265256 144220 265308 144226
rect 265256 144162 265308 144168
rect 265360 143614 265388 144463
rect 265348 143608 265400 143614
rect 265348 143550 265400 143556
rect 265530 143576 265586 143585
rect 265530 143511 265586 143520
rect 265162 143168 265218 143177
rect 265162 143103 265218 143112
rect 265176 142186 265204 143103
rect 265164 142180 265216 142186
rect 265164 142122 265216 142128
rect 265544 139602 265572 143511
rect 265532 139596 265584 139602
rect 265532 139538 265584 139544
rect 265438 138408 265494 138417
rect 265438 138343 265494 138352
rect 265452 138174 265480 138343
rect 265440 138168 265492 138174
rect 265440 138110 265492 138116
rect 265530 138136 265586 138145
rect 265530 138071 265532 138080
rect 265584 138071 265586 138080
rect 265532 138042 265584 138048
rect 265438 137592 265494 137601
rect 265438 137527 265494 137536
rect 265452 136678 265480 137527
rect 265530 137184 265586 137193
rect 265530 137119 265586 137128
rect 265544 136814 265572 137119
rect 265532 136808 265584 136814
rect 265532 136750 265584 136756
rect 265440 136672 265492 136678
rect 265440 136614 265492 136620
rect 265254 136368 265310 136377
rect 265254 136303 265310 136312
rect 265268 135522 265296 136303
rect 265256 135516 265308 135522
rect 265256 135458 265308 135464
rect 265254 134600 265310 134609
rect 265254 134535 265310 134544
rect 265268 133958 265296 134535
rect 265256 133952 265308 133958
rect 265256 133894 265308 133900
rect 265162 132832 265218 132841
rect 265162 132767 265218 132776
rect 265176 132666 265204 132767
rect 265164 132660 265216 132666
rect 265164 132602 265216 132608
rect 265530 129432 265586 129441
rect 265530 129367 265586 129376
rect 265346 129024 265402 129033
rect 265346 128959 265402 128968
rect 265360 128450 265388 128959
rect 265348 128444 265400 128450
rect 265348 128386 265400 128392
rect 265544 128382 265572 129367
rect 265532 128376 265584 128382
rect 265532 128318 265584 128324
rect 265530 127256 265586 127265
rect 265530 127191 265586 127200
rect 265544 127090 265572 127191
rect 265532 127084 265584 127090
rect 265532 127026 265584 127032
rect 265532 125724 265584 125730
rect 265532 125666 265584 125672
rect 265544 125633 265572 125666
rect 265530 125624 265586 125633
rect 265530 125559 265586 125568
rect 264704 124908 264756 124914
rect 264704 124850 264756 124856
rect 265162 124672 265218 124681
rect 265162 124607 265218 124616
rect 265176 124234 265204 124607
rect 265348 124296 265400 124302
rect 265346 124264 265348 124273
rect 265400 124264 265402 124273
rect 265164 124228 265216 124234
rect 265346 124199 265402 124208
rect 265164 124170 265216 124176
rect 265438 123448 265494 123457
rect 265438 123383 265494 123392
rect 265162 123040 265218 123049
rect 265162 122975 265164 122984
rect 265216 122975 265218 122984
rect 265164 122946 265216 122952
rect 265452 122874 265480 123383
rect 265440 122868 265492 122874
rect 265440 122810 265492 122816
rect 265530 121680 265586 121689
rect 264704 121644 264756 121650
rect 265530 121615 265586 121624
rect 264704 121586 264756 121592
rect 264612 121440 264664 121446
rect 264612 121382 264664 121388
rect 264716 121281 264744 121586
rect 265544 121514 265572 121615
rect 265532 121508 265584 121514
rect 265532 121450 265584 121456
rect 264702 121272 264758 121281
rect 264702 121207 264758 121216
rect 265530 120864 265586 120873
rect 265530 120799 265586 120808
rect 265544 120290 265572 120799
rect 265532 120284 265584 120290
rect 265532 120226 265584 120232
rect 265438 120184 265494 120193
rect 265438 120119 265440 120128
rect 265492 120119 265494 120128
rect 265440 120090 265492 120096
rect 265530 119096 265586 119105
rect 265530 119031 265586 119040
rect 265438 118824 265494 118833
rect 265438 118759 265440 118768
rect 265492 118759 265494 118768
rect 265440 118730 265492 118736
rect 265544 118726 265572 119031
rect 265532 118720 265584 118726
rect 265532 118662 265584 118668
rect 265530 118280 265586 118289
rect 265530 118215 265586 118224
rect 265440 118040 265492 118046
rect 265440 117982 265492 117988
rect 265348 117564 265400 117570
rect 265348 117506 265400 117512
rect 264612 116068 264664 116074
rect 264612 116010 264664 116016
rect 264624 115977 264652 116010
rect 264610 115968 264666 115977
rect 264610 115903 264666 115912
rect 265360 115258 265388 117506
rect 265452 116618 265480 117982
rect 265544 117502 265572 118215
rect 265532 117496 265584 117502
rect 265532 117438 265584 117444
rect 265440 116612 265492 116618
rect 265440 116554 265492 116560
rect 265348 115252 265400 115258
rect 265348 115194 265400 115200
rect 265530 112296 265586 112305
rect 265530 112231 265586 112240
rect 265544 111926 265572 112231
rect 265532 111920 265584 111926
rect 265532 111862 265584 111868
rect 265162 110936 265218 110945
rect 265162 110871 265218 110880
rect 265176 110634 265204 110871
rect 265164 110628 265216 110634
rect 265164 110570 265216 110576
rect 265346 109304 265402 109313
rect 265346 109239 265402 109248
rect 265360 109070 265388 109239
rect 265348 109064 265400 109070
rect 265348 109006 265400 109012
rect 264610 108760 264666 108769
rect 264610 108695 264666 108704
rect 264624 79422 264652 108695
rect 265530 108352 265586 108361
rect 265530 108287 265586 108296
rect 265544 107846 265572 108287
rect 265532 107840 265584 107846
rect 265532 107782 265584 107788
rect 265438 107128 265494 107137
rect 265438 107063 265494 107072
rect 265452 106418 265480 107063
rect 265440 106412 265492 106418
rect 265440 106354 265492 106360
rect 265438 105360 265494 105369
rect 265438 105295 265494 105304
rect 264794 104952 264850 104961
rect 265452 104922 265480 105295
rect 264794 104887 264850 104896
rect 265440 104916 265492 104922
rect 264702 103184 264758 103193
rect 264702 103119 264758 103128
rect 264716 84862 264744 103119
rect 264808 87718 264836 104887
rect 265440 104858 265492 104864
rect 265346 104544 265402 104553
rect 265346 104479 265402 104488
rect 265162 104000 265218 104009
rect 265162 103935 265218 103944
rect 265176 103766 265204 103935
rect 265164 103760 265216 103766
rect 265164 103702 265216 103708
rect 265360 103562 265388 104479
rect 265348 103556 265400 103562
rect 265348 103498 265400 103504
rect 265438 102776 265494 102785
rect 265438 102711 265494 102720
rect 265452 102406 265480 102711
rect 265440 102400 265492 102406
rect 265440 102342 265492 102348
rect 265530 101008 265586 101017
rect 265530 100943 265586 100952
rect 265544 100910 265572 100943
rect 265532 100904 265584 100910
rect 265532 100846 265584 100852
rect 265530 99512 265586 99521
rect 265530 99447 265532 99456
rect 265584 99447 265586 99456
rect 265532 99418 265584 99424
rect 265636 99374 265664 285874
rect 265714 285832 265770 285841
rect 265714 285767 265770 285776
rect 265452 99346 265664 99374
rect 265452 95130 265480 99346
rect 265728 98954 265756 285767
rect 267096 255332 267148 255338
rect 267096 255274 267148 255280
rect 267004 236768 267056 236774
rect 267004 236710 267056 236716
rect 265898 175400 265954 175409
rect 265898 175335 265954 175344
rect 265912 174554 265940 175335
rect 266082 174992 266138 175001
rect 266082 174927 266138 174936
rect 265990 174584 266046 174593
rect 265900 174548 265952 174554
rect 265990 174519 266046 174528
rect 265900 174490 265952 174496
rect 265806 174176 265862 174185
rect 265806 174111 265862 174120
rect 265820 174078 265848 174111
rect 265808 174072 265860 174078
rect 265808 174014 265860 174020
rect 266004 174010 266032 174519
rect 265992 174004 266044 174010
rect 265992 173946 266044 173952
rect 265990 173768 266046 173777
rect 265990 173703 266046 173712
rect 265898 173360 265954 173369
rect 265898 173295 265954 173304
rect 265806 172816 265862 172825
rect 265806 172751 265862 172760
rect 265820 172718 265848 172751
rect 265808 172712 265860 172718
rect 265808 172654 265860 172660
rect 265912 172582 265940 173295
rect 266004 172650 266032 173703
rect 266096 172922 266124 174927
rect 266084 172916 266136 172922
rect 266084 172858 266136 172864
rect 265992 172644 266044 172650
rect 265992 172586 266044 172592
rect 265900 172576 265952 172582
rect 265900 172518 265952 172524
rect 265808 169924 265860 169930
rect 265808 169866 265860 169872
rect 265820 169833 265848 169866
rect 265806 169824 265862 169833
rect 265806 169759 265862 169768
rect 265898 169416 265954 169425
rect 265898 169351 265954 169360
rect 265806 168600 265862 168609
rect 265912 168570 265940 169351
rect 265990 169008 266046 169017
rect 265990 168943 266046 168952
rect 265806 168535 265862 168544
rect 265900 168564 265952 168570
rect 265820 168502 265848 168535
rect 265900 168506 265952 168512
rect 265808 168496 265860 168502
rect 265808 168438 265860 168444
rect 265898 168464 265954 168473
rect 266004 168434 266032 168943
rect 265898 168399 265954 168408
rect 265992 168428 266044 168434
rect 265806 167240 265862 167249
rect 265806 167175 265862 167184
rect 265820 167142 265848 167175
rect 265808 167136 265860 167142
rect 265808 167078 265860 167084
rect 265912 166994 265940 168399
rect 265992 168370 266044 168376
rect 265912 166966 266124 166994
rect 265806 166424 265862 166433
rect 265806 166359 265862 166368
rect 265820 165782 265848 166359
rect 265808 165776 265860 165782
rect 265808 165718 265860 165724
rect 265898 164656 265954 164665
rect 265898 164591 265954 164600
rect 265808 164416 265860 164422
rect 265808 164358 265860 164364
rect 265820 164257 265848 164358
rect 265912 164354 265940 164591
rect 265900 164348 265952 164354
rect 265900 164290 265952 164296
rect 265806 164248 265862 164257
rect 265806 164183 265862 164192
rect 265806 163024 265862 163033
rect 265806 162959 265808 162968
rect 265860 162959 265862 162968
rect 265808 162930 265860 162936
rect 265806 161664 265862 161673
rect 265806 161599 265862 161608
rect 265820 161498 265848 161599
rect 265808 161492 265860 161498
rect 265808 161434 265860 161440
rect 265990 160848 266046 160857
rect 265990 160783 266046 160792
rect 265898 160440 265954 160449
rect 265898 160375 265954 160384
rect 265912 160138 265940 160375
rect 266004 160206 266032 160783
rect 265992 160200 266044 160206
rect 265992 160142 266044 160148
rect 265900 160132 265952 160138
rect 265900 160074 265952 160080
rect 265898 159488 265954 159497
rect 265898 159423 265954 159432
rect 265912 158778 265940 159423
rect 265900 158772 265952 158778
rect 265900 158714 265952 158720
rect 265898 158264 265954 158273
rect 265898 158199 265954 158208
rect 265912 157486 265940 158199
rect 266096 158098 266124 166966
rect 266266 161528 266322 161537
rect 266266 161463 266322 161472
rect 266280 159322 266308 161463
rect 266268 159316 266320 159322
rect 266268 159258 266320 159264
rect 266084 158092 266136 158098
rect 266084 158034 266136 158040
rect 265900 157480 265952 157486
rect 265806 157448 265862 157457
rect 265900 157422 265952 157428
rect 265806 157383 265808 157392
rect 265860 157383 265862 157392
rect 265808 157354 265860 157360
rect 265898 156904 265954 156913
rect 265898 156839 265954 156848
rect 265806 156496 265862 156505
rect 265806 156431 265862 156440
rect 265820 155990 265848 156431
rect 265912 156058 265940 156839
rect 266082 156088 266138 156097
rect 265900 156052 265952 156058
rect 266082 156023 266138 156032
rect 265900 155994 265952 156000
rect 265808 155984 265860 155990
rect 265808 155926 265860 155932
rect 265806 154864 265862 154873
rect 265806 154799 265862 154808
rect 265820 154766 265848 154799
rect 265808 154760 265860 154766
rect 265808 154702 265860 154708
rect 265990 154728 266046 154737
rect 265990 154663 266046 154672
rect 265806 153504 265862 153513
rect 265806 153439 265862 153448
rect 265820 153406 265848 153439
rect 265808 153400 265860 153406
rect 265808 153342 265860 153348
rect 265898 152144 265954 152153
rect 265898 152079 265954 152088
rect 265806 151872 265862 151881
rect 265806 151807 265808 151816
rect 265860 151807 265862 151816
rect 265808 151778 265860 151784
rect 265806 151328 265862 151337
rect 265806 151263 265862 151272
rect 265820 150618 265848 151263
rect 265912 151094 265940 152079
rect 265900 151088 265952 151094
rect 265900 151030 265952 151036
rect 265808 150612 265860 150618
rect 265808 150554 265860 150560
rect 265806 149288 265862 149297
rect 265806 149223 265862 149232
rect 265820 149190 265848 149223
rect 265808 149184 265860 149190
rect 265808 149126 265860 149132
rect 266004 149002 266032 154663
rect 265820 148974 266032 149002
rect 265820 146946 265848 148974
rect 266096 148866 266124 156023
rect 266004 148838 266124 148866
rect 265898 148336 265954 148345
rect 265898 148271 265954 148280
rect 265912 147694 265940 148271
rect 265900 147688 265952 147694
rect 265900 147630 265952 147636
rect 265808 146940 265860 146946
rect 265808 146882 265860 146888
rect 265898 146704 265954 146713
rect 265898 146639 265954 146648
rect 265806 146568 265862 146577
rect 265806 146503 265862 146512
rect 265820 146470 265848 146503
rect 265808 146464 265860 146470
rect 265808 146406 265860 146412
rect 265912 146334 265940 146639
rect 265900 146328 265952 146334
rect 265900 146270 265952 146276
rect 265898 145752 265954 145761
rect 265898 145687 265954 145696
rect 265808 145104 265860 145110
rect 265808 145046 265860 145052
rect 265820 144945 265848 145046
rect 265912 145042 265940 145687
rect 265900 145036 265952 145042
rect 265900 144978 265952 144984
rect 265806 144936 265862 144945
rect 265806 144871 265862 144880
rect 265806 144120 265862 144129
rect 265806 144055 265862 144064
rect 265820 143682 265848 144055
rect 265808 143676 265860 143682
rect 265808 143618 265860 143624
rect 266004 142882 266032 148838
rect 266082 148744 266138 148753
rect 266082 148679 266138 148688
rect 266096 147762 266124 148679
rect 266084 147756 266136 147762
rect 266084 147698 266136 147704
rect 266004 142854 266308 142882
rect 266174 142760 266230 142769
rect 266174 142695 266230 142704
rect 266082 142352 266138 142361
rect 266082 142287 266138 142296
rect 265806 141400 265862 141409
rect 265806 141335 265862 141344
rect 265820 140894 265848 141335
rect 265898 140992 265954 141001
rect 265898 140927 265954 140936
rect 265808 140888 265860 140894
rect 265808 140830 265860 140836
rect 265912 140826 265940 140927
rect 265990 140856 266046 140865
rect 265900 140820 265952 140826
rect 265990 140791 266046 140800
rect 265900 140762 265952 140768
rect 265898 139768 265954 139777
rect 265898 139703 265954 139712
rect 265912 139534 265940 139703
rect 265900 139528 265952 139534
rect 265806 139496 265862 139505
rect 265900 139470 265952 139476
rect 265806 139431 265808 139440
rect 265860 139431 265862 139440
rect 265808 139402 265860 139408
rect 266004 139346 266032 140791
rect 265820 139318 266032 139346
rect 266096 139346 266124 142287
rect 266188 139466 266216 142695
rect 266280 140078 266308 142854
rect 266268 140072 266320 140078
rect 266268 140014 266320 140020
rect 266176 139460 266228 139466
rect 266176 139402 266228 139408
rect 266096 139318 266308 139346
rect 265820 117570 265848 139318
rect 265900 139256 265952 139262
rect 265900 139198 265952 139204
rect 265912 118046 265940 139198
rect 265990 138816 266046 138825
rect 265990 138751 266046 138760
rect 266004 138038 266032 138751
rect 265992 138032 266044 138038
rect 266280 138014 266308 139318
rect 265992 137974 266044 137980
rect 266096 137986 266308 138014
rect 265990 136776 266046 136785
rect 265990 136711 265992 136720
rect 266044 136711 266046 136720
rect 265992 136682 266044 136688
rect 265990 135416 266046 135425
rect 265990 135351 266046 135360
rect 266004 135318 266032 135351
rect 265992 135312 266044 135318
rect 265992 135254 266044 135260
rect 265990 134192 266046 134201
rect 265990 134127 266046 134136
rect 266004 134094 266032 134127
rect 265992 134088 266044 134094
rect 265992 134030 266044 134036
rect 265992 132592 266044 132598
rect 265990 132560 265992 132569
rect 266044 132560 266046 132569
rect 265990 132495 266046 132504
rect 265990 131608 266046 131617
rect 265990 131543 266046 131552
rect 266004 131306 266032 131543
rect 265992 131300 266044 131306
rect 265992 131242 266044 131248
rect 265992 129940 266044 129946
rect 265992 129882 266044 129888
rect 266004 129849 266032 129882
rect 265990 129840 266046 129849
rect 265990 129775 266046 129784
rect 265990 128616 266046 128625
rect 265990 128551 266046 128560
rect 266004 128518 266032 128551
rect 265992 128512 266044 128518
rect 265992 128454 266044 128460
rect 265992 128376 266044 128382
rect 265992 128318 266044 128324
rect 265900 118040 265952 118046
rect 265900 117982 265952 117988
rect 265898 117872 265954 117881
rect 265898 117807 265954 117816
rect 265808 117564 265860 117570
rect 265808 117506 265860 117512
rect 265806 117464 265862 117473
rect 265912 117434 265940 117807
rect 265806 117399 265862 117408
rect 265900 117428 265952 117434
rect 265820 117366 265848 117399
rect 265900 117370 265952 117376
rect 265808 117360 265860 117366
rect 265808 117302 265860 117308
rect 265898 116512 265954 116521
rect 265898 116447 265954 116456
rect 265912 116210 265940 116447
rect 265900 116204 265952 116210
rect 265900 116146 265952 116152
rect 265808 116136 265860 116142
rect 265806 116104 265808 116113
rect 265860 116104 265862 116113
rect 265806 116039 265862 116048
rect 265898 115288 265954 115297
rect 265898 115223 265954 115232
rect 265806 114744 265862 114753
rect 265806 114679 265862 114688
rect 265820 114646 265848 114679
rect 265808 114640 265860 114646
rect 265808 114582 265860 114588
rect 265912 114578 265940 115223
rect 265900 114572 265952 114578
rect 265900 114514 265952 114520
rect 265898 113928 265954 113937
rect 265898 113863 265954 113872
rect 265806 113520 265862 113529
rect 265806 113455 265862 113464
rect 265820 113354 265848 113455
rect 265808 113348 265860 113354
rect 265808 113290 265860 113296
rect 265912 113286 265940 113863
rect 265900 113280 265952 113286
rect 265806 113248 265862 113257
rect 265900 113222 265952 113228
rect 265806 113183 265808 113192
rect 265860 113183 265862 113192
rect 265808 113154 265860 113160
rect 265898 112704 265954 112713
rect 265898 112639 265954 112648
rect 265806 112160 265862 112169
rect 265806 112095 265862 112104
rect 265820 111994 265848 112095
rect 265808 111988 265860 111994
rect 265808 111930 265860 111936
rect 265912 111858 265940 112639
rect 265900 111852 265952 111858
rect 265900 111794 265952 111800
rect 265898 111344 265954 111353
rect 265898 111279 265954 111288
rect 265808 110560 265860 110566
rect 265806 110528 265808 110537
rect 265860 110528 265862 110537
rect 265912 110498 265940 111279
rect 265806 110463 265862 110472
rect 265900 110492 265952 110498
rect 265900 110434 265952 110440
rect 265898 110120 265954 110129
rect 265898 110055 265954 110064
rect 265806 109712 265862 109721
rect 265806 109647 265862 109656
rect 265820 109206 265848 109647
rect 265808 109200 265860 109206
rect 265808 109142 265860 109148
rect 265912 109138 265940 110055
rect 265900 109132 265952 109138
rect 265900 109074 265952 109080
rect 265806 107944 265862 107953
rect 265806 107879 265808 107888
rect 265860 107879 265862 107888
rect 265808 107850 265860 107856
rect 265808 107772 265860 107778
rect 265808 107714 265860 107720
rect 265820 107681 265848 107714
rect 265806 107672 265862 107681
rect 265806 107607 265862 107616
rect 265806 106720 265862 106729
rect 265806 106655 265862 106664
rect 265820 106486 265848 106655
rect 265898 106584 265954 106593
rect 265898 106519 265954 106528
rect 265808 106480 265860 106486
rect 265808 106422 265860 106428
rect 265912 106350 265940 106519
rect 265900 106344 265952 106350
rect 265900 106286 265952 106292
rect 265806 105768 265862 105777
rect 265806 105703 265862 105712
rect 265820 105058 265848 105703
rect 265808 105052 265860 105058
rect 265808 104994 265860 105000
rect 265808 103624 265860 103630
rect 265806 103592 265808 103601
rect 265860 103592 265862 103601
rect 265806 103527 265862 103536
rect 265806 102368 265862 102377
rect 265806 102303 265862 102312
rect 265820 102270 265848 102303
rect 265808 102264 265860 102270
rect 265808 102206 265860 102212
rect 265898 101416 265954 101425
rect 265898 101351 265954 101360
rect 265806 100872 265862 100881
rect 265912 100842 265940 101351
rect 265806 100807 265862 100816
rect 265900 100836 265952 100842
rect 265820 100774 265848 100807
rect 265900 100778 265952 100784
rect 265808 100768 265860 100774
rect 265808 100710 265860 100716
rect 265898 100192 265954 100201
rect 265898 100127 265954 100136
rect 265806 99784 265862 99793
rect 265806 99719 265862 99728
rect 265820 99550 265848 99719
rect 265808 99544 265860 99550
rect 265808 99486 265860 99492
rect 265912 99414 265940 100127
rect 265900 99408 265952 99414
rect 265900 99350 265952 99356
rect 265636 98926 265756 98954
rect 265636 98002 265664 98926
rect 265714 98832 265770 98841
rect 265714 98767 265770 98776
rect 265728 98122 265756 98767
rect 266004 98546 266032 128318
rect 266096 117978 266124 137986
rect 266174 133240 266230 133249
rect 266174 133175 266230 133184
rect 266188 132530 266216 133175
rect 266176 132524 266228 132530
rect 266176 132466 266228 132472
rect 266176 131232 266228 131238
rect 266174 131200 266176 131209
rect 266228 131200 266230 131209
rect 266174 131135 266230 131144
rect 266174 130656 266230 130665
rect 266174 130591 266230 130600
rect 266188 129878 266216 130591
rect 266176 129872 266228 129878
rect 266176 129814 266228 129820
rect 266174 128480 266230 128489
rect 266174 128415 266230 128424
rect 266188 128382 266216 128415
rect 266176 128376 266228 128382
rect 266176 128318 266228 128324
rect 266174 127664 266230 127673
rect 266174 127599 266230 127608
rect 266188 127022 266216 127599
rect 266176 127016 266228 127022
rect 266176 126958 266228 126964
rect 266174 126440 266230 126449
rect 266174 126375 266230 126384
rect 266188 125798 266216 126375
rect 266266 126032 266322 126041
rect 266266 125967 266322 125976
rect 266176 125792 266228 125798
rect 266176 125734 266228 125740
rect 266280 125662 266308 125967
rect 266268 125656 266320 125662
rect 266268 125598 266320 125604
rect 266174 125080 266230 125089
rect 266174 125015 266230 125024
rect 266188 124370 266216 125015
rect 266176 124364 266228 124370
rect 266176 124306 266228 124312
rect 266174 123856 266230 123865
rect 266174 123791 266230 123800
rect 266188 122942 266216 123791
rect 266176 122936 266228 122942
rect 266176 122878 266228 122884
rect 266174 120456 266230 120465
rect 266174 120391 266230 120400
rect 266188 120222 266216 120391
rect 266176 120216 266228 120222
rect 266176 120158 266228 120164
rect 266174 119504 266230 119513
rect 266174 119439 266230 119448
rect 266188 118862 266216 119439
rect 266176 118856 266228 118862
rect 266176 118798 266228 118804
rect 266084 117972 266136 117978
rect 266084 117914 266136 117920
rect 266082 116920 266138 116929
rect 266082 116855 266138 116864
rect 266096 116006 266124 116855
rect 266084 116000 266136 116006
rect 266084 115942 266136 115948
rect 266082 114880 266138 114889
rect 266082 114815 266138 114824
rect 266096 98666 266124 114815
rect 266084 98660 266136 98666
rect 266084 98602 266136 98608
rect 266004 98518 266124 98546
rect 265990 98424 266046 98433
rect 265990 98359 266046 98368
rect 265716 98116 265768 98122
rect 265716 98058 265768 98064
rect 265808 98048 265860 98054
rect 265806 98016 265808 98025
rect 265860 98016 265862 98025
rect 265636 97974 265756 98002
rect 265622 97200 265678 97209
rect 265622 97135 265678 97144
rect 265532 96824 265584 96830
rect 265530 96792 265532 96801
rect 265584 96792 265586 96801
rect 265636 96762 265664 97135
rect 265530 96727 265586 96736
rect 265624 96756 265676 96762
rect 265624 96698 265676 96704
rect 265728 96286 265756 97974
rect 265806 97951 265862 97960
rect 265898 97608 265954 97617
rect 265898 97543 265954 97552
rect 265806 96928 265862 96937
rect 265806 96863 265862 96872
rect 265716 96280 265768 96286
rect 265716 96222 265768 96228
rect 265714 95704 265770 95713
rect 265714 95639 265770 95648
rect 265728 95266 265756 95639
rect 265716 95260 265768 95266
rect 265716 95202 265768 95208
rect 265440 95124 265492 95130
rect 265440 95066 265492 95072
rect 264796 87712 264848 87718
rect 264796 87654 264848 87660
rect 264704 84856 264756 84862
rect 264704 84798 264756 84804
rect 264612 79416 264664 79422
rect 264612 79358 264664 79364
rect 264520 58676 264572 58682
rect 264520 58618 264572 58624
rect 264428 49088 264480 49094
rect 264428 49030 264480 49036
rect 264336 39364 264388 39370
rect 264336 39306 264388 39312
rect 264244 8968 264296 8974
rect 264244 8910 264296 8916
rect 260104 6180 260156 6186
rect 260104 6122 260156 6128
rect 265820 4826 265848 96863
rect 265912 96694 265940 97543
rect 265900 96688 265952 96694
rect 265900 96630 265952 96636
rect 266004 89714 266032 98359
rect 266096 91798 266124 98518
rect 266084 91792 266136 91798
rect 266084 91734 266136 91740
rect 265912 89686 266032 89714
rect 265912 60042 265940 89686
rect 265900 60036 265952 60042
rect 265900 59978 265952 59984
rect 267016 6866 267044 236710
rect 267108 96150 267136 255274
rect 278056 175846 278084 286146
rect 280804 286000 280856 286006
rect 280804 285942 280856 285948
rect 280160 245676 280212 245682
rect 280160 245618 280212 245624
rect 279148 180396 279200 180402
rect 279148 180338 279200 180344
rect 278780 176656 278832 176662
rect 278780 176598 278832 176604
rect 278792 176089 278820 176598
rect 278778 176080 278834 176089
rect 278778 176015 278834 176024
rect 278044 175840 278096 175846
rect 278044 175782 278096 175788
rect 279160 171134 279188 180338
rect 279160 171106 279372 171134
rect 279344 149841 279372 171106
rect 279330 149832 279386 149841
rect 279330 149767 279386 149776
rect 280172 125497 280200 245618
rect 280344 181552 280396 181558
rect 280344 181494 280396 181500
rect 280250 180432 280306 180441
rect 280250 180367 280306 180376
rect 280158 125488 280214 125497
rect 280158 125423 280214 125432
rect 280264 106321 280292 180367
rect 280356 120873 280384 181494
rect 280528 178832 280580 178838
rect 280528 178774 280580 178780
rect 280436 175908 280488 175914
rect 280436 175850 280488 175856
rect 280448 121689 280476 175850
rect 280434 121680 280490 121689
rect 280434 121615 280490 121624
rect 280342 120864 280398 120873
rect 280342 120799 280398 120808
rect 280540 119377 280568 178774
rect 280712 176112 280764 176118
rect 280712 176054 280764 176060
rect 280620 176044 280672 176050
rect 280620 175986 280672 175992
rect 280632 141681 280660 175986
rect 280724 160177 280752 176054
rect 280816 162858 280844 285942
rect 280908 167618 280936 286554
rect 283196 286476 283248 286482
rect 283196 286418 283248 286424
rect 283104 284708 283156 284714
rect 283104 284650 283156 284656
rect 282184 283892 282236 283898
rect 282184 283834 282236 283840
rect 280988 252612 281040 252618
rect 280988 252554 281040 252560
rect 280896 167612 280948 167618
rect 280896 167554 280948 167560
rect 280804 162852 280856 162858
rect 280804 162794 280856 162800
rect 280710 160168 280766 160177
rect 280710 160103 280766 160112
rect 280618 141672 280674 141681
rect 280618 141607 280674 141616
rect 281000 136610 281028 252554
rect 281724 239488 281776 239494
rect 281724 239430 281776 239436
rect 281080 182980 281132 182986
rect 281080 182922 281132 182928
rect 281092 175914 281120 182922
rect 281540 177472 281592 177478
rect 281540 177414 281592 177420
rect 281080 175908 281132 175914
rect 281080 175850 281132 175856
rect 281552 172417 281580 177414
rect 281632 177404 281684 177410
rect 281632 177346 281684 177352
rect 281538 172408 281594 172417
rect 281538 172343 281594 172352
rect 281644 170105 281672 177346
rect 281630 170096 281686 170105
rect 281630 170031 281686 170040
rect 281736 168609 281764 239430
rect 281816 235272 281868 235278
rect 281816 235214 281868 235220
rect 281722 168600 281778 168609
rect 281722 168535 281778 168544
rect 281828 167793 281856 235214
rect 282000 184340 282052 184346
rect 282000 184282 282052 184288
rect 281906 181520 281962 181529
rect 281906 181455 281962 181464
rect 281814 167784 281870 167793
rect 281814 167719 281870 167728
rect 281540 162852 281592 162858
rect 281540 162794 281592 162800
rect 280988 136604 281040 136610
rect 280988 136546 281040 136552
rect 281552 122505 281580 162794
rect 281920 161474 281948 181455
rect 282012 164801 282040 184282
rect 282092 175840 282144 175846
rect 282092 175782 282144 175788
rect 281998 164792 282054 164801
rect 281998 164727 282054 164736
rect 282104 162489 282132 175782
rect 282196 170921 282224 283834
rect 282368 283620 282420 283626
rect 282368 283562 282420 283568
rect 282274 177440 282330 177449
rect 282274 177375 282330 177384
rect 282182 170912 282238 170921
rect 282182 170847 282238 170856
rect 282288 167113 282316 177375
rect 282380 173233 282408 283562
rect 282920 180124 282972 180130
rect 282920 180066 282972 180072
rect 282366 173224 282422 173233
rect 282366 173159 282422 173168
rect 282552 167612 282604 167618
rect 282552 167554 282604 167560
rect 282274 167104 282330 167113
rect 282274 167039 282330 167048
rect 282090 162480 282146 162489
rect 282090 162415 282146 162424
rect 281828 161446 281948 161474
rect 281828 154737 281856 161446
rect 282184 161220 282236 161226
rect 282184 161162 282236 161168
rect 282196 160857 282224 161162
rect 282182 160848 282238 160857
rect 282182 160783 282238 160792
rect 281906 158536 281962 158545
rect 281906 158471 281962 158480
rect 281920 157894 281948 158471
rect 282000 157956 282052 157962
rect 282000 157898 282052 157904
rect 281908 157888 281960 157894
rect 282012 157865 282040 157898
rect 281908 157830 281960 157836
rect 281998 157856 282054 157865
rect 281998 157791 282054 157800
rect 282460 156596 282512 156602
rect 282460 156538 282512 156544
rect 282472 156369 282500 156538
rect 282458 156360 282514 156369
rect 282458 156295 282514 156304
rect 282184 155780 282236 155786
rect 282184 155722 282236 155728
rect 281814 154728 281870 154737
rect 281814 154663 281870 154672
rect 282092 154148 282144 154154
rect 282092 154090 282144 154096
rect 282104 154057 282132 154090
rect 282090 154048 282146 154057
rect 282090 153983 282146 153992
rect 282092 153196 282144 153202
rect 282092 153138 282144 153144
rect 282104 152425 282132 153138
rect 282090 152416 282146 152425
rect 282090 152351 282146 152360
rect 281632 151020 281684 151026
rect 281632 150962 281684 150968
rect 281644 150929 281672 150962
rect 281630 150920 281686 150929
rect 281630 150855 281686 150864
rect 281722 150512 281778 150521
rect 281722 150447 281778 150456
rect 281632 137896 281684 137902
rect 281630 137864 281632 137873
rect 281684 137864 281686 137873
rect 281630 137799 281686 137808
rect 281632 136604 281684 136610
rect 281632 136546 281684 136552
rect 281644 123185 281672 136546
rect 281630 123176 281686 123185
rect 281630 123111 281686 123120
rect 281538 122496 281594 122505
rect 281538 122431 281594 122440
rect 281736 120193 281764 150447
rect 282092 148912 282144 148918
rect 282092 148854 282144 148860
rect 282104 147801 282132 148854
rect 282090 147792 282146 147801
rect 282090 147727 282146 147736
rect 281908 144492 281960 144498
rect 281908 144434 281960 144440
rect 281920 143993 281948 144434
rect 281906 143984 281962 143993
rect 281906 143919 281962 143928
rect 282196 135561 282224 155722
rect 282276 153332 282328 153338
rect 282276 153274 282328 153280
rect 282288 153241 282316 153274
rect 282274 153232 282330 153241
rect 282274 153167 282330 153176
rect 282276 151768 282328 151774
rect 282274 151736 282276 151745
rect 282328 151736 282330 151745
rect 282274 151671 282330 151680
rect 282276 137964 282328 137970
rect 282276 137906 282328 137912
rect 282288 137057 282316 137906
rect 282274 137048 282330 137057
rect 282274 136983 282330 136992
rect 282182 135552 282238 135561
rect 282182 135487 282238 135496
rect 281816 135176 281868 135182
rect 281816 135118 281868 135124
rect 281828 134065 281856 135118
rect 282564 134745 282592 167554
rect 282826 165472 282882 165481
rect 282932 165458 282960 180066
rect 283012 177812 283064 177818
rect 283012 177754 283064 177760
rect 282882 165430 282960 165458
rect 282826 165407 282882 165416
rect 282826 161664 282882 161673
rect 283024 161650 283052 177754
rect 282882 161622 283052 161650
rect 282826 161599 282882 161608
rect 282826 159352 282882 159361
rect 282826 159287 282882 159296
rect 282840 159186 282868 159287
rect 282828 159180 282880 159186
rect 282828 159122 282880 159128
rect 282828 157344 282880 157350
rect 282828 157286 282880 157292
rect 282840 157049 282868 157286
rect 282826 157040 282882 157049
rect 282826 156975 282882 156984
rect 282828 155916 282880 155922
rect 282828 155858 282880 155864
rect 282840 155553 282868 155858
rect 282826 155544 282882 155553
rect 282826 155479 282882 155488
rect 282826 150104 282882 150113
rect 282826 150039 282882 150048
rect 282840 149258 282868 150039
rect 282828 149252 282880 149258
rect 282828 149194 282880 149200
rect 282828 149048 282880 149054
rect 282828 148990 282880 148996
rect 282840 148617 282868 148990
rect 282826 148608 282882 148617
rect 282826 148543 282882 148552
rect 282826 146296 282882 146305
rect 282826 146231 282882 146240
rect 282840 145110 282868 146231
rect 282828 145104 282880 145110
rect 282828 145046 282880 145052
rect 282828 143540 282880 143546
rect 282828 143482 282880 143488
rect 282840 142497 282868 143482
rect 282826 142488 282882 142497
rect 282826 142423 282882 142432
rect 283116 142154 283144 284650
rect 283208 155786 283236 286418
rect 283656 286408 283708 286414
rect 283656 286350 283708 286356
rect 283288 181620 283340 181626
rect 283288 181562 283340 181568
rect 283196 155780 283248 155786
rect 283196 155722 283248 155728
rect 282932 142126 283144 142154
rect 282826 140176 282882 140185
rect 282826 140111 282882 140120
rect 282840 139874 282868 140111
rect 282828 139868 282880 139874
rect 282828 139810 282880 139816
rect 282932 139482 282960 142126
rect 282748 139454 282960 139482
rect 282748 139369 282776 139454
rect 282828 139392 282880 139398
rect 282734 139360 282790 139369
rect 282828 139334 282880 139340
rect 282734 139295 282790 139304
rect 282840 138553 282868 139334
rect 282826 138544 282882 138553
rect 282826 138479 282882 138488
rect 282828 136604 282880 136610
rect 282828 136546 282880 136552
rect 282840 136377 282868 136546
rect 282826 136368 282882 136377
rect 282826 136303 282882 136312
rect 282550 134736 282606 134745
rect 282550 134671 282606 134680
rect 281814 134056 281870 134065
rect 281814 133991 281870 134000
rect 282276 133884 282328 133890
rect 282276 133826 282328 133832
rect 282288 133249 282316 133826
rect 282274 133240 282330 133249
rect 282274 133175 282330 133184
rect 282092 132456 282144 132462
rect 282092 132398 282144 132404
rect 282550 132424 282606 132433
rect 282104 131753 282132 132398
rect 282550 132359 282552 132368
rect 282604 132359 282606 132368
rect 282552 132330 282604 132336
rect 282090 131744 282146 131753
rect 282090 131679 282146 131688
rect 281908 131096 281960 131102
rect 281908 131038 281960 131044
rect 281920 130937 281948 131038
rect 282092 131028 282144 131034
rect 282092 130970 282144 130976
rect 281906 130928 281962 130937
rect 281906 130863 281962 130872
rect 282104 130121 282132 130970
rect 282090 130112 282146 130121
rect 282090 130047 282146 130056
rect 282092 129668 282144 129674
rect 282092 129610 282144 129616
rect 281908 129600 281960 129606
rect 281908 129542 281960 129548
rect 281920 129441 281948 129542
rect 281906 129432 281962 129441
rect 281906 129367 281962 129376
rect 282104 128625 282132 129610
rect 282090 128616 282146 128625
rect 282090 128551 282146 128560
rect 281908 128240 281960 128246
rect 281908 128182 281960 128188
rect 281920 127809 281948 128182
rect 281906 127800 281962 127809
rect 281906 127735 281962 127744
rect 281908 127696 281960 127702
rect 281908 127638 281960 127644
rect 281920 127129 281948 127638
rect 281906 127120 281962 127129
rect 281906 127055 281962 127064
rect 282828 126744 282880 126750
rect 282828 126686 282880 126692
rect 282840 126313 282868 126686
rect 282826 126304 282882 126313
rect 282826 126239 282882 126248
rect 282826 124808 282882 124817
rect 282826 124743 282882 124752
rect 282840 124506 282868 124743
rect 282828 124500 282880 124506
rect 282828 124442 282880 124448
rect 282826 123992 282882 124001
rect 282826 123927 282882 123936
rect 282840 123554 282868 123927
rect 282828 123548 282880 123554
rect 282828 123490 282880 123496
rect 281722 120184 281778 120193
rect 281722 120119 281778 120128
rect 280526 119368 280582 119377
rect 280526 119303 280582 119312
rect 282828 118652 282880 118658
rect 282828 118594 282880 118600
rect 282736 118584 282788 118590
rect 282734 118552 282736 118561
rect 282788 118552 282790 118561
rect 282734 118487 282790 118496
rect 282840 117881 282868 118594
rect 282826 117872 282882 117881
rect 282826 117807 282882 117816
rect 282828 117292 282880 117298
rect 282828 117234 282880 117240
rect 282840 117065 282868 117234
rect 282826 117056 282882 117065
rect 282826 116991 282882 117000
rect 282828 116476 282880 116482
rect 282828 116418 282880 116424
rect 282840 116385 282868 116418
rect 282826 116376 282882 116385
rect 282826 116311 282882 116320
rect 282828 114844 282880 114850
rect 282828 114786 282880 114792
rect 282840 114753 282868 114786
rect 282826 114744 282882 114753
rect 282826 114679 282882 114688
rect 282736 114368 282788 114374
rect 282736 114310 282788 114316
rect 282748 114073 282776 114310
rect 282734 114064 282790 114073
rect 282734 113999 282790 114008
rect 282828 113484 282880 113490
rect 282828 113426 282880 113432
rect 282840 113257 282868 113426
rect 282826 113248 282882 113257
rect 282826 113183 282882 113192
rect 282828 112736 282880 112742
rect 282828 112678 282880 112684
rect 282840 112441 282868 112678
rect 282826 112432 282882 112441
rect 282826 112367 282882 112376
rect 281998 111752 282054 111761
rect 281998 111687 282054 111696
rect 282012 111110 282040 111687
rect 282828 111172 282880 111178
rect 282828 111114 282880 111120
rect 282000 111104 282052 111110
rect 282000 111046 282052 111052
rect 282840 110945 282868 111114
rect 282826 110936 282882 110945
rect 282826 110871 282882 110880
rect 282274 110120 282330 110129
rect 282274 110055 282330 110064
rect 282828 110084 282880 110090
rect 282288 109954 282316 110055
rect 282828 110026 282880 110032
rect 282276 109948 282328 109954
rect 282276 109890 282328 109896
rect 282840 109449 282868 110026
rect 282826 109440 282882 109449
rect 282826 109375 282882 109384
rect 282368 108996 282420 109002
rect 282368 108938 282420 108944
rect 281540 108656 281592 108662
rect 281538 108624 281540 108633
rect 281592 108624 281594 108633
rect 281538 108559 281594 108568
rect 282380 107817 282408 108938
rect 282366 107808 282422 107817
rect 282366 107743 282422 107752
rect 281724 107636 281776 107642
rect 281724 107578 281776 107584
rect 281736 107137 281764 107578
rect 281722 107128 281778 107137
rect 281722 107063 281778 107072
rect 280250 106312 280306 106321
rect 280250 106247 280306 106256
rect 282826 105496 282882 105505
rect 282826 105431 282882 105440
rect 282840 105126 282868 105431
rect 282828 105120 282880 105126
rect 282828 105062 282880 105068
rect 281540 104848 281592 104854
rect 281538 104816 281540 104825
rect 281592 104816 281594 104825
rect 281538 104751 281594 104760
rect 283300 104582 283328 181562
rect 283380 178764 283432 178770
rect 283380 178706 283432 178712
rect 283392 108662 283420 178706
rect 283564 178696 283616 178702
rect 283564 178638 283616 178644
rect 283472 177880 283524 177886
rect 283472 177822 283524 177828
rect 283484 137902 283512 177822
rect 283576 151026 283604 178638
rect 283564 151020 283616 151026
rect 283564 150962 283616 150968
rect 283472 137896 283524 137902
rect 283472 137838 283524 137844
rect 283668 135182 283696 286350
rect 285864 286068 285916 286074
rect 285864 286010 285916 286016
rect 284300 284980 284352 284986
rect 284300 284922 284352 284928
rect 283748 284096 283800 284102
rect 283748 284038 283800 284044
rect 283656 135176 283708 135182
rect 283656 135118 283708 135124
rect 283380 108656 283432 108662
rect 283380 108598 283432 108604
rect 283760 104854 283788 284038
rect 284312 157962 284340 284922
rect 285772 273284 285824 273290
rect 285772 273226 285824 273232
rect 284392 266484 284444 266490
rect 284392 266426 284444 266432
rect 284300 157956 284352 157962
rect 284300 157898 284352 157904
rect 284404 144498 284432 266426
rect 284484 249824 284536 249830
rect 284484 249766 284536 249772
rect 284392 144492 284444 144498
rect 284392 144434 284444 144440
rect 284496 131102 284524 249766
rect 284576 188352 284628 188358
rect 284576 188294 284628 188300
rect 284484 131096 284536 131102
rect 284484 131038 284536 131044
rect 284588 128246 284616 188294
rect 285680 187060 285732 187066
rect 285680 187002 285732 187008
rect 284668 186992 284720 186998
rect 284668 186934 284720 186940
rect 284680 129606 284708 186934
rect 284944 184204 284996 184210
rect 284944 184146 284996 184152
rect 284852 181688 284904 181694
rect 284852 181630 284904 181636
rect 284760 180192 284812 180198
rect 284760 180134 284812 180140
rect 284668 129600 284720 129606
rect 284668 129542 284720 129548
rect 284576 128240 284628 128246
rect 284576 128182 284628 128188
rect 284772 127702 284800 180134
rect 284864 129674 284892 181630
rect 284956 148918 284984 184146
rect 285128 181484 285180 181490
rect 285128 181426 285180 181432
rect 285036 180328 285088 180334
rect 285036 180270 285088 180276
rect 285048 151774 285076 180270
rect 285036 151768 285088 151774
rect 285036 151710 285088 151716
rect 284944 148912 284996 148918
rect 284944 148854 284996 148860
rect 285140 131034 285168 181426
rect 285692 156602 285720 187002
rect 285680 156596 285732 156602
rect 285680 156538 285732 156544
rect 285784 132394 285812 273226
rect 285876 161226 285904 286010
rect 286336 256698 286364 484366
rect 287060 288448 287112 288454
rect 287060 288390 287112 288396
rect 286508 259480 286560 259486
rect 286508 259422 286560 259428
rect 286324 256692 286376 256698
rect 286324 256634 286376 256640
rect 286324 198008 286376 198014
rect 286324 197950 286376 197956
rect 286232 184408 286284 184414
rect 286232 184350 286284 184356
rect 285956 184272 286008 184278
rect 285956 184214 286008 184220
rect 285864 161220 285916 161226
rect 285864 161162 285916 161168
rect 285772 132388 285824 132394
rect 285772 132330 285824 132336
rect 285128 131028 285180 131034
rect 285128 130970 285180 130976
rect 284852 129668 284904 129674
rect 284852 129610 284904 129616
rect 284760 127696 284812 127702
rect 284760 127638 284812 127644
rect 283748 104848 283800 104854
rect 283748 104790 283800 104796
rect 281540 104576 281592 104582
rect 281540 104518 281592 104524
rect 283288 104576 283340 104582
rect 283288 104518 283340 104524
rect 281552 104009 281580 104518
rect 281538 104000 281594 104009
rect 281538 103935 281594 103944
rect 282828 103488 282880 103494
rect 282828 103430 282880 103436
rect 282000 103284 282052 103290
rect 282000 103226 282052 103232
rect 282012 102513 282040 103226
rect 282840 103193 282868 103430
rect 282826 103184 282882 103193
rect 282826 103119 282882 103128
rect 281998 102504 282054 102513
rect 281998 102439 282054 102448
rect 281630 101688 281686 101697
rect 281630 101623 281686 101632
rect 281538 99376 281594 99385
rect 281538 99311 281594 99320
rect 279422 98152 279478 98161
rect 279422 98087 279478 98096
rect 267556 97368 267608 97374
rect 267556 97310 267608 97316
rect 267280 97300 267332 97306
rect 267280 97242 267332 97248
rect 267096 96144 267148 96150
rect 267096 96086 267148 96092
rect 267292 95198 267320 97242
rect 267280 95192 267332 95198
rect 267280 95134 267332 95140
rect 267568 93838 267596 97310
rect 279330 96656 279386 96665
rect 279330 96591 279386 96600
rect 279344 96354 279372 96591
rect 279436 96422 279464 98087
rect 279514 97336 279570 97345
rect 279514 97271 279570 97280
rect 279424 96416 279476 96422
rect 279424 96358 279476 96364
rect 279332 96348 279384 96354
rect 279332 96290 279384 96296
rect 279240 96280 279292 96286
rect 279240 96222 279292 96228
rect 279252 96121 279280 96222
rect 279528 96150 279556 97271
rect 279516 96144 279568 96150
rect 279238 96112 279294 96121
rect 279516 96086 279568 96092
rect 279238 96047 279294 96056
rect 270972 95198 271000 96016
rect 270960 95192 271012 95198
rect 270960 95134 271012 95140
rect 276952 93838 276980 96016
rect 281552 95130 281580 99311
rect 281540 95124 281592 95130
rect 281540 95066 281592 95072
rect 281644 95062 281672 101623
rect 285968 100298 285996 184214
rect 286048 180260 286100 180266
rect 286048 180202 286100 180208
rect 286060 114374 286088 180202
rect 286140 177540 286192 177546
rect 286140 177482 286192 177488
rect 286152 118590 286180 177482
rect 286244 133890 286272 184350
rect 286336 153338 286364 197950
rect 286416 191140 286468 191146
rect 286416 191082 286468 191088
rect 286428 154154 286456 191082
rect 286416 154148 286468 154154
rect 286416 154090 286468 154096
rect 286324 153332 286376 153338
rect 286324 153274 286376 153280
rect 286232 133884 286284 133890
rect 286232 133826 286284 133832
rect 286140 118584 286192 118590
rect 286140 118526 286192 118532
rect 286048 114368 286100 114374
rect 286048 114310 286100 114316
rect 286520 112742 286548 259422
rect 286508 112736 286560 112742
rect 286508 112678 286560 112684
rect 287072 110090 287100 288390
rect 287336 287972 287388 287978
rect 287336 287914 287388 287920
rect 287152 287292 287204 287298
rect 287152 287234 287204 287240
rect 287060 110084 287112 110090
rect 287060 110026 287112 110032
rect 287164 109954 287192 287234
rect 287244 287224 287296 287230
rect 287244 287166 287296 287172
rect 287256 111110 287284 287166
rect 287348 114850 287376 287914
rect 289820 287904 289872 287910
rect 289820 287846 289872 287852
rect 288716 284640 288768 284646
rect 288716 284582 288768 284588
rect 287428 280288 287480 280294
rect 287428 280230 287480 280236
rect 287440 139874 287468 280230
rect 288532 271992 288584 271998
rect 288532 271934 288584 271940
rect 287520 238060 287572 238066
rect 287520 238002 287572 238008
rect 287532 159186 287560 238002
rect 287610 180296 287666 180305
rect 287610 180231 287666 180240
rect 287520 159180 287572 159186
rect 287520 159122 287572 159128
rect 287428 139868 287480 139874
rect 287428 139810 287480 139816
rect 287336 114844 287388 114850
rect 287336 114786 287388 114792
rect 287624 113490 287652 180231
rect 287888 177744 287940 177750
rect 287888 177686 287940 177692
rect 287796 177608 287848 177614
rect 287796 177550 287848 177556
rect 287704 177336 287756 177342
rect 287704 177278 287756 177284
rect 287612 113484 287664 113490
rect 287612 113426 287664 113432
rect 287716 111178 287744 177278
rect 287808 116482 287836 177550
rect 287900 124506 287928 177686
rect 288440 175976 288492 175982
rect 288440 175918 288492 175924
rect 288452 149258 288480 175918
rect 288440 149252 288492 149258
rect 288440 149194 288492 149200
rect 287888 124500 287940 124506
rect 287888 124442 287940 124448
rect 288544 123554 288572 271934
rect 288624 269136 288676 269142
rect 288624 269078 288676 269084
rect 288636 126750 288664 269078
rect 288728 145110 288756 284582
rect 289268 284504 289320 284510
rect 289268 284446 289320 284452
rect 288808 258188 288860 258194
rect 288808 258130 288860 258136
rect 288820 157894 288848 258130
rect 289176 182844 289228 182850
rect 289176 182786 289228 182792
rect 288898 180568 288954 180577
rect 288898 180503 288954 180512
rect 288808 157888 288860 157894
rect 288808 157830 288860 157836
rect 288716 145104 288768 145110
rect 288716 145046 288768 145052
rect 288624 126744 288676 126750
rect 288624 126686 288676 126692
rect 288532 123548 288584 123554
rect 288532 123490 288584 123496
rect 287796 116476 287848 116482
rect 287796 116418 287848 116424
rect 287704 111172 287756 111178
rect 287704 111114 287756 111120
rect 287244 111104 287296 111110
rect 287244 111046 287296 111052
rect 287152 109948 287204 109954
rect 287152 109890 287204 109896
rect 288912 105126 288940 180503
rect 289082 180024 289138 180033
rect 289082 179959 289138 179968
rect 288992 177676 289044 177682
rect 288992 177618 289044 177624
rect 289004 109002 289032 177618
rect 289096 117298 289124 179959
rect 289188 139398 289216 182786
rect 289176 139392 289228 139398
rect 289176 139334 289228 139340
rect 289084 117292 289136 117298
rect 289084 117234 289136 117240
rect 288992 108996 289044 109002
rect 288992 108938 289044 108944
rect 288900 105120 288952 105126
rect 288900 105062 288952 105068
rect 289280 103290 289308 284446
rect 289832 107642 289860 287846
rect 291200 287428 291252 287434
rect 291200 287370 291252 287376
rect 289912 280220 289964 280226
rect 289912 280162 289964 280168
rect 289924 143546 289952 280162
rect 290096 238264 290148 238270
rect 290096 238206 290148 238212
rect 290004 238196 290056 238202
rect 290004 238138 290056 238144
rect 289912 143540 289964 143546
rect 289912 143482 289964 143488
rect 289820 107636 289872 107642
rect 289820 107578 289872 107584
rect 290016 103494 290044 238138
rect 290108 118658 290136 238206
rect 290188 238128 290240 238134
rect 290188 238070 290240 238076
rect 290200 137970 290228 238070
rect 290280 182912 290332 182918
rect 290280 182854 290332 182860
rect 290188 137964 290240 137970
rect 290188 137906 290240 137912
rect 290292 136610 290320 182854
rect 290280 136604 290332 136610
rect 290280 136546 290332 136552
rect 291212 132462 291240 287370
rect 292580 287360 292632 287366
rect 292580 287302 292632 287308
rect 291292 267844 291344 267850
rect 291292 267786 291344 267792
rect 291304 155922 291332 267786
rect 291936 267776 291988 267782
rect 291936 267718 291988 267724
rect 291844 251252 291896 251258
rect 291844 251194 291896 251200
rect 291856 167006 291884 251194
rect 291948 233238 291976 267718
rect 291936 233232 291988 233238
rect 291936 233174 291988 233180
rect 291844 167000 291896 167006
rect 291844 166942 291896 166948
rect 292592 157350 292620 287302
rect 292672 258120 292724 258126
rect 292672 258062 292724 258068
rect 292580 157344 292632 157350
rect 292580 157286 292632 157292
rect 291292 155916 291344 155922
rect 291292 155858 291344 155864
rect 292684 149054 292712 258062
rect 292764 242956 292816 242962
rect 292764 242898 292816 242904
rect 292776 153202 292804 242898
rect 294616 241466 294644 524418
rect 295996 244254 296024 683130
rect 305644 378208 305696 378214
rect 305644 378150 305696 378156
rect 298744 284368 298796 284374
rect 298744 284310 298796 284316
rect 295984 244248 296036 244254
rect 295984 244190 296036 244196
rect 294604 241460 294656 241466
rect 294604 241402 294656 241408
rect 292764 153196 292816 153202
rect 292764 153138 292816 153144
rect 292672 149048 292724 149054
rect 292672 148990 292724 148996
rect 298756 139398 298784 284310
rect 305656 282878 305684 378150
rect 316684 311908 316736 311914
rect 316684 311850 316736 311856
rect 305644 282872 305696 282878
rect 305644 282814 305696 282820
rect 316696 266354 316724 311850
rect 347056 296002 347084 699654
rect 347044 295996 347096 296002
rect 347044 295938 347096 295944
rect 316684 266348 316736 266354
rect 316684 266290 316736 266296
rect 364352 239698 364380 702406
rect 397472 700466 397500 703520
rect 413664 700534 413692 703520
rect 413652 700528 413704 700534
rect 413652 700470 413704 700476
rect 397460 700460 397512 700466
rect 397460 700402 397512 700408
rect 429856 699718 429884 703520
rect 422944 699712 422996 699718
rect 422944 699654 422996 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 422956 289134 422984 699654
rect 422944 289128 422996 289134
rect 422944 289070 422996 289076
rect 454684 278792 454736 278798
rect 454684 278734 454736 278740
rect 364340 239692 364392 239698
rect 364340 239634 364392 239640
rect 298744 139392 298796 139398
rect 298744 139334 298796 139340
rect 291200 132456 291252 132462
rect 291200 132398 291252 132404
rect 454696 126954 454724 278734
rect 462332 240922 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 462320 240916 462372 240922
rect 462320 240858 462372 240864
rect 494072 239630 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 699718 527220 703520
rect 529204 700392 529256 700398
rect 529204 700334 529256 700340
rect 526444 699712 526496 699718
rect 526444 699654 526496 699660
rect 527180 699712 527232 699718
rect 527180 699654 527232 699660
rect 526456 276010 526484 699654
rect 526444 276004 526496 276010
rect 526444 275946 526496 275952
rect 529216 240106 529244 700334
rect 543476 700330 543504 703520
rect 559668 700398 559696 703520
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580262 591016 580318 591025
rect 580262 590951 580318 590960
rect 579894 564360 579950 564369
rect 579894 564295 579950 564304
rect 579908 563106 579936 564295
rect 579896 563100 579948 563106
rect 579896 563042 579948 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580184 470626 580212 471407
rect 580172 470620 580224 470626
rect 580172 470562 580224 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 579986 404968 580042 404977
rect 579986 404903 580042 404912
rect 580000 404394 580028 404903
rect 579988 404388 580040 404394
rect 579988 404330 580040 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 579618 325272 579674 325281
rect 579618 325207 579674 325216
rect 579632 324358 579660 325207
rect 579620 324352 579672 324358
rect 579620 324294 579672 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 565084 266416 565136 266422
rect 565084 266358 565136 266364
rect 529204 240100 529256 240106
rect 529204 240042 529256 240048
rect 494060 239624 494112 239630
rect 494060 239566 494112 239572
rect 454684 126948 454736 126954
rect 454684 126890 454736 126896
rect 290096 118652 290148 118658
rect 290096 118594 290148 118600
rect 290004 103488 290056 103494
rect 290004 103430 290056 103436
rect 289268 103284 289320 103290
rect 289268 103226 289320 103232
rect 565096 100706 565124 266358
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 579802 245576 579858 245585
rect 579802 245511 579858 245520
rect 579816 244322 579844 245511
rect 579804 244316 579856 244322
rect 579804 244258 579856 244264
rect 580276 240854 580304 590951
rect 580354 577688 580410 577697
rect 580354 577623 580410 577632
rect 580368 242214 580396 577623
rect 580446 365120 580502 365129
rect 580446 365055 580502 365064
rect 580356 242208 580408 242214
rect 580356 242150 580408 242156
rect 580264 240848 580316 240854
rect 580264 240790 580316 240796
rect 580460 240786 580488 365055
rect 580448 240780 580500 240786
rect 580448 240722 580500 240728
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580264 199436 580316 199442
rect 580264 199378 580316 199384
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 579988 179376 580040 179382
rect 579988 179318 580040 179324
rect 580000 179217 580028 179318
rect 579986 179208 580042 179217
rect 579986 179143 580042 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 565084 100700 565136 100706
rect 565084 100642 565136 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 282276 100292 282328 100298
rect 282276 100234 282328 100240
rect 285956 100292 286008 100298
rect 285956 100234 286008 100240
rect 282288 100201 282316 100234
rect 282274 100192 282330 100201
rect 282274 100127 282330 100136
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 281632 95056 281684 95062
rect 281632 94998 281684 95004
rect 267556 93832 267608 93838
rect 267556 93774 267608 93780
rect 276940 93832 276992 93838
rect 276940 93774 276992 93780
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580276 46345 580304 199378
rect 580262 46336 580318 46345
rect 580262 46271 580318 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 267004 6860 267056 6866
rect 267004 6802 267056 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 265808 4820 265860 4826
rect 265808 4762 265860 4768
rect 235816 3528 235868 3534
rect 235816 3470 235868 3476
rect 233884 3460 233936 3466
rect 233884 3402 233936 3408
rect 235828 480 235856 3470
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3330 553832 3386 553888
rect 2962 527856 3018 527912
rect 3330 501744 3386 501800
rect 3054 475632 3110 475688
rect 3330 462576 3386 462632
rect 3330 449520 3386 449576
rect 3146 423544 3202 423600
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3054 306176 3110 306232
rect 3330 293120 3386 293176
rect 3514 514800 3570 514856
rect 3330 267144 3386 267200
rect 3422 254088 3478 254144
rect 3054 241032 3110 241088
rect 3606 410488 3662 410544
rect 3330 214920 3386 214976
rect 3054 201864 3110 201920
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3698 149776 3754 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 3422 97588 3424 97608
rect 3424 97588 3476 97608
rect 3476 97588 3478 97608
rect 3422 97552 3478 97588
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 97814 176704 97870 176760
rect 103334 176704 103390 176760
rect 107014 176704 107070 176760
rect 108118 176704 108174 176760
rect 110050 176704 110106 176760
rect 110694 176704 110750 176760
rect 112626 176704 112682 176760
rect 114006 176704 114062 176760
rect 114374 176704 114430 176760
rect 115846 176724 115902 176760
rect 115846 176704 115848 176724
rect 115848 176704 115900 176724
rect 115900 176704 115902 176724
rect 116950 176740 116952 176760
rect 116952 176740 117004 176760
rect 117004 176740 117006 176760
rect 116950 176704 117006 176740
rect 118422 176704 118478 176760
rect 120814 176704 120870 176760
rect 122286 176704 122342 176760
rect 124494 176704 124550 176760
rect 127990 176704 128046 176760
rect 129462 176704 129518 176760
rect 98366 175344 98422 175400
rect 99470 175344 99526 175400
rect 100758 175344 100814 175400
rect 102046 175344 102102 175400
rect 104622 175344 104678 175400
rect 105726 175344 105782 175400
rect 130934 176704 130990 176760
rect 133142 176704 133198 176760
rect 134522 176704 134578 176760
rect 148230 176704 148286 176760
rect 135718 175480 135774 175536
rect 128174 175344 128230 175400
rect 132038 175344 132094 175400
rect 158902 175344 158958 175400
rect 119434 174936 119490 174992
rect 123114 174936 123170 174992
rect 125690 174936 125746 174992
rect 66166 129240 66222 129296
rect 66074 128016 66130 128072
rect 65982 126248 66038 126304
rect 65890 123528 65946 123584
rect 65798 122576 65854 122632
rect 65982 102312 66038 102368
rect 67638 125160 67694 125216
rect 66166 100680 66222 100736
rect 67822 120808 67878 120864
rect 67822 94832 67878 94888
rect 67638 94696 67694 94752
rect 66166 94560 66222 94616
rect 65982 94424 66038 94480
rect 102966 93608 103022 93664
rect 104254 93608 104310 93664
rect 105542 93608 105598 93664
rect 106462 93608 106518 93664
rect 107750 93628 107806 93664
rect 107750 93608 107752 93628
rect 107752 93608 107804 93628
rect 107804 93608 107806 93628
rect 90270 93472 90326 93528
rect 101862 93472 101918 93528
rect 109222 93644 109224 93664
rect 109224 93644 109276 93664
rect 109276 93644 109278 93664
rect 109222 93608 109278 93644
rect 110142 93200 110198 93256
rect 84382 92404 84438 92440
rect 84382 92384 84384 92404
rect 84384 92384 84436 92404
rect 84436 92384 84438 92404
rect 86682 92384 86738 92440
rect 88062 92384 88118 92440
rect 89074 92384 89130 92440
rect 91466 92384 91522 92440
rect 94962 92384 95018 92440
rect 100022 92384 100078 92440
rect 105726 92384 105782 92440
rect 108118 92384 108174 92440
rect 109958 92384 110014 92440
rect 75734 91704 75790 91760
rect 86774 91160 86830 91216
rect 93214 91568 93270 91624
rect 95054 91704 95110 91760
rect 97814 91704 97870 91760
rect 100574 91704 100630 91760
rect 96342 91568 96398 91624
rect 97538 91568 97594 91624
rect 99286 91568 99342 91624
rect 99102 91160 99158 91216
rect 104622 91160 104678 91216
rect 124126 94152 124182 94208
rect 117134 94036 117190 94072
rect 117134 94016 117136 94036
rect 117136 94016 117188 94036
rect 117188 94016 117190 94036
rect 122102 94016 122158 94072
rect 118238 93900 118294 93936
rect 118238 93880 118240 93900
rect 118240 93880 118292 93900
rect 118292 93880 118294 93900
rect 119710 93608 119766 93664
rect 111798 93472 111854 93528
rect 125414 93472 125470 93528
rect 128174 93200 128230 93256
rect 126058 93064 126114 93120
rect 113178 92520 113234 92576
rect 110970 92384 111026 92440
rect 111982 92384 112038 92440
rect 112350 92384 112406 92440
rect 113362 92384 113418 92440
rect 114374 92384 114430 92440
rect 115202 92384 115258 92440
rect 115846 92384 115902 92440
rect 118054 92420 118056 92440
rect 118056 92420 118108 92440
rect 118108 92420 118110 92440
rect 118054 92384 118110 92420
rect 120262 92384 120318 92440
rect 121182 92384 121238 92440
rect 125782 92384 125838 92440
rect 115478 91432 115534 91488
rect 121918 91840 121974 91896
rect 126610 91840 126666 91896
rect 122838 91432 122894 91488
rect 125322 91432 125378 91488
rect 123574 91160 123630 91216
rect 126702 91160 126758 91216
rect 151634 94288 151690 94344
rect 151542 93880 151598 93936
rect 135718 93336 135774 93392
rect 151726 94016 151782 94072
rect 129462 92384 129518 92440
rect 132406 92384 132462 92440
rect 134430 92384 134486 92440
rect 153106 92404 153162 92440
rect 153106 92384 153108 92404
rect 153108 92384 153160 92404
rect 153160 92384 153162 92404
rect 130750 91160 130806 91216
rect 165526 94424 165582 94480
rect 133326 91160 133382 91216
rect 169022 171536 169078 171592
rect 167550 110064 167606 110120
rect 167550 108704 167606 108760
rect 167826 92248 167882 92304
rect 168286 111732 168288 111752
rect 168288 111732 168340 111752
rect 168340 111732 168342 111752
rect 168286 111696 168342 111732
rect 169022 93744 169078 93800
rect 169206 91976 169262 92032
rect 171782 92112 171838 92168
rect 180154 91296 180210 91352
rect 192850 179968 192906 180024
rect 194230 180104 194286 180160
rect 195150 177520 195206 177576
rect 196806 257352 196862 257408
rect 198278 282920 198334 282976
rect 197358 281580 197414 281616
rect 197358 281560 197360 281580
rect 197360 281560 197412 281580
rect 197412 281560 197414 281580
rect 197358 280220 197414 280256
rect 197358 280200 197360 280220
rect 197360 280200 197412 280220
rect 197412 280200 197414 280220
rect 197358 279384 197414 279440
rect 197450 277208 197506 277264
rect 197358 275848 197414 275904
rect 198186 274488 198242 274544
rect 197450 272856 197506 272912
rect 197358 272312 197414 272368
rect 197358 269320 197414 269376
rect 197450 268776 197506 268832
rect 197358 267960 197414 268016
rect 197450 267144 197506 267200
rect 197358 266600 197414 266656
rect 197450 265784 197506 265840
rect 197358 265240 197414 265296
rect 197358 264424 197414 264480
rect 197358 263628 197414 263664
rect 197358 263608 197360 263628
rect 197360 263608 197412 263628
rect 197412 263608 197414 263628
rect 197358 261432 197414 261488
rect 197450 259256 197506 259312
rect 197358 258712 197414 258768
rect 197358 257896 197414 257952
rect 198094 256536 198150 256592
rect 197450 255176 197506 255232
rect 197358 254360 197414 254416
rect 197726 253544 197782 253600
rect 197358 253000 197414 253056
rect 197358 250008 197414 250064
rect 197634 249464 197690 249520
rect 197542 248648 197598 248704
rect 197266 247288 197322 247344
rect 197358 245928 197414 245984
rect 197358 243752 197414 243808
rect 197450 242936 197506 242992
rect 197174 241576 197230 241632
rect 197910 251640 197966 251696
rect 198002 247832 198058 247888
rect 198002 242120 198058 242176
rect 197910 233824 197966 233880
rect 200762 285776 200818 285832
rect 206650 284688 206706 284744
rect 215850 285640 215906 285696
rect 219714 284416 219770 284472
rect 221554 286048 221610 286104
rect 221186 285912 221242 285968
rect 226890 286184 226946 286240
rect 233698 284552 233754 284608
rect 239034 284280 239090 284336
rect 240782 284824 240838 284880
rect 243358 284008 243414 284064
rect 198646 283736 198702 283792
rect 199566 282376 199622 282432
rect 198554 280744 198610 280800
rect 199474 278568 199530 278624
rect 198646 278024 198702 278080
rect 198554 270952 198610 271008
rect 198462 263064 198518 263120
rect 198370 255720 198426 255776
rect 198370 252184 198426 252240
rect 198278 232600 198334 232656
rect 198094 232464 198150 232520
rect 198554 186904 198610 186960
rect 198462 182824 198518 182880
rect 199290 262248 199346 262304
rect 199198 245112 199254 245168
rect 198646 181328 198702 181384
rect 199382 260072 199438 260128
rect 199658 276664 199714 276720
rect 199750 275032 199806 275088
rect 200026 273672 200082 273728
rect 199934 271496 199990 271552
rect 199842 270136 199898 270192
rect 199750 182960 199806 183016
rect 244278 278840 244334 278896
rect 244370 278024 244426 278080
rect 244370 271496 244426 271552
rect 244094 250552 244150 250608
rect 244002 244296 244058 244352
rect 243910 240488 243966 240544
rect 200118 240080 200174 240136
rect 200118 180240 200174 180296
rect 198370 177248 198426 177304
rect 207938 237904 207994 237960
rect 210698 180376 210754 180432
rect 225786 180512 225842 180568
rect 213918 176160 213974 176216
rect 227718 176160 227774 176216
rect 213918 175072 213974 175128
rect 214010 174664 214066 174720
rect 213918 173712 213974 173768
rect 214010 173304 214066 173360
rect 213918 172388 213920 172408
rect 213920 172388 213972 172408
rect 213972 172388 213974 172408
rect 213918 172352 213974 172388
rect 214010 171944 214066 172000
rect 213918 170720 213974 170776
rect 213918 169652 213974 169688
rect 213918 169632 213920 169652
rect 213920 169632 213972 169652
rect 213972 169632 213974 169652
rect 214010 169360 214066 169416
rect 213918 168000 213974 168056
rect 214010 167864 214066 167920
rect 213918 166948 213920 166968
rect 213920 166948 213972 166968
rect 213972 166948 213974 166968
rect 213918 166912 213974 166948
rect 214010 166640 214066 166696
rect 214102 166096 214158 166152
rect 213918 165452 213920 165472
rect 213920 165452 213972 165472
rect 213972 165452 213974 165472
rect 213918 165416 213974 165452
rect 214010 164736 214066 164792
rect 213918 163920 213974 163976
rect 214010 163376 214066 163432
rect 213918 162560 213974 162616
rect 214010 162016 214066 162072
rect 214654 170992 214710 171048
rect 213918 161372 213920 161392
rect 213920 161372 213972 161392
rect 213972 161372 213974 161392
rect 213918 161336 213974 161372
rect 213918 159840 213974 159896
rect 214010 159432 214066 159488
rect 214746 160792 214802 160848
rect 214470 158616 214526 158672
rect 213918 158072 213974 158128
rect 213918 157276 213974 157312
rect 213918 157256 213920 157276
rect 213920 157256 213972 157276
rect 213972 157256 213974 157276
rect 214010 156848 214066 156904
rect 213918 155916 213974 155952
rect 213918 155896 213920 155916
rect 213920 155896 213972 155916
rect 213972 155896 213974 155916
rect 214010 155352 214066 155408
rect 214010 153856 214066 153912
rect 213918 153448 213974 153504
rect 213918 152632 213974 152688
rect 214746 152088 214802 152144
rect 214838 151952 214894 152008
rect 214010 150864 214066 150920
rect 213182 150184 213238 150240
rect 213918 149504 213974 149560
rect 213918 148688 213974 148744
rect 213918 148008 213974 148064
rect 214010 146648 214066 146704
rect 213918 146396 213974 146432
rect 213918 146376 213920 146396
rect 213920 146376 213972 146396
rect 213972 146376 213974 146396
rect 214010 145288 214066 145344
rect 213918 144916 213920 144936
rect 213920 144916 213972 144936
rect 213972 144916 213974 144936
rect 213918 144880 213974 144916
rect 214470 143928 214526 143984
rect 213918 143556 213920 143576
rect 213920 143556 213972 143576
rect 213972 143556 213974 143576
rect 213918 143520 213974 143556
rect 214010 142704 214066 142760
rect 213918 142296 213974 142352
rect 214010 141344 214066 141400
rect 213918 140936 213974 140992
rect 214010 139984 214066 140040
rect 213918 139576 213974 139632
rect 213918 136720 213974 136776
rect 214010 136040 214066 136096
rect 214102 135632 214158 135688
rect 213918 135380 213974 135416
rect 213918 135360 213920 135380
rect 213920 135360 213972 135380
rect 213972 135360 213974 135380
rect 213918 134272 213974 134328
rect 214746 150728 214802 150784
rect 229190 169496 229246 169552
rect 229374 174256 229430 174312
rect 229282 154264 229338 154320
rect 229558 168952 229614 169008
rect 229466 161472 229522 161528
rect 229374 153312 229430 153368
rect 229098 150592 229154 150648
rect 214838 138080 214894 138136
rect 214010 132776 214066 132832
rect 213918 132540 213920 132560
rect 213920 132540 213972 132560
rect 213972 132540 213974 132560
rect 213918 132504 213974 132540
rect 214010 131416 214066 131472
rect 213918 131164 213974 131200
rect 213918 131144 213920 131164
rect 213920 131144 213972 131164
rect 213972 131144 213974 131164
rect 214010 130056 214066 130112
rect 213918 129820 213920 129840
rect 213920 129820 213972 129840
rect 213972 129820 213974 129840
rect 213918 129784 213974 129820
rect 214010 128832 214066 128888
rect 213918 128444 213974 128480
rect 213918 128424 213920 128444
rect 213920 128424 213972 128444
rect 213972 128424 213974 128444
rect 214010 127472 214066 127528
rect 213918 127084 213974 127120
rect 213918 127064 213920 127084
rect 213920 127064 213972 127084
rect 213972 127064 213974 127084
rect 214010 126112 214066 126168
rect 213918 125724 213974 125760
rect 213918 125704 213920 125724
rect 213920 125704 213972 125724
rect 213972 125704 213974 125724
rect 214010 124752 214066 124808
rect 213918 124228 213974 124264
rect 213918 124208 213920 124228
rect 213920 124208 213972 124228
rect 213972 124208 213974 124228
rect 214010 123528 214066 123584
rect 213918 123120 213974 123176
rect 214010 122168 214066 122224
rect 213918 121760 213974 121816
rect 214010 120808 214066 120864
rect 213918 120400 213974 120456
rect 213918 119584 213974 119640
rect 214010 118904 214066 118960
rect 213182 118768 213238 118824
rect 213918 117308 213920 117328
rect 213920 117308 213972 117328
rect 213972 117308 213974 117328
rect 213918 117272 213974 117308
rect 214010 116184 214066 116240
rect 213918 115912 213974 115968
rect 214010 114960 214066 115016
rect 213918 114572 213974 114608
rect 213918 114552 213920 114572
rect 213920 114552 213972 114572
rect 213972 114552 213974 114572
rect 214010 113600 214066 113656
rect 213918 113212 213974 113248
rect 213918 113192 213920 113212
rect 213920 113192 213972 113212
rect 213972 113192 213974 113212
rect 214010 112240 214066 112296
rect 213918 111868 213920 111888
rect 213920 111868 213972 111888
rect 213972 111868 213974 111888
rect 213918 111832 213974 111868
rect 213918 110492 213974 110528
rect 213918 110472 213920 110492
rect 213920 110472 213972 110492
rect 213972 110472 213974 110492
rect 214010 109656 214066 109712
rect 213918 109132 213974 109168
rect 213918 109112 213920 109132
rect 213920 109112 213972 109132
rect 213972 109112 213974 109132
rect 213918 108296 213974 108352
rect 214010 106936 214066 106992
rect 213918 106528 213974 106584
rect 214102 105712 214158 105768
rect 214010 105304 214066 105360
rect 213918 105052 213974 105088
rect 213918 105032 213920 105052
rect 213920 105032 213972 105052
rect 213972 105032 213974 105052
rect 213918 103672 213974 103728
rect 214010 102584 214066 102640
rect 213918 102312 213974 102368
rect 214194 99728 214250 99784
rect 214102 99456 214158 99512
rect 213918 98368 213974 98424
rect 214010 97960 214066 98016
rect 213918 97008 213974 97064
rect 213918 95784 213974 95840
rect 214378 100816 214434 100872
rect 230478 158616 230534 158672
rect 230754 174664 230810 174720
rect 230662 173712 230718 173768
rect 230662 159568 230718 159624
rect 230478 155796 230480 155816
rect 230480 155796 230532 155816
rect 230532 155796 230534 155816
rect 230478 155760 230534 155796
rect 230478 155252 230480 155272
rect 230480 155252 230532 155272
rect 230532 155252 230534 155272
rect 230478 155216 230534 155252
rect 230570 154808 230626 154864
rect 230846 153856 230902 153912
rect 230754 151000 230810 151056
rect 230754 149640 230810 149696
rect 230570 146784 230626 146840
rect 230846 145832 230902 145888
rect 231122 173304 231178 173360
rect 231398 177656 231454 177712
rect 231214 170484 231216 170504
rect 231216 170484 231268 170504
rect 231268 170484 231270 170504
rect 231030 161880 231086 161936
rect 231030 157664 231086 157720
rect 231214 170448 231270 170484
rect 231490 172760 231546 172816
rect 231490 171808 231546 171864
rect 231306 169904 231362 169960
rect 231490 167592 231546 167648
rect 231398 167048 231454 167104
rect 231306 166676 231308 166696
rect 231308 166676 231360 166696
rect 231360 166676 231362 166696
rect 231306 166640 231362 166676
rect 231398 164772 231400 164792
rect 231400 164772 231452 164792
rect 231452 164772 231454 164792
rect 231398 164736 231454 164772
rect 231398 163820 231400 163840
rect 231400 163820 231452 163840
rect 231452 163820 231454 163840
rect 231398 163784 231454 163820
rect 231490 162832 231546 162888
rect 231214 159024 231270 159080
rect 231490 156712 231546 156768
rect 231122 156168 231178 156224
rect 231122 152496 231178 152552
rect 231306 151952 231362 152008
rect 231766 175208 231822 175264
rect 231766 172352 231822 172408
rect 231674 171400 231730 171456
rect 231582 151544 231638 151600
rect 231214 148724 231216 148744
rect 231216 148724 231268 148744
rect 231268 148724 231270 148744
rect 231214 148688 231270 148724
rect 231766 170856 231822 170912
rect 231766 168544 231822 168600
rect 231766 168000 231822 168056
rect 231766 166096 231822 166152
rect 231766 165724 231768 165744
rect 231768 165724 231820 165744
rect 231820 165724 231822 165744
rect 231766 165688 231822 165724
rect 231766 165144 231822 165200
rect 231766 164328 231822 164384
rect 231766 163412 231768 163432
rect 231768 163412 231820 163432
rect 231820 163412 231822 163432
rect 231766 163376 231822 163412
rect 231766 160928 231822 160984
rect 231766 160556 231768 160576
rect 231768 160556 231820 160576
rect 231820 160556 231822 160576
rect 231766 160520 231822 160556
rect 231766 159976 231822 160032
rect 231766 158072 231822 158128
rect 231766 157120 231822 157176
rect 231766 152904 231822 152960
rect 231766 150048 231822 150104
rect 231766 148144 231822 148200
rect 231766 147192 231822 147248
rect 231674 146240 231730 146296
rect 231306 145288 231362 145344
rect 231122 144880 231178 144936
rect 231306 144336 231362 144392
rect 231306 142976 231362 143032
rect 231766 143928 231822 143984
rect 231766 143420 231768 143440
rect 231768 143420 231820 143440
rect 231820 143420 231822 143440
rect 231766 143384 231822 143420
rect 231674 142432 231730 142488
rect 231766 142060 231768 142080
rect 231768 142060 231820 142080
rect 231820 142060 231822 142080
rect 231766 142024 231822 142060
rect 231766 141652 231768 141672
rect 231768 141652 231820 141672
rect 231820 141652 231822 141672
rect 231766 141616 231822 141652
rect 231398 141072 231454 141128
rect 231214 140120 231270 140176
rect 230938 138216 230994 138272
rect 229650 136856 229706 136912
rect 215114 134136 215170 134192
rect 214838 117544 214894 117600
rect 215022 110880 215078 110936
rect 214930 107616 214986 107672
rect 214746 93064 214802 93120
rect 230662 133456 230718 133512
rect 231030 130600 231086 130656
rect 230938 129784 230994 129840
rect 231122 124480 231178 124536
rect 230846 124072 230902 124128
rect 230754 123120 230810 123176
rect 230570 118904 230626 118960
rect 230570 118396 230572 118416
rect 230572 118396 230624 118416
rect 230624 118396 230626 118416
rect 230570 118360 230626 118396
rect 231122 122168 231178 122224
rect 230754 117408 230810 117464
rect 230938 115096 230994 115152
rect 231030 114144 231086 114200
rect 230938 109792 230994 109848
rect 231030 107888 231086 107944
rect 230754 105576 230810 105632
rect 230754 104660 230756 104680
rect 230756 104660 230808 104680
rect 230808 104660 230810 104680
rect 230754 104624 230810 104660
rect 230938 104216 230994 104272
rect 230570 102720 230626 102776
rect 230662 101768 230718 101824
rect 231766 139712 231822 139768
rect 231766 139168 231822 139224
rect 231950 147736 232006 147792
rect 231306 138796 231308 138816
rect 231308 138796 231360 138816
rect 231360 138796 231362 138816
rect 231306 138760 231362 138796
rect 231766 137844 231768 137864
rect 231768 137844 231820 137864
rect 231820 137844 231822 137864
rect 231766 137808 231822 137844
rect 231674 137264 231730 137320
rect 231398 135904 231454 135960
rect 231766 135360 231822 135416
rect 231766 134952 231822 135008
rect 231674 134408 231730 134464
rect 231582 134000 231638 134056
rect 231766 133048 231822 133104
rect 231674 132504 231730 132560
rect 231766 132096 231822 132152
rect 231674 131552 231730 131608
rect 231582 131144 231638 131200
rect 231490 130192 231546 130248
rect 231674 129240 231730 129296
rect 231766 128832 231822 128888
rect 231674 128288 231730 128344
rect 231766 127880 231822 127936
rect 231582 127336 231638 127392
rect 231674 126928 231730 126984
rect 231766 126384 231822 126440
rect 231582 125976 231638 126032
rect 231766 125432 231822 125488
rect 231306 125024 231362 125080
rect 231766 123528 231822 123584
rect 231398 121624 231454 121680
rect 231490 121216 231546 121272
rect 231398 120264 231454 120320
rect 231766 122576 231822 122632
rect 231766 120672 231822 120728
rect 231766 119720 231822 119776
rect 231582 119312 231638 119368
rect 231490 116456 231546 116512
rect 231766 117952 231822 118008
rect 231766 117000 231822 117056
rect 231674 116048 231730 116104
rect 231766 115504 231822 115560
rect 231306 114552 231362 114608
rect 231490 113600 231546 113656
rect 231766 113192 231822 113248
rect 231214 106528 231270 106584
rect 231122 100816 231178 100872
rect 230846 99456 230902 99512
rect 231030 98912 231086 98968
rect 231766 112648 231822 112704
rect 231674 112240 231730 112296
rect 231766 111716 231822 111752
rect 231766 111696 231768 111716
rect 231768 111696 231820 111716
rect 231820 111696 231822 111716
rect 231582 111288 231638 111344
rect 231490 110744 231546 110800
rect 231766 110372 231768 110392
rect 231768 110372 231820 110392
rect 231820 110372 231822 110392
rect 231766 110336 231822 110372
rect 231766 109420 231768 109440
rect 231768 109420 231820 109440
rect 231820 109420 231822 109440
rect 231766 109384 231822 109420
rect 231674 108876 231676 108896
rect 231676 108876 231728 108896
rect 231728 108876 231730 108896
rect 231674 108840 231730 108876
rect 231766 108432 231822 108488
rect 231766 107480 231822 107536
rect 231490 107072 231546 107128
rect 231766 106156 231768 106176
rect 231768 106156 231820 106176
rect 231820 106156 231822 106176
rect 231766 106120 231822 106156
rect 231674 105168 231730 105224
rect 231766 103672 231822 103728
rect 231766 103264 231822 103320
rect 231490 102312 231546 102368
rect 231766 101360 231822 101416
rect 231674 100408 231730 100464
rect 231766 99900 231768 99920
rect 231768 99900 231820 99920
rect 231820 99900 231822 99920
rect 231766 99864 231822 99900
rect 231306 98504 231362 98560
rect 230754 97960 230810 98016
rect 230754 97008 230810 97064
rect 230662 96600 230718 96656
rect 230570 95784 230626 95840
rect 231582 97588 231584 97608
rect 231584 97588 231636 97608
rect 231636 97588 231638 97608
rect 231582 97552 231638 97588
rect 231766 97008 231822 97064
rect 231306 96600 231362 96656
rect 243910 239944 243966 240000
rect 244186 241848 244242 241904
rect 244646 273672 244702 273728
rect 244554 273128 244610 273184
rect 244738 270136 244794 270192
rect 244830 264424 244886 264480
rect 246026 284824 246082 284880
rect 245658 283736 245714 283792
rect 245198 283192 245254 283248
rect 245014 262248 245070 262304
rect 244922 260616 244978 260672
rect 244922 255176 244978 255232
rect 245106 260888 245162 260944
rect 245842 282376 245898 282432
rect 245658 281016 245714 281072
rect 245658 279384 245714 279440
rect 245750 275884 245752 275904
rect 245752 275884 245804 275904
rect 245804 275884 245806 275904
rect 245750 275848 245806 275884
rect 245750 274488 245806 274544
rect 245750 272312 245806 272368
rect 245750 269592 245806 269648
rect 245658 268776 245714 268832
rect 245750 267960 245806 268016
rect 245750 267416 245806 267472
rect 245750 265784 245806 265840
rect 245750 265104 245806 265160
rect 245658 263880 245714 263936
rect 245750 263064 245806 263120
rect 245658 261704 245714 261760
rect 245934 281560 245990 281616
rect 245934 280220 245990 280256
rect 245934 280200 245936 280220
rect 245936 280200 245988 280220
rect 245988 280200 245990 280220
rect 245934 266600 245990 266656
rect 245934 259528 245990 259584
rect 245750 258712 245806 258768
rect 245750 256536 245806 256592
rect 245658 252456 245714 252512
rect 245750 248648 245806 248704
rect 245658 247288 245714 247344
rect 245658 242936 245714 242992
rect 245658 241576 245714 241632
rect 245290 239944 245346 240000
rect 246118 275304 246174 275360
rect 246118 265240 246174 265296
rect 246118 265104 246174 265160
rect 246026 255992 246082 256048
rect 246026 253816 246082 253872
rect 246026 251640 246082 251696
rect 246026 250280 246082 250336
rect 246026 248140 246028 248160
rect 246028 248140 246080 248160
rect 246080 248140 246082 248160
rect 246026 248104 246082 248140
rect 246026 246472 246082 246528
rect 246026 245928 246082 245984
rect 246026 243752 246082 243808
rect 246026 240216 246082 240272
rect 246302 276664 246358 276720
rect 246210 254360 246266 254416
rect 246394 270952 246450 271008
rect 246486 258188 246542 258224
rect 246486 258168 246488 258188
rect 246488 258168 246540 258188
rect 246540 258168 246542 258188
rect 246670 257352 246726 257408
rect 246578 253000 246634 253056
rect 246486 252184 246542 252240
rect 246394 177520 246450 177576
rect 246854 249464 246910 249520
rect 246670 242392 246726 242448
rect 248418 286184 248474 286240
rect 253294 284280 253350 284336
rect 260194 284552 260250 284608
rect 264426 174392 264482 174448
rect 262954 159840 263010 159896
rect 261574 141888 261630 141944
rect 262586 135768 262642 135824
rect 261666 100544 261722 100600
rect 265254 171944 265310 172000
rect 265438 171536 265494 171592
rect 265530 171148 265586 171184
rect 265530 171128 265532 171148
rect 265532 171128 265584 171148
rect 265584 171128 265586 171148
rect 265530 170584 265586 170640
rect 265162 170176 265218 170232
rect 265346 167592 265402 167648
rect 265162 167048 265218 167104
rect 265438 165960 265494 166016
rect 264426 165688 264482 165744
rect 264242 140120 264298 140176
rect 264150 126792 264206 126848
rect 264334 130192 264390 130248
rect 265438 165008 265494 165064
rect 265162 163784 265218 163840
rect 264702 163376 264758 163432
rect 264518 153040 264574 153096
rect 264518 135904 264574 135960
rect 264518 133728 264574 133784
rect 264518 131960 264574 132016
rect 264426 122576 264482 122632
rect 264426 122032 264482 122088
rect 265438 162016 265494 162072
rect 265530 160112 265586 160168
rect 265438 159024 265494 159080
rect 265346 158752 265402 158808
rect 265162 157800 265218 157856
rect 265438 155624 265494 155680
rect 265530 155216 265586 155272
rect 265530 153856 265586 153912
rect 265254 152632 265310 152688
rect 265346 150864 265402 150920
rect 265070 150476 265126 150512
rect 265070 150456 265072 150476
rect 265072 150456 265124 150476
rect 265124 150456 265126 150476
rect 265346 150048 265402 150104
rect 265530 149640 265586 149696
rect 265254 147872 265310 147928
rect 265530 147056 265586 147112
rect 265346 146104 265402 146160
rect 265162 145288 265218 145344
rect 265346 144472 265402 144528
rect 265530 143520 265586 143576
rect 265162 143112 265218 143168
rect 265438 138352 265494 138408
rect 265530 138100 265586 138136
rect 265530 138080 265532 138100
rect 265532 138080 265584 138100
rect 265584 138080 265586 138100
rect 265438 137536 265494 137592
rect 265530 137128 265586 137184
rect 265254 136312 265310 136368
rect 265254 134544 265310 134600
rect 265162 132776 265218 132832
rect 265530 129376 265586 129432
rect 265346 128968 265402 129024
rect 265530 127200 265586 127256
rect 265530 125568 265586 125624
rect 265162 124616 265218 124672
rect 265346 124244 265348 124264
rect 265348 124244 265400 124264
rect 265400 124244 265402 124264
rect 265346 124208 265402 124244
rect 265438 123392 265494 123448
rect 265162 123004 265218 123040
rect 265162 122984 265164 123004
rect 265164 122984 265216 123004
rect 265216 122984 265218 123004
rect 265530 121624 265586 121680
rect 264702 121216 264758 121272
rect 265530 120808 265586 120864
rect 265438 120148 265494 120184
rect 265438 120128 265440 120148
rect 265440 120128 265492 120148
rect 265492 120128 265494 120148
rect 265530 119040 265586 119096
rect 265438 118788 265494 118824
rect 265438 118768 265440 118788
rect 265440 118768 265492 118788
rect 265492 118768 265494 118788
rect 265530 118224 265586 118280
rect 264610 115912 264666 115968
rect 265530 112240 265586 112296
rect 265162 110880 265218 110936
rect 265346 109248 265402 109304
rect 264610 108704 264666 108760
rect 265530 108296 265586 108352
rect 265438 107072 265494 107128
rect 265438 105304 265494 105360
rect 264794 104896 264850 104952
rect 264702 103128 264758 103184
rect 265346 104488 265402 104544
rect 265162 103944 265218 104000
rect 265438 102720 265494 102776
rect 265530 100952 265586 101008
rect 265530 99476 265586 99512
rect 265530 99456 265532 99476
rect 265532 99456 265584 99476
rect 265584 99456 265586 99476
rect 265714 285776 265770 285832
rect 265898 175344 265954 175400
rect 266082 174936 266138 174992
rect 265990 174528 266046 174584
rect 265806 174120 265862 174176
rect 265990 173712 266046 173768
rect 265898 173304 265954 173360
rect 265806 172760 265862 172816
rect 265806 169768 265862 169824
rect 265898 169360 265954 169416
rect 265806 168544 265862 168600
rect 265990 168952 266046 169008
rect 265898 168408 265954 168464
rect 265806 167184 265862 167240
rect 265806 166368 265862 166424
rect 265898 164600 265954 164656
rect 265806 164192 265862 164248
rect 265806 162988 265862 163024
rect 265806 162968 265808 162988
rect 265808 162968 265860 162988
rect 265860 162968 265862 162988
rect 265806 161608 265862 161664
rect 265990 160792 266046 160848
rect 265898 160384 265954 160440
rect 265898 159432 265954 159488
rect 265898 158208 265954 158264
rect 266266 161472 266322 161528
rect 265806 157412 265862 157448
rect 265806 157392 265808 157412
rect 265808 157392 265860 157412
rect 265860 157392 265862 157412
rect 265898 156848 265954 156904
rect 265806 156440 265862 156496
rect 266082 156032 266138 156088
rect 265806 154808 265862 154864
rect 265990 154672 266046 154728
rect 265806 153448 265862 153504
rect 265898 152088 265954 152144
rect 265806 151836 265862 151872
rect 265806 151816 265808 151836
rect 265808 151816 265860 151836
rect 265860 151816 265862 151836
rect 265806 151272 265862 151328
rect 265806 149232 265862 149288
rect 265898 148280 265954 148336
rect 265898 146648 265954 146704
rect 265806 146512 265862 146568
rect 265898 145696 265954 145752
rect 265806 144880 265862 144936
rect 265806 144064 265862 144120
rect 266082 148688 266138 148744
rect 266174 142704 266230 142760
rect 266082 142296 266138 142352
rect 265806 141344 265862 141400
rect 265898 140936 265954 140992
rect 265990 140800 266046 140856
rect 265898 139712 265954 139768
rect 265806 139460 265862 139496
rect 265806 139440 265808 139460
rect 265808 139440 265860 139460
rect 265860 139440 265862 139460
rect 265990 138760 266046 138816
rect 265990 136740 266046 136776
rect 265990 136720 265992 136740
rect 265992 136720 266044 136740
rect 266044 136720 266046 136740
rect 265990 135360 266046 135416
rect 265990 134136 266046 134192
rect 265990 132540 265992 132560
rect 265992 132540 266044 132560
rect 266044 132540 266046 132560
rect 265990 132504 266046 132540
rect 265990 131552 266046 131608
rect 265990 129784 266046 129840
rect 265990 128560 266046 128616
rect 265898 117816 265954 117872
rect 265806 117408 265862 117464
rect 265898 116456 265954 116512
rect 265806 116084 265808 116104
rect 265808 116084 265860 116104
rect 265860 116084 265862 116104
rect 265806 116048 265862 116084
rect 265898 115232 265954 115288
rect 265806 114688 265862 114744
rect 265898 113872 265954 113928
rect 265806 113464 265862 113520
rect 265806 113212 265862 113248
rect 265806 113192 265808 113212
rect 265808 113192 265860 113212
rect 265860 113192 265862 113212
rect 265898 112648 265954 112704
rect 265806 112104 265862 112160
rect 265898 111288 265954 111344
rect 265806 110508 265808 110528
rect 265808 110508 265860 110528
rect 265860 110508 265862 110528
rect 265806 110472 265862 110508
rect 265898 110064 265954 110120
rect 265806 109656 265862 109712
rect 265806 107908 265862 107944
rect 265806 107888 265808 107908
rect 265808 107888 265860 107908
rect 265860 107888 265862 107908
rect 265806 107616 265862 107672
rect 265806 106664 265862 106720
rect 265898 106528 265954 106584
rect 265806 105712 265862 105768
rect 265806 103572 265808 103592
rect 265808 103572 265860 103592
rect 265860 103572 265862 103592
rect 265806 103536 265862 103572
rect 265806 102312 265862 102368
rect 265898 101360 265954 101416
rect 265806 100816 265862 100872
rect 265898 100136 265954 100192
rect 265806 99728 265862 99784
rect 265714 98776 265770 98832
rect 266174 133184 266230 133240
rect 266174 131180 266176 131200
rect 266176 131180 266228 131200
rect 266228 131180 266230 131200
rect 266174 131144 266230 131180
rect 266174 130600 266230 130656
rect 266174 128424 266230 128480
rect 266174 127608 266230 127664
rect 266174 126384 266230 126440
rect 266266 125976 266322 126032
rect 266174 125024 266230 125080
rect 266174 123800 266230 123856
rect 266174 120400 266230 120456
rect 266174 119448 266230 119504
rect 266082 116864 266138 116920
rect 266082 114824 266138 114880
rect 265990 98368 266046 98424
rect 265622 97144 265678 97200
rect 265530 96772 265532 96792
rect 265532 96772 265584 96792
rect 265584 96772 265586 96792
rect 265530 96736 265586 96772
rect 265806 97996 265808 98016
rect 265808 97996 265860 98016
rect 265860 97996 265862 98016
rect 265806 97960 265862 97996
rect 265898 97552 265954 97608
rect 265806 96872 265862 96928
rect 265714 95648 265770 95704
rect 278778 176024 278834 176080
rect 279330 149776 279386 149832
rect 280250 180376 280306 180432
rect 280158 125432 280214 125488
rect 280434 121624 280490 121680
rect 280342 120808 280398 120864
rect 280710 160112 280766 160168
rect 280618 141616 280674 141672
rect 281538 172352 281594 172408
rect 281630 170040 281686 170096
rect 281722 168544 281778 168600
rect 281906 181464 281962 181520
rect 281814 167728 281870 167784
rect 281998 164736 282054 164792
rect 282274 177384 282330 177440
rect 282182 170856 282238 170912
rect 282366 173168 282422 173224
rect 282274 167048 282330 167104
rect 282090 162424 282146 162480
rect 282182 160792 282238 160848
rect 281906 158480 281962 158536
rect 281998 157800 282054 157856
rect 282458 156304 282514 156360
rect 281814 154672 281870 154728
rect 282090 153992 282146 154048
rect 282090 152360 282146 152416
rect 281630 150864 281686 150920
rect 281722 150456 281778 150512
rect 281630 137844 281632 137864
rect 281632 137844 281684 137864
rect 281684 137844 281686 137864
rect 281630 137808 281686 137844
rect 281630 123120 281686 123176
rect 281538 122440 281594 122496
rect 282090 147736 282146 147792
rect 281906 143928 281962 143984
rect 282274 153176 282330 153232
rect 282274 151716 282276 151736
rect 282276 151716 282328 151736
rect 282328 151716 282330 151736
rect 282274 151680 282330 151716
rect 282274 136992 282330 137048
rect 282182 135496 282238 135552
rect 282826 165416 282882 165472
rect 282826 161608 282882 161664
rect 282826 159296 282882 159352
rect 282826 156984 282882 157040
rect 282826 155488 282882 155544
rect 282826 150048 282882 150104
rect 282826 148552 282882 148608
rect 282826 146240 282882 146296
rect 282826 142432 282882 142488
rect 282826 140120 282882 140176
rect 282734 139304 282790 139360
rect 282826 138488 282882 138544
rect 282826 136312 282882 136368
rect 282550 134680 282606 134736
rect 281814 134000 281870 134056
rect 282274 133184 282330 133240
rect 282550 132388 282606 132424
rect 282550 132368 282552 132388
rect 282552 132368 282604 132388
rect 282604 132368 282606 132388
rect 282090 131688 282146 131744
rect 281906 130872 281962 130928
rect 282090 130056 282146 130112
rect 281906 129376 281962 129432
rect 282090 128560 282146 128616
rect 281906 127744 281962 127800
rect 281906 127064 281962 127120
rect 282826 126248 282882 126304
rect 282826 124752 282882 124808
rect 282826 123936 282882 123992
rect 281722 120128 281778 120184
rect 280526 119312 280582 119368
rect 282734 118532 282736 118552
rect 282736 118532 282788 118552
rect 282788 118532 282790 118552
rect 282734 118496 282790 118532
rect 282826 117816 282882 117872
rect 282826 117000 282882 117056
rect 282826 116320 282882 116376
rect 282826 114688 282882 114744
rect 282734 114008 282790 114064
rect 282826 113192 282882 113248
rect 282826 112376 282882 112432
rect 281998 111696 282054 111752
rect 282826 110880 282882 110936
rect 282274 110064 282330 110120
rect 282826 109384 282882 109440
rect 281538 108604 281540 108624
rect 281540 108604 281592 108624
rect 281592 108604 281594 108624
rect 281538 108568 281594 108604
rect 282366 107752 282422 107808
rect 281722 107072 281778 107128
rect 280250 106256 280306 106312
rect 282826 105440 282882 105496
rect 281538 104796 281540 104816
rect 281540 104796 281592 104816
rect 281592 104796 281594 104816
rect 281538 104760 281594 104796
rect 281538 103944 281594 104000
rect 282826 103128 282882 103184
rect 281998 102448 282054 102504
rect 281630 101632 281686 101688
rect 281538 99320 281594 99376
rect 279422 98096 279478 98152
rect 279330 96600 279386 96656
rect 279514 97280 279570 97336
rect 279238 96056 279294 96112
rect 287610 180240 287666 180296
rect 288898 180512 288954 180568
rect 289082 179968 289138 180024
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 580262 590960 580318 591016
rect 579894 564304 579950 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 579986 404912 580042 404968
rect 580170 378392 580226 378448
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 579618 325216 579674 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 579802 245520 579858 245576
rect 580354 577632 580410 577688
rect 580446 365064 580502 365120
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 579986 179152 580042 179208
rect 580170 165824 580226 165880
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 282274 100136 282330 100192
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580262 46280 580318 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580257 591018 580323 591021
rect 583520 591018 584960 591108
rect 580257 591016 584960 591018
rect 580257 590960 580262 591016
rect 580318 590960 584960 591016
rect 580257 590958 584960 590960
rect 580257 590955 580323 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580349 577690 580415 577693
rect 583520 577690 584960 577780
rect 580349 577688 584960 577690
rect 580349 577632 580354 577688
rect 580410 577632 584960 577688
rect 580349 577630 584960 577632
rect 580349 577627 580415 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579889 564362 579955 564365
rect 583520 564362 584960 564452
rect 579889 564360 584960 564362
rect 579889 564304 579894 564360
rect 579950 564304 584960 564360
rect 579889 564302 584960 564304
rect 579889 564299 579955 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3049 475690 3115 475693
rect -960 475688 3115 475690
rect -960 475632 3054 475688
rect 3110 475632 3115 475688
rect -960 475630 3115 475632
rect -960 475540 480 475630
rect 3049 475627 3115 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3601 410546 3667 410549
rect -960 410544 3667 410546
rect -960 410488 3606 410544
rect 3662 410488 3667 410544
rect -960 410486 3667 410488
rect -960 410396 480 410486
rect 3601 410483 3667 410486
rect 579981 404970 580047 404973
rect 583520 404970 584960 405060
rect 579981 404968 584960 404970
rect 579981 404912 579986 404968
rect 580042 404912 584960 404968
rect 579981 404910 584960 404912
rect 579981 404907 580047 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580441 365122 580507 365125
rect 583520 365122 584960 365212
rect 580441 365120 584960 365122
rect 580441 365064 580446 365120
rect 580502 365064 584960 365120
rect 580441 365062 584960 365064
rect 580441 365059 580507 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579613 325274 579679 325277
rect 583520 325274 584960 325364
rect 579613 325272 584960 325274
rect 579613 325216 579618 325272
rect 579674 325216 584960 325272
rect 579613 325214 584960 325216
rect 579613 325211 579679 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3049 306234 3115 306237
rect -960 306232 3115 306234
rect -960 306176 3054 306232
rect 3110 306176 3115 306232
rect -960 306174 3115 306176
rect -960 306084 480 306174
rect 3049 306171 3115 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 226885 286242 226951 286245
rect 248413 286242 248479 286245
rect 226885 286240 248479 286242
rect 226885 286184 226890 286240
rect 226946 286184 248418 286240
rect 248474 286184 248479 286240
rect 226885 286182 248479 286184
rect 226885 286179 226951 286182
rect 248413 286179 248479 286182
rect 221549 286106 221615 286109
rect 280654 286106 280660 286108
rect 221549 286104 280660 286106
rect 221549 286048 221554 286104
rect 221610 286048 280660 286104
rect 221549 286046 280660 286048
rect 221549 286043 221615 286046
rect 280654 286044 280660 286046
rect 280724 286044 280730 286108
rect 221181 285970 221247 285973
rect 285622 285970 285628 285972
rect 221181 285968 285628 285970
rect 221181 285912 221186 285968
rect 221242 285912 285628 285968
rect 221181 285910 285628 285912
rect 221181 285907 221247 285910
rect 285622 285908 285628 285910
rect 285692 285908 285698 285972
rect 200757 285834 200823 285837
rect 265709 285834 265775 285837
rect 200757 285832 265775 285834
rect 200757 285776 200762 285832
rect 200818 285776 265714 285832
rect 265770 285776 265775 285832
rect 200757 285774 265775 285776
rect 200757 285771 200823 285774
rect 265709 285771 265775 285774
rect 215845 285698 215911 285701
rect 284334 285698 284340 285700
rect 215845 285696 284340 285698
rect 215845 285640 215850 285696
rect 215906 285640 284340 285696
rect 215845 285638 284340 285640
rect 215845 285635 215911 285638
rect 284334 285636 284340 285638
rect 284404 285636 284410 285700
rect 583520 285276 584960 285516
rect 240777 284882 240843 284885
rect 246021 284882 246087 284885
rect 240777 284880 246087 284882
rect 240777 284824 240782 284880
rect 240838 284824 246026 284880
rect 246082 284824 246087 284880
rect 240777 284822 246087 284824
rect 240777 284819 240843 284822
rect 246021 284819 246087 284822
rect 206645 284746 206711 284749
rect 287646 284746 287652 284748
rect 206645 284744 287652 284746
rect 206645 284688 206650 284744
rect 206706 284688 287652 284744
rect 206645 284686 287652 284688
rect 206645 284683 206711 284686
rect 287646 284684 287652 284686
rect 287716 284684 287722 284748
rect 233693 284610 233759 284613
rect 260189 284610 260255 284613
rect 233693 284608 260255 284610
rect 233693 284552 233698 284608
rect 233754 284552 260194 284608
rect 260250 284552 260255 284608
rect 233693 284550 260255 284552
rect 233693 284547 233759 284550
rect 260189 284547 260255 284550
rect 219709 284474 219775 284477
rect 278814 284474 278820 284476
rect 219709 284472 278820 284474
rect 219709 284416 219714 284472
rect 219770 284416 278820 284472
rect 219709 284414 278820 284416
rect 219709 284411 219775 284414
rect 278814 284412 278820 284414
rect 278884 284412 278890 284476
rect 239029 284338 239095 284341
rect 253289 284338 253355 284341
rect 239029 284336 253355 284338
rect 239029 284280 239034 284336
rect 239090 284280 253294 284336
rect 253350 284280 253355 284336
rect 239029 284278 253355 284280
rect 239029 284275 239095 284278
rect 253289 284275 253355 284278
rect 243353 284068 243419 284069
rect 243302 284066 243308 284068
rect 243262 284006 243308 284066
rect 243372 284064 243419 284068
rect 243414 284008 243419 284064
rect 243302 284004 243308 284006
rect 243372 284004 243419 284008
rect 243353 284003 243419 284004
rect 198641 283794 198707 283797
rect 245653 283794 245719 283797
rect 198641 283792 200284 283794
rect 198641 283736 198646 283792
rect 198702 283736 200284 283792
rect 198641 283734 200284 283736
rect 244076 283792 245719 283794
rect 244076 283736 245658 283792
rect 245714 283736 245719 283792
rect 244076 283734 245719 283736
rect 198641 283731 198707 283734
rect 245653 283731 245719 283734
rect 245193 283250 245259 283253
rect 244076 283248 245259 283250
rect 244076 283192 245198 283248
rect 245254 283192 245259 283248
rect 244076 283190 245259 283192
rect 245193 283187 245259 283190
rect 198273 282978 198339 282981
rect 198273 282976 200284 282978
rect 198273 282920 198278 282976
rect 198334 282920 200284 282976
rect 198273 282918 200284 282920
rect 198273 282915 198339 282918
rect 199561 282434 199627 282437
rect 245837 282434 245903 282437
rect 199561 282432 200284 282434
rect 199561 282376 199566 282432
rect 199622 282376 200284 282432
rect 199561 282374 200284 282376
rect 244076 282432 245903 282434
rect 244076 282376 245842 282432
rect 245898 282376 245903 282432
rect 244076 282374 245903 282376
rect 199561 282371 199627 282374
rect 245837 282371 245903 282374
rect 197353 281618 197419 281621
rect 245929 281618 245995 281621
rect 197353 281616 200284 281618
rect 197353 281560 197358 281616
rect 197414 281560 200284 281616
rect 197353 281558 200284 281560
rect 244076 281616 245995 281618
rect 244076 281560 245934 281616
rect 245990 281560 245995 281616
rect 244076 281558 245995 281560
rect 197353 281555 197419 281558
rect 245929 281555 245995 281558
rect 245653 281074 245719 281077
rect 244076 281072 245719 281074
rect 244076 281016 245658 281072
rect 245714 281016 245719 281072
rect 244076 281014 245719 281016
rect 245653 281011 245719 281014
rect 198549 280802 198615 280805
rect 198549 280800 200284 280802
rect 198549 280744 198554 280800
rect 198610 280744 200284 280800
rect 198549 280742 200284 280744
rect 198549 280739 198615 280742
rect 197353 280258 197419 280261
rect 245929 280258 245995 280261
rect 197353 280256 200284 280258
rect -960 279972 480 280212
rect 197353 280200 197358 280256
rect 197414 280200 200284 280256
rect 197353 280198 200284 280200
rect 244076 280256 245995 280258
rect 244076 280200 245934 280256
rect 245990 280200 245995 280256
rect 244076 280198 245995 280200
rect 197353 280195 197419 280198
rect 245929 280195 245995 280198
rect 197353 279442 197419 279445
rect 245653 279442 245719 279445
rect 197353 279440 200284 279442
rect 197353 279384 197358 279440
rect 197414 279384 200284 279440
rect 197353 279382 200284 279384
rect 244076 279440 245719 279442
rect 244076 279384 245658 279440
rect 245714 279384 245719 279440
rect 244076 279382 245719 279384
rect 197353 279379 197419 279382
rect 245653 279379 245719 279382
rect 244273 278898 244339 278901
rect 244076 278896 244339 278898
rect 244076 278840 244278 278896
rect 244334 278840 244339 278896
rect 244076 278838 244339 278840
rect 244273 278835 244339 278838
rect 199469 278626 199535 278629
rect 199469 278624 200284 278626
rect 199469 278568 199474 278624
rect 199530 278568 200284 278624
rect 199469 278566 200284 278568
rect 199469 278563 199535 278566
rect 198641 278082 198707 278085
rect 244365 278082 244431 278085
rect 198641 278080 200284 278082
rect 198641 278024 198646 278080
rect 198702 278024 200284 278080
rect 198641 278022 200284 278024
rect 244076 278080 244431 278082
rect 244076 278024 244370 278080
rect 244426 278024 244431 278080
rect 244076 278022 244431 278024
rect 198641 278019 198707 278022
rect 244365 278019 244431 278022
rect 288934 277538 288940 277540
rect 244076 277478 288940 277538
rect 288934 277476 288940 277478
rect 289004 277476 289010 277540
rect 197445 277266 197511 277269
rect 197445 277264 200284 277266
rect 197445 277208 197450 277264
rect 197506 277208 200284 277264
rect 197445 277206 200284 277208
rect 197445 277203 197511 277206
rect 199653 276722 199719 276725
rect 246297 276722 246363 276725
rect 199653 276720 200284 276722
rect 199653 276664 199658 276720
rect 199714 276664 200284 276720
rect 199653 276662 200284 276664
rect 244076 276720 246363 276722
rect 244076 276664 246302 276720
rect 246358 276664 246363 276720
rect 244076 276662 246363 276664
rect 199653 276659 199719 276662
rect 246297 276659 246363 276662
rect 197353 275906 197419 275909
rect 245745 275906 245811 275909
rect 197353 275904 200284 275906
rect 197353 275848 197358 275904
rect 197414 275848 200284 275904
rect 197353 275846 200284 275848
rect 244076 275904 245811 275906
rect 244076 275848 245750 275904
rect 245806 275848 245811 275904
rect 244076 275846 245811 275848
rect 197353 275843 197419 275846
rect 245745 275843 245811 275846
rect 246113 275362 246179 275365
rect 244076 275360 246179 275362
rect 244076 275304 246118 275360
rect 246174 275304 246179 275360
rect 244076 275302 246179 275304
rect 246113 275299 246179 275302
rect 199745 275090 199811 275093
rect 199745 275088 200284 275090
rect 199745 275032 199750 275088
rect 199806 275032 200284 275088
rect 199745 275030 200284 275032
rect 199745 275027 199811 275030
rect 198181 274546 198247 274549
rect 245745 274546 245811 274549
rect 198181 274544 200284 274546
rect 198181 274488 198186 274544
rect 198242 274488 200284 274544
rect 198181 274486 200284 274488
rect 244076 274544 245811 274546
rect 244076 274488 245750 274544
rect 245806 274488 245811 274544
rect 244076 274486 245811 274488
rect 198181 274483 198247 274486
rect 245745 274483 245811 274486
rect 200021 273730 200087 273733
rect 244641 273730 244707 273733
rect 200021 273728 200284 273730
rect 200021 273672 200026 273728
rect 200082 273672 200284 273728
rect 200021 273670 200284 273672
rect 244076 273728 244707 273730
rect 244076 273672 244646 273728
rect 244702 273672 244707 273728
rect 244076 273670 244707 273672
rect 200021 273667 200087 273670
rect 244641 273667 244707 273670
rect 244549 273186 244615 273189
rect 244076 273184 244615 273186
rect 244076 273128 244554 273184
rect 244610 273128 244615 273184
rect 244076 273126 244615 273128
rect 244549 273123 244615 273126
rect 197445 272914 197511 272917
rect 197445 272912 200284 272914
rect 197445 272856 197450 272912
rect 197506 272856 200284 272912
rect 197445 272854 200284 272856
rect 197445 272851 197511 272854
rect 197353 272370 197419 272373
rect 245745 272370 245811 272373
rect 197353 272368 200284 272370
rect 197353 272312 197358 272368
rect 197414 272312 200284 272368
rect 197353 272310 200284 272312
rect 244076 272368 245811 272370
rect 244076 272312 245750 272368
rect 245806 272312 245811 272368
rect 244076 272310 245811 272312
rect 197353 272307 197419 272310
rect 245745 272307 245811 272310
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 199929 271554 199995 271557
rect 244365 271554 244431 271557
rect 199929 271552 200284 271554
rect 199929 271496 199934 271552
rect 199990 271496 200284 271552
rect 199929 271494 200284 271496
rect 244076 271552 244431 271554
rect 244076 271496 244370 271552
rect 244426 271496 244431 271552
rect 244076 271494 244431 271496
rect 199929 271491 199995 271494
rect 244365 271491 244431 271494
rect 198549 271010 198615 271013
rect 246389 271010 246455 271013
rect 198549 271008 200284 271010
rect 198549 270952 198554 271008
rect 198610 270952 200284 271008
rect 198549 270950 200284 270952
rect 244076 271008 246455 271010
rect 244076 270952 246394 271008
rect 246450 270952 246455 271008
rect 244076 270950 246455 270952
rect 198549 270947 198615 270950
rect 246389 270947 246455 270950
rect 199837 270194 199903 270197
rect 244733 270194 244799 270197
rect 199837 270192 200284 270194
rect 199837 270136 199842 270192
rect 199898 270136 200284 270192
rect 199837 270134 200284 270136
rect 244076 270192 244799 270194
rect 244076 270136 244738 270192
rect 244794 270136 244799 270192
rect 244076 270134 244799 270136
rect 199837 270131 199903 270134
rect 244733 270131 244799 270134
rect 245745 269650 245811 269653
rect 244076 269648 245811 269650
rect 244076 269592 245750 269648
rect 245806 269592 245811 269648
rect 244076 269590 245811 269592
rect 245745 269587 245811 269590
rect 197353 269378 197419 269381
rect 197353 269376 200284 269378
rect 197353 269320 197358 269376
rect 197414 269320 200284 269376
rect 197353 269318 200284 269320
rect 197353 269315 197419 269318
rect 197445 268834 197511 268837
rect 245653 268834 245719 268837
rect 197445 268832 200284 268834
rect 197445 268776 197450 268832
rect 197506 268776 200284 268832
rect 197445 268774 200284 268776
rect 244076 268832 245719 268834
rect 244076 268776 245658 268832
rect 245714 268776 245719 268832
rect 244076 268774 245719 268776
rect 197445 268771 197511 268774
rect 245653 268771 245719 268774
rect 197353 268018 197419 268021
rect 245745 268018 245811 268021
rect 197353 268016 200284 268018
rect 197353 267960 197358 268016
rect 197414 267960 200284 268016
rect 197353 267958 200284 267960
rect 244076 268016 245811 268018
rect 244076 267960 245750 268016
rect 245806 267960 245811 268016
rect 244076 267958 245811 267960
rect 197353 267955 197419 267958
rect 245745 267955 245811 267958
rect 245745 267474 245811 267477
rect 244076 267472 245811 267474
rect 244076 267416 245750 267472
rect 245806 267416 245811 267472
rect 244076 267414 245811 267416
rect 245745 267411 245811 267414
rect -960 267202 480 267292
rect 3325 267202 3391 267205
rect -960 267200 3391 267202
rect -960 267144 3330 267200
rect 3386 267144 3391 267200
rect -960 267142 3391 267144
rect -960 267052 480 267142
rect 3325 267139 3391 267142
rect 197445 267202 197511 267205
rect 197445 267200 200284 267202
rect 197445 267144 197450 267200
rect 197506 267144 200284 267200
rect 197445 267142 200284 267144
rect 197445 267139 197511 267142
rect 197353 266658 197419 266661
rect 245929 266658 245995 266661
rect 197353 266656 200284 266658
rect 197353 266600 197358 266656
rect 197414 266600 200284 266656
rect 197353 266598 200284 266600
rect 244076 266656 245995 266658
rect 244076 266600 245934 266656
rect 245990 266600 245995 266656
rect 244076 266598 245995 266600
rect 197353 266595 197419 266598
rect 245929 266595 245995 266598
rect 197445 265842 197511 265845
rect 245745 265842 245811 265845
rect 197445 265840 200284 265842
rect 197445 265784 197450 265840
rect 197506 265784 200284 265840
rect 197445 265782 200284 265784
rect 244076 265840 245811 265842
rect 244076 265784 245750 265840
rect 245806 265784 245811 265840
rect 244076 265782 245811 265784
rect 197445 265779 197511 265782
rect 245745 265779 245811 265782
rect 197353 265298 197419 265301
rect 246113 265298 246179 265301
rect 197353 265296 200284 265298
rect 197353 265240 197358 265296
rect 197414 265240 200284 265296
rect 197353 265238 200284 265240
rect 244076 265296 246179 265298
rect 244076 265240 246118 265296
rect 246174 265240 246179 265296
rect 244076 265238 246179 265240
rect 197353 265235 197419 265238
rect 246113 265235 246179 265238
rect 245745 265162 245811 265165
rect 246113 265162 246179 265165
rect 245745 265160 246179 265162
rect 245745 265104 245750 265160
rect 245806 265104 246118 265160
rect 246174 265104 246179 265160
rect 245745 265102 246179 265104
rect 245745 265099 245811 265102
rect 246113 265099 246179 265102
rect 197353 264482 197419 264485
rect 244825 264482 244891 264485
rect 197353 264480 200284 264482
rect 197353 264424 197358 264480
rect 197414 264424 200284 264480
rect 197353 264422 200284 264424
rect 244076 264480 244891 264482
rect 244076 264424 244830 264480
rect 244886 264424 244891 264480
rect 244076 264422 244891 264424
rect 197353 264419 197419 264422
rect 244825 264419 244891 264422
rect 245653 263938 245719 263941
rect 244076 263936 245719 263938
rect 244076 263880 245658 263936
rect 245714 263880 245719 263936
rect 244076 263878 245719 263880
rect 245653 263875 245719 263878
rect 197353 263666 197419 263669
rect 197353 263664 200284 263666
rect 197353 263608 197358 263664
rect 197414 263608 200284 263664
rect 197353 263606 200284 263608
rect 197353 263603 197419 263606
rect 198457 263122 198523 263125
rect 245745 263122 245811 263125
rect 198457 263120 200284 263122
rect 198457 263064 198462 263120
rect 198518 263064 200284 263120
rect 198457 263062 200284 263064
rect 244076 263120 245811 263122
rect 244076 263064 245750 263120
rect 245806 263064 245811 263120
rect 244076 263062 245811 263064
rect 198457 263059 198523 263062
rect 245745 263059 245811 263062
rect 199285 262306 199351 262309
rect 245009 262306 245075 262309
rect 199285 262304 200284 262306
rect 199285 262248 199290 262304
rect 199346 262248 200284 262304
rect 199285 262246 200284 262248
rect 244076 262304 245075 262306
rect 244076 262248 245014 262304
rect 245070 262248 245075 262304
rect 244076 262246 245075 262248
rect 199285 262243 199351 262246
rect 245009 262243 245075 262246
rect 245653 261762 245719 261765
rect 244076 261760 245719 261762
rect 244076 261704 245658 261760
rect 245714 261704 245719 261760
rect 244076 261702 245719 261704
rect 245653 261699 245719 261702
rect 197353 261490 197419 261493
rect 197353 261488 200284 261490
rect 197353 261432 197358 261488
rect 197414 261432 200284 261488
rect 197353 261430 200284 261432
rect 197353 261427 197419 261430
rect 199510 260884 199516 260948
rect 199580 260946 199586 260948
rect 245101 260946 245167 260949
rect 199580 260886 200284 260946
rect 244076 260944 245167 260946
rect 244076 260888 245106 260944
rect 245162 260888 245167 260944
rect 244076 260886 245167 260888
rect 199580 260884 199586 260886
rect 245101 260883 245167 260886
rect 244917 260674 244983 260677
rect 244046 260672 244983 260674
rect 244046 260616 244922 260672
rect 244978 260616 244983 260672
rect 244046 260614 244983 260616
rect 199377 260130 199443 260133
rect 199377 260128 200284 260130
rect 199377 260072 199382 260128
rect 199438 260072 200284 260128
rect 244046 260100 244106 260614
rect 244917 260611 244983 260614
rect 199377 260070 200284 260072
rect 199377 260067 199443 260070
rect 245929 259586 245995 259589
rect 244076 259584 245995 259586
rect 244076 259528 245934 259584
rect 245990 259528 245995 259584
rect 244076 259526 245995 259528
rect 245929 259523 245995 259526
rect 197445 259314 197511 259317
rect 197445 259312 200284 259314
rect 197445 259256 197450 259312
rect 197506 259256 200284 259312
rect 197445 259254 200284 259256
rect 197445 259251 197511 259254
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 197353 258770 197419 258773
rect 245745 258770 245811 258773
rect 197353 258768 200284 258770
rect 197353 258712 197358 258768
rect 197414 258712 200284 258768
rect 197353 258710 200284 258712
rect 244076 258768 245811 258770
rect 244076 258712 245750 258768
rect 245806 258712 245811 258768
rect 583520 258756 584960 258846
rect 244076 258710 245811 258712
rect 197353 258707 197419 258710
rect 245745 258707 245811 258710
rect 246481 258226 246547 258229
rect 244076 258224 246547 258226
rect 244076 258168 246486 258224
rect 246542 258168 246547 258224
rect 244076 258166 246547 258168
rect 246481 258163 246547 258166
rect 197353 257954 197419 257957
rect 197353 257952 200284 257954
rect 197353 257896 197358 257952
rect 197414 257896 200284 257952
rect 197353 257894 200284 257896
rect 197353 257891 197419 257894
rect 196801 257410 196867 257413
rect 246665 257410 246731 257413
rect 196801 257408 200284 257410
rect 196801 257352 196806 257408
rect 196862 257352 200284 257408
rect 196801 257350 200284 257352
rect 244076 257408 246731 257410
rect 244076 257352 246670 257408
rect 246726 257352 246731 257408
rect 244076 257350 246731 257352
rect 196801 257347 196867 257350
rect 246665 257347 246731 257350
rect 198089 256594 198155 256597
rect 245745 256594 245811 256597
rect 198089 256592 200284 256594
rect 198089 256536 198094 256592
rect 198150 256536 200284 256592
rect 198089 256534 200284 256536
rect 244076 256592 245811 256594
rect 244076 256536 245750 256592
rect 245806 256536 245811 256592
rect 244076 256534 245811 256536
rect 198089 256531 198155 256534
rect 245745 256531 245811 256534
rect 246021 256050 246087 256053
rect 244076 256048 246087 256050
rect 244076 255992 246026 256048
rect 246082 255992 246087 256048
rect 244076 255990 246087 255992
rect 246021 255987 246087 255990
rect 198365 255778 198431 255781
rect 198365 255776 200284 255778
rect 198365 255720 198370 255776
rect 198426 255720 200284 255776
rect 198365 255718 200284 255720
rect 198365 255715 198431 255718
rect 197445 255234 197511 255237
rect 244917 255234 244983 255237
rect 197445 255232 200284 255234
rect 197445 255176 197450 255232
rect 197506 255176 200284 255232
rect 197445 255174 200284 255176
rect 244076 255232 244983 255234
rect 244076 255176 244922 255232
rect 244978 255176 244983 255232
rect 244076 255174 244983 255176
rect 197445 255171 197511 255174
rect 244917 255171 244983 255174
rect 197353 254418 197419 254421
rect 246205 254418 246271 254421
rect 197353 254416 200284 254418
rect 197353 254360 197358 254416
rect 197414 254360 200284 254416
rect 197353 254358 200284 254360
rect 244076 254416 246271 254418
rect 244076 254360 246210 254416
rect 246266 254360 246271 254416
rect 244076 254358 246271 254360
rect 197353 254355 197419 254358
rect 246205 254355 246271 254358
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 246021 253874 246087 253877
rect 244076 253872 246087 253874
rect 244076 253816 246026 253872
rect 246082 253816 246087 253872
rect 244076 253814 246087 253816
rect 246021 253811 246087 253814
rect 197721 253602 197787 253605
rect 197721 253600 200284 253602
rect 197721 253544 197726 253600
rect 197782 253544 200284 253600
rect 197721 253542 200284 253544
rect 197721 253539 197787 253542
rect 197353 253058 197419 253061
rect 246573 253058 246639 253061
rect 197353 253056 200284 253058
rect 197353 253000 197358 253056
rect 197414 253000 200284 253056
rect 197353 252998 200284 253000
rect 244076 253056 246639 253058
rect 244076 253000 246578 253056
rect 246634 253000 246639 253056
rect 244076 252998 246639 253000
rect 197353 252995 197419 252998
rect 246573 252995 246639 252998
rect 244038 252452 244044 252516
rect 244108 252514 244114 252516
rect 245653 252514 245719 252517
rect 244108 252512 245719 252514
rect 244108 252456 245658 252512
rect 245714 252456 245719 252512
rect 244108 252454 245719 252456
rect 244108 252452 244114 252454
rect 245653 252451 245719 252454
rect 198365 252242 198431 252245
rect 246481 252242 246547 252245
rect 198365 252240 200284 252242
rect 198365 252184 198370 252240
rect 198426 252184 200284 252240
rect 198365 252182 200284 252184
rect 244076 252240 246547 252242
rect 244076 252184 246486 252240
rect 246542 252184 246547 252240
rect 244076 252182 246547 252184
rect 198365 252179 198431 252182
rect 246481 252179 246547 252182
rect 197905 251698 197971 251701
rect 246021 251698 246087 251701
rect 197905 251696 200284 251698
rect 197905 251640 197910 251696
rect 197966 251640 200284 251696
rect 197905 251638 200284 251640
rect 244076 251696 246087 251698
rect 244076 251640 246026 251696
rect 246082 251640 246087 251696
rect 244076 251638 246087 251640
rect 197905 251635 197971 251638
rect 246021 251635 246087 251638
rect 200622 250340 200682 250852
rect 244046 250613 244106 250852
rect 244046 250608 244155 250613
rect 244046 250552 244094 250608
rect 244150 250552 244155 250608
rect 244046 250550 244155 250552
rect 244089 250547 244155 250550
rect 200614 250276 200620 250340
rect 200684 250276 200690 250340
rect 246021 250338 246087 250341
rect 244076 250336 246087 250338
rect 244076 250280 246026 250336
rect 246082 250280 246087 250336
rect 244076 250278 246087 250280
rect 246021 250275 246087 250278
rect 197353 250066 197419 250069
rect 197353 250064 200284 250066
rect 197353 250008 197358 250064
rect 197414 250008 200284 250064
rect 197353 250006 200284 250008
rect 197353 250003 197419 250006
rect 197629 249522 197695 249525
rect 246849 249522 246915 249525
rect 197629 249520 200284 249522
rect 197629 249464 197634 249520
rect 197690 249464 200284 249520
rect 197629 249462 200284 249464
rect 244076 249520 246915 249522
rect 244076 249464 246854 249520
rect 246910 249464 246915 249520
rect 244076 249462 246915 249464
rect 197629 249459 197695 249462
rect 246849 249459 246915 249462
rect 197537 248706 197603 248709
rect 245745 248706 245811 248709
rect 197537 248704 200284 248706
rect 197537 248648 197542 248704
rect 197598 248648 200284 248704
rect 197537 248646 200284 248648
rect 244076 248704 245811 248706
rect 244076 248648 245750 248704
rect 245806 248648 245811 248704
rect 244076 248646 245811 248648
rect 197537 248643 197603 248646
rect 245745 248643 245811 248646
rect 246021 248162 246087 248165
rect 244076 248160 246087 248162
rect 244076 248104 246026 248160
rect 246082 248104 246087 248160
rect 244076 248102 246087 248104
rect 246021 248099 246087 248102
rect 197997 247890 198063 247893
rect 197997 247888 200284 247890
rect 197997 247832 198002 247888
rect 198058 247832 200284 247888
rect 197997 247830 200284 247832
rect 197997 247827 198063 247830
rect 197261 247346 197327 247349
rect 245653 247346 245719 247349
rect 197261 247344 200284 247346
rect 197261 247288 197266 247344
rect 197322 247288 200284 247344
rect 197261 247286 200284 247288
rect 244076 247344 245719 247346
rect 244076 247288 245658 247344
rect 245714 247288 245719 247344
rect 244076 247286 245719 247288
rect 197261 247283 197327 247286
rect 245653 247283 245719 247286
rect 246021 246530 246087 246533
rect 244076 246528 246087 246530
rect 200806 246260 200866 246500
rect 244076 246472 246026 246528
rect 246082 246472 246087 246528
rect 244076 246470 246087 246472
rect 246021 246467 246087 246470
rect 200798 246196 200804 246260
rect 200868 246196 200874 246260
rect 197353 245986 197419 245989
rect 246021 245986 246087 245989
rect 197353 245984 200284 245986
rect 197353 245928 197358 245984
rect 197414 245928 200284 245984
rect 197353 245926 200284 245928
rect 244076 245984 246087 245986
rect 244076 245928 246026 245984
rect 246082 245928 246087 245984
rect 244076 245926 246087 245928
rect 197353 245923 197419 245926
rect 246021 245923 246087 245926
rect 579797 245578 579863 245581
rect 583520 245578 584960 245668
rect 579797 245576 584960 245578
rect 579797 245520 579802 245576
rect 579858 245520 584960 245576
rect 579797 245518 584960 245520
rect 579797 245515 579863 245518
rect 583520 245428 584960 245518
rect 199193 245170 199259 245173
rect 199193 245168 200284 245170
rect 199193 245112 199198 245168
rect 199254 245112 200284 245168
rect 199193 245110 200284 245112
rect 199193 245107 199259 245110
rect 243494 244900 243554 245140
rect 243486 244836 243492 244900
rect 243556 244836 243562 244900
rect 200798 244564 200804 244628
rect 200868 244564 200874 244628
rect 200806 244324 200866 244564
rect 244046 244357 244106 244596
rect 243997 244352 244106 244357
rect 243997 244296 244002 244352
rect 244058 244296 244106 244352
rect 243997 244294 244106 244296
rect 243997 244291 244063 244294
rect 197353 243810 197419 243813
rect 246021 243810 246087 243813
rect 197353 243808 200284 243810
rect 197353 243752 197358 243808
rect 197414 243752 200284 243808
rect 197353 243750 200284 243752
rect 244076 243808 246087 243810
rect 244076 243752 246026 243808
rect 246082 243752 246087 243808
rect 244076 243750 246087 243752
rect 197353 243747 197419 243750
rect 246021 243747 246087 243750
rect 197445 242994 197511 242997
rect 245653 242994 245719 242997
rect 197445 242992 200284 242994
rect 197445 242936 197450 242992
rect 197506 242936 200284 242992
rect 197445 242934 200284 242936
rect 244076 242992 245719 242994
rect 244076 242936 245658 242992
rect 245714 242936 245719 242992
rect 244076 242934 245719 242936
rect 197445 242931 197511 242934
rect 245653 242931 245719 242934
rect 246665 242450 246731 242453
rect 244076 242448 246731 242450
rect 244076 242392 246670 242448
rect 246726 242392 246731 242448
rect 244076 242390 246731 242392
rect 246665 242387 246731 242390
rect 197997 242178 198063 242181
rect 197997 242176 200284 242178
rect 197997 242120 198002 242176
rect 198058 242120 200284 242176
rect 197997 242118 200284 242120
rect 197997 242115 198063 242118
rect 243670 241844 243676 241908
rect 243740 241906 243746 241908
rect 244181 241906 244247 241909
rect 243740 241904 244247 241906
rect 243740 241848 244186 241904
rect 244242 241848 244247 241904
rect 243740 241846 244247 241848
rect 243740 241844 243746 241846
rect 244181 241843 244247 241846
rect 197169 241634 197235 241637
rect 245653 241634 245719 241637
rect 197169 241632 200284 241634
rect 197169 241576 197174 241632
rect 197230 241576 200284 241632
rect 197169 241574 200284 241576
rect 244076 241632 245719 241634
rect 244076 241576 245658 241632
rect 245714 241576 245719 241632
rect 244076 241574 245719 241576
rect 197169 241571 197235 241574
rect 245653 241571 245719 241574
rect -960 241090 480 241180
rect 3049 241090 3115 241093
rect -960 241088 3115 241090
rect -960 241032 3054 241088
rect 3110 241032 3115 241088
rect -960 241030 3115 241032
rect -960 240940 480 241030
rect 3049 241027 3115 241030
rect 200113 240138 200179 240141
rect 200254 240138 200314 240788
rect 243862 240549 243922 240788
rect 243862 240544 243971 240549
rect 243862 240488 243910 240544
rect 243966 240488 243971 240544
rect 243862 240486 243971 240488
rect 243905 240483 243971 240486
rect 246021 240274 246087 240277
rect 244076 240272 246087 240274
rect 244076 240216 246026 240272
rect 246082 240216 246087 240272
rect 244076 240214 246087 240216
rect 246021 240211 246087 240214
rect 200113 240136 200314 240138
rect 200113 240080 200118 240136
rect 200174 240080 200314 240136
rect 200113 240078 200314 240080
rect 200113 240075 200179 240078
rect 243905 240002 243971 240005
rect 245285 240002 245351 240005
rect 243905 240000 245351 240002
rect 243905 239944 243910 240000
rect 243966 239944 245290 240000
rect 245346 239944 245351 240000
rect 243905 239942 245351 239944
rect 243905 239939 243971 239942
rect 245285 239939 245351 239942
rect 207933 237962 207999 237965
rect 278998 237962 279004 237964
rect 207933 237960 279004 237962
rect 207933 237904 207938 237960
rect 207994 237904 279004 237960
rect 207933 237902 279004 237904
rect 207933 237899 207999 237902
rect 278998 237900 279004 237902
rect 279068 237900 279074 237964
rect 197905 233882 197971 233885
rect 284702 233882 284708 233884
rect 197905 233880 284708 233882
rect 197905 233824 197910 233880
rect 197966 233824 284708 233880
rect 197905 233822 284708 233824
rect 197905 233819 197971 233822
rect 284702 233820 284708 233822
rect 284772 233820 284778 233884
rect 198273 232658 198339 232661
rect 284518 232658 284524 232660
rect 198273 232656 284524 232658
rect 198273 232600 198278 232656
rect 198334 232600 284524 232656
rect 198273 232598 284524 232600
rect 198273 232595 198339 232598
rect 284518 232596 284524 232598
rect 284588 232596 284594 232660
rect 198089 232522 198155 232525
rect 284886 232522 284892 232524
rect 198089 232520 284892 232522
rect 198089 232464 198094 232520
rect 198150 232464 284892 232520
rect 198089 232462 284892 232464
rect 198089 232459 198155 232462
rect 284886 232460 284892 232462
rect 284956 232460 284962 232524
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect 199510 231100 199516 231164
rect 199580 231162 199586 231164
rect 281574 231162 281580 231164
rect 199580 231102 281580 231162
rect 199580 231100 199586 231102
rect 281574 231100 281580 231102
rect 281644 231100 281650 231164
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 198549 186962 198615 186965
rect 281758 186962 281764 186964
rect 198549 186960 281764 186962
rect 198549 186904 198554 186960
rect 198610 186904 281764 186960
rect 198549 186902 281764 186904
rect 198549 186899 198615 186902
rect 281758 186900 281764 186902
rect 281828 186900 281834 186964
rect 199745 183018 199811 183021
rect 230422 183018 230428 183020
rect 199745 183016 230428 183018
rect 199745 182960 199750 183016
rect 199806 182960 230428 183016
rect 199745 182958 230428 182960
rect 199745 182955 199811 182958
rect 230422 182956 230428 182958
rect 230492 182956 230498 183020
rect 198457 182882 198523 182885
rect 282126 182882 282132 182884
rect 198457 182880 282132 182882
rect 198457 182824 198462 182880
rect 198518 182824 282132 182880
rect 198457 182822 282132 182824
rect 198457 182819 198523 182822
rect 282126 182820 282132 182822
rect 282196 182820 282202 182884
rect 200982 181460 200988 181524
rect 201052 181522 201058 181524
rect 281901 181522 281967 181525
rect 201052 181520 281967 181522
rect 201052 181464 281906 181520
rect 281962 181464 281967 181520
rect 201052 181462 281967 181464
rect 201052 181460 201058 181462
rect 281901 181459 281967 181462
rect 198641 181386 198707 181389
rect 281942 181386 281948 181388
rect 198641 181384 281948 181386
rect 198641 181328 198646 181384
rect 198702 181328 281948 181384
rect 198641 181326 281948 181328
rect 198641 181323 198707 181326
rect 281942 181324 281948 181326
rect 282012 181324 282018 181388
rect 225781 180570 225847 180573
rect 288893 180570 288959 180573
rect 225781 180568 288959 180570
rect 225781 180512 225786 180568
rect 225842 180512 288898 180568
rect 288954 180512 288959 180568
rect 225781 180510 288959 180512
rect 225781 180507 225847 180510
rect 288893 180507 288959 180510
rect 210693 180434 210759 180437
rect 280245 180434 280311 180437
rect 210693 180432 280311 180434
rect 210693 180376 210698 180432
rect 210754 180376 280250 180432
rect 280306 180376 280311 180432
rect 210693 180374 280311 180376
rect 210693 180371 210759 180374
rect 280245 180371 280311 180374
rect 200113 180298 200179 180301
rect 287605 180298 287671 180301
rect 200113 180296 287671 180298
rect 200113 180240 200118 180296
rect 200174 180240 287610 180296
rect 287666 180240 287671 180296
rect 200113 180238 287671 180240
rect 200113 180235 200179 180238
rect 287605 180235 287671 180238
rect 194225 180162 194291 180165
rect 285806 180162 285812 180164
rect 194225 180160 285812 180162
rect 194225 180104 194230 180160
rect 194286 180104 285812 180160
rect 194225 180102 285812 180104
rect 194225 180099 194291 180102
rect 285806 180100 285812 180102
rect 285876 180100 285882 180164
rect 192845 180026 192911 180029
rect 289077 180026 289143 180029
rect 192845 180024 289143 180026
rect 192845 179968 192850 180024
rect 192906 179968 289082 180024
rect 289138 179968 289143 180024
rect 192845 179966 289143 179968
rect 192845 179963 192911 179966
rect 289077 179963 289143 179966
rect 579981 179210 580047 179213
rect 583520 179210 584960 179300
rect 579981 179208 584960 179210
rect 579981 179152 579986 179208
rect 580042 179152 584960 179208
rect 579981 179150 584960 179152
rect 579981 179147 580047 179150
rect 583520 179060 584960 179150
rect 200614 177652 200620 177716
rect 200684 177714 200690 177716
rect 231393 177714 231459 177717
rect 200684 177712 231459 177714
rect 200684 177656 231398 177712
rect 231454 177656 231459 177712
rect 200684 177654 231459 177656
rect 200684 177652 200690 177654
rect 231393 177651 231459 177654
rect 195145 177578 195211 177581
rect 233182 177578 233188 177580
rect 195145 177576 233188 177578
rect 195145 177520 195150 177576
rect 195206 177520 233188 177576
rect 195145 177518 233188 177520
rect 195145 177515 195211 177518
rect 233182 177516 233188 177518
rect 233252 177516 233258 177580
rect 246389 177578 246455 177581
rect 279734 177578 279740 177580
rect 246389 177576 279740 177578
rect 246389 177520 246394 177576
rect 246450 177520 279740 177576
rect 246389 177518 279740 177520
rect 246389 177515 246455 177518
rect 279734 177516 279740 177518
rect 279804 177516 279810 177580
rect 200798 177380 200804 177444
rect 200868 177442 200874 177444
rect 282269 177442 282335 177445
rect 200868 177440 282335 177442
rect 200868 177384 282274 177440
rect 282330 177384 282335 177440
rect 200868 177382 282335 177384
rect 200868 177380 200874 177382
rect 282269 177379 282335 177382
rect 198365 177306 198431 177309
rect 280286 177306 280292 177308
rect 198365 177304 280292 177306
rect 198365 177248 198370 177304
rect 198426 177248 280292 177304
rect 198365 177246 280292 177248
rect 198365 177243 198431 177246
rect 280286 177244 280292 177246
rect 280356 177244 280362 177308
rect 97022 176700 97028 176764
rect 97092 176762 97098 176764
rect 97809 176762 97875 176765
rect 103329 176762 103395 176765
rect 107009 176764 107075 176765
rect 108113 176764 108179 176765
rect 106958 176762 106964 176764
rect 97092 176760 97875 176762
rect 97092 176704 97814 176760
rect 97870 176704 97875 176760
rect 97092 176702 97875 176704
rect 97092 176700 97098 176702
rect 97809 176699 97875 176702
rect 103286 176760 103395 176762
rect 103286 176704 103334 176760
rect 103390 176704 103395 176760
rect 103286 176699 103395 176704
rect 106918 176702 106964 176762
rect 107028 176760 107075 176764
rect 108062 176762 108068 176764
rect 107070 176704 107075 176760
rect 106958 176700 106964 176702
rect 107028 176700 107075 176704
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 108174 176704 108179 176760
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 109534 176700 109540 176764
rect 109604 176762 109610 176764
rect 110045 176762 110111 176765
rect 110689 176764 110755 176765
rect 110638 176762 110644 176764
rect 109604 176760 110111 176762
rect 109604 176704 110050 176760
rect 110106 176704 110111 176760
rect 109604 176702 110111 176704
rect 110598 176702 110644 176762
rect 110708 176760 110755 176764
rect 110750 176704 110755 176760
rect 109604 176700 109610 176702
rect 107009 176699 107075 176700
rect 108113 176699 108179 176700
rect 110045 176699 110111 176702
rect 110638 176700 110644 176702
rect 110708 176700 110755 176704
rect 112110 176700 112116 176764
rect 112180 176762 112186 176764
rect 112621 176762 112687 176765
rect 112180 176760 112687 176762
rect 112180 176704 112626 176760
rect 112682 176704 112687 176760
rect 112180 176702 112687 176704
rect 112180 176700 112186 176702
rect 110689 176699 110755 176700
rect 112621 176699 112687 176702
rect 113214 176700 113220 176764
rect 113284 176762 113290 176764
rect 114001 176762 114067 176765
rect 114369 176764 114435 176765
rect 115841 176764 115907 176765
rect 116945 176764 117011 176765
rect 118417 176764 118483 176765
rect 120809 176764 120875 176765
rect 114318 176762 114324 176764
rect 113284 176760 114067 176762
rect 113284 176704 114006 176760
rect 114062 176704 114067 176760
rect 113284 176702 114067 176704
rect 114278 176702 114324 176762
rect 114388 176760 114435 176764
rect 115790 176762 115796 176764
rect 114430 176704 114435 176760
rect 113284 176700 113290 176702
rect 114001 176699 114067 176702
rect 114318 176700 114324 176702
rect 114388 176700 114435 176704
rect 115750 176702 115796 176762
rect 115860 176760 115907 176764
rect 116894 176762 116900 176764
rect 115902 176704 115907 176760
rect 115790 176700 115796 176702
rect 115860 176700 115907 176704
rect 116854 176702 116900 176762
rect 116964 176760 117011 176764
rect 118366 176762 118372 176764
rect 117006 176704 117011 176760
rect 116894 176700 116900 176702
rect 116964 176700 117011 176704
rect 118326 176702 118372 176762
rect 118436 176760 118483 176764
rect 120758 176762 120764 176764
rect 118478 176704 118483 176760
rect 118366 176700 118372 176702
rect 118436 176700 118483 176704
rect 120718 176702 120764 176762
rect 120828 176760 120875 176764
rect 120870 176704 120875 176760
rect 120758 176700 120764 176702
rect 120828 176700 120875 176704
rect 121862 176700 121868 176764
rect 121932 176762 121938 176764
rect 122281 176762 122347 176765
rect 124489 176764 124555 176765
rect 124438 176762 124444 176764
rect 121932 176760 122347 176762
rect 121932 176704 122286 176760
rect 122342 176704 122347 176760
rect 121932 176702 122347 176704
rect 124398 176702 124444 176762
rect 124508 176760 124555 176764
rect 124550 176704 124555 176760
rect 121932 176700 121938 176702
rect 114369 176699 114435 176700
rect 115841 176699 115907 176700
rect 116945 176699 117011 176700
rect 118417 176699 118483 176700
rect 120809 176699 120875 176700
rect 122281 176699 122347 176702
rect 124438 176700 124444 176702
rect 124508 176700 124555 176704
rect 127014 176700 127020 176764
rect 127084 176762 127090 176764
rect 127985 176762 128051 176765
rect 129457 176764 129523 176765
rect 129406 176762 129412 176764
rect 127084 176760 128051 176762
rect 127084 176704 127990 176760
rect 128046 176704 128051 176760
rect 127084 176702 128051 176704
rect 129366 176702 129412 176762
rect 129476 176760 129523 176764
rect 129518 176704 129523 176760
rect 127084 176700 127090 176702
rect 124489 176699 124555 176700
rect 127985 176699 128051 176702
rect 129406 176700 129412 176702
rect 129476 176700 129523 176704
rect 130694 176700 130700 176764
rect 130764 176762 130770 176764
rect 130929 176762 130995 176765
rect 133137 176764 133203 176765
rect 133086 176762 133092 176764
rect 130764 176760 130995 176762
rect 130764 176704 130934 176760
rect 130990 176704 130995 176760
rect 130764 176702 130995 176704
rect 133046 176702 133092 176762
rect 133156 176760 133203 176764
rect 133198 176704 133203 176760
rect 130764 176700 130770 176702
rect 129457 176699 129523 176700
rect 130929 176699 130995 176702
rect 133086 176700 133092 176702
rect 133156 176700 133203 176704
rect 134374 176700 134380 176764
rect 134444 176762 134450 176764
rect 134517 176762 134583 176765
rect 148225 176764 148291 176765
rect 148174 176762 148180 176764
rect 134444 176760 134583 176762
rect 134444 176704 134522 176760
rect 134578 176704 134583 176760
rect 134444 176702 134583 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 134444 176700 134450 176702
rect 133137 176699 133203 176700
rect 134517 176699 134583 176702
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 148225 176699 148291 176700
rect 103286 176492 103346 176699
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 213913 176218 213979 176221
rect 227713 176218 227779 176221
rect 213913 176216 217242 176218
rect 213913 176160 213918 176216
rect 213974 176160 217242 176216
rect 213913 176158 217242 176160
rect 213913 176155 213979 176158
rect -960 175796 480 176036
rect 217182 175644 217242 176158
rect 227713 176216 228282 176218
rect 227713 176160 227718 176216
rect 227774 176160 228282 176216
rect 227713 176158 228282 176160
rect 227713 176155 227779 176158
rect 228222 175644 228282 176158
rect 278773 176082 278839 176085
rect 278773 176080 279434 176082
rect 278773 176024 278778 176080
rect 278834 176024 279434 176080
rect 278773 176022 279434 176024
rect 278773 176019 278839 176022
rect 135713 175540 135779 175541
rect 135662 175538 135668 175540
rect 135622 175478 135668 175538
rect 135732 175536 135779 175540
rect 135774 175480 135779 175536
rect 135662 175476 135668 175478
rect 135732 175476 135779 175480
rect 135713 175475 135779 175476
rect 98361 175404 98427 175405
rect 99465 175404 99531 175405
rect 100753 175404 100819 175405
rect 102041 175404 102107 175405
rect 104617 175404 104683 175405
rect 105721 175404 105787 175405
rect 128169 175404 128235 175405
rect 132033 175404 132099 175405
rect 158897 175404 158963 175405
rect 98310 175402 98316 175404
rect 98270 175342 98316 175402
rect 98380 175400 98427 175404
rect 99414 175402 99420 175404
rect 98422 175344 98427 175400
rect 98310 175340 98316 175342
rect 98380 175340 98427 175344
rect 99374 175342 99420 175402
rect 99484 175400 99531 175404
rect 100702 175402 100708 175404
rect 99526 175344 99531 175400
rect 99414 175340 99420 175342
rect 99484 175340 99531 175344
rect 100662 175342 100708 175402
rect 100772 175400 100819 175404
rect 101990 175402 101996 175404
rect 100814 175344 100819 175400
rect 100702 175340 100708 175342
rect 100772 175340 100819 175344
rect 101950 175342 101996 175402
rect 102060 175400 102107 175404
rect 104566 175402 104572 175404
rect 102102 175344 102107 175400
rect 101990 175340 101996 175342
rect 102060 175340 102107 175344
rect 104526 175342 104572 175402
rect 104636 175400 104683 175404
rect 105670 175402 105676 175404
rect 104678 175344 104683 175400
rect 104566 175340 104572 175342
rect 104636 175340 104683 175344
rect 105630 175342 105676 175402
rect 105740 175400 105787 175404
rect 128118 175402 128124 175404
rect 105782 175344 105787 175400
rect 105670 175340 105676 175342
rect 105740 175340 105787 175344
rect 128078 175342 128124 175402
rect 128188 175400 128235 175404
rect 131982 175402 131988 175404
rect 128230 175344 128235 175400
rect 128118 175340 128124 175342
rect 128188 175340 128235 175344
rect 131942 175342 131988 175402
rect 132052 175400 132099 175404
rect 158846 175402 158852 175404
rect 132094 175344 132099 175400
rect 131982 175340 131988 175342
rect 132052 175340 132099 175344
rect 158806 175342 158852 175402
rect 158916 175400 158963 175404
rect 158958 175344 158963 175400
rect 158846 175340 158852 175342
rect 158916 175340 158963 175344
rect 98361 175339 98427 175340
rect 99465 175339 99531 175340
rect 100753 175339 100819 175340
rect 102041 175339 102107 175340
rect 104617 175339 104683 175340
rect 105721 175339 105787 175340
rect 128169 175339 128235 175340
rect 132033 175339 132099 175340
rect 158897 175339 158963 175340
rect 265893 175402 265959 175405
rect 268150 175402 268210 175644
rect 279374 175508 279434 176022
rect 265893 175400 268210 175402
rect 265893 175344 265898 175400
rect 265954 175344 268210 175400
rect 265893 175342 268210 175344
rect 265893 175339 265959 175342
rect 231761 175266 231827 175269
rect 228968 175264 231827 175266
rect 228968 175208 231766 175264
rect 231822 175208 231827 175264
rect 228968 175206 231827 175208
rect 231761 175203 231827 175206
rect 213913 175130 213979 175133
rect 213913 175128 217242 175130
rect 213913 175072 213918 175128
rect 213974 175072 217242 175128
rect 213913 175070 217242 175072
rect 213913 175067 213979 175070
rect 119429 174996 119495 174997
rect 123109 174996 123175 174997
rect 125685 174996 125751 174997
rect 119392 174994 119398 174996
rect 119338 174934 119398 174994
rect 119462 174992 119495 174996
rect 123064 174994 123070 174996
rect 119490 174936 119495 174992
rect 119392 174932 119398 174934
rect 119462 174932 119495 174936
rect 123018 174934 123070 174994
rect 123134 174992 123175 174996
rect 125648 174994 125654 174996
rect 123170 174936 123175 174992
rect 123064 174932 123070 174934
rect 123134 174932 123175 174936
rect 125594 174934 125654 174994
rect 125718 174992 125751 174996
rect 125746 174936 125751 174992
rect 217182 174964 217242 175070
rect 266077 174994 266143 174997
rect 268150 174994 268210 175236
rect 279734 175204 279740 175268
rect 279804 175204 279810 175268
rect 266077 174992 268210 174994
rect 125648 174932 125654 174934
rect 125718 174932 125751 174936
rect 119429 174931 119495 174932
rect 123109 174931 123175 174932
rect 125685 174931 125751 174932
rect 266077 174936 266082 174992
rect 266138 174936 268210 174992
rect 266077 174934 268210 174936
rect 266077 174931 266143 174934
rect 214005 174722 214071 174725
rect 230749 174722 230815 174725
rect 214005 174720 217242 174722
rect 214005 174664 214010 174720
rect 214066 174664 217242 174720
rect 214005 174662 217242 174664
rect 228968 174720 230815 174722
rect 228968 174664 230754 174720
rect 230810 174664 230815 174720
rect 228968 174662 230815 174664
rect 214005 174659 214071 174662
rect 217182 174284 217242 174662
rect 230749 174659 230815 174662
rect 265985 174586 266051 174589
rect 268150 174586 268210 174828
rect 279742 174692 279802 175204
rect 265985 174584 268210 174586
rect 265985 174528 265990 174584
rect 266046 174528 268210 174584
rect 265985 174526 268210 174528
rect 265985 174523 266051 174526
rect 268326 174524 268332 174588
rect 268396 174524 268402 174588
rect 264421 174450 264487 174453
rect 267774 174450 267780 174452
rect 264421 174448 267780 174450
rect 264421 174392 264426 174448
rect 264482 174392 267780 174448
rect 264421 174390 267780 174392
rect 264421 174387 264487 174390
rect 267774 174388 267780 174390
rect 267844 174388 267850 174452
rect 268334 174420 268394 174524
rect 229369 174314 229435 174317
rect 228968 174312 229435 174314
rect 228968 174256 229374 174312
rect 229430 174256 229435 174312
rect 228968 174254 229435 174256
rect 229369 174251 229435 174254
rect 265801 174178 265867 174181
rect 265801 174176 268210 174178
rect 265801 174120 265806 174176
rect 265862 174120 268210 174176
rect 265801 174118 268210 174120
rect 265801 174115 265867 174118
rect 268150 174012 268210 174118
rect 281942 174042 281948 174044
rect 279956 173982 281948 174042
rect 281942 173980 281948 173982
rect 282012 173980 282018 174044
rect 213913 173770 213979 173773
rect 230657 173770 230723 173773
rect 213913 173768 217242 173770
rect 213913 173712 213918 173768
rect 213974 173712 217242 173768
rect 213913 173710 217242 173712
rect 228968 173768 230723 173770
rect 228968 173712 230662 173768
rect 230718 173712 230723 173768
rect 228968 173710 230723 173712
rect 213913 173707 213979 173710
rect 217182 173604 217242 173710
rect 230657 173707 230723 173710
rect 265985 173770 266051 173773
rect 265985 173768 268210 173770
rect 265985 173712 265990 173768
rect 266046 173712 268210 173768
rect 265985 173710 268210 173712
rect 265985 173707 266051 173710
rect 268150 173604 268210 173710
rect 214005 173362 214071 173365
rect 231117 173362 231183 173365
rect 214005 173360 217242 173362
rect 214005 173304 214010 173360
rect 214066 173304 217242 173360
rect 214005 173302 217242 173304
rect 228968 173360 231183 173362
rect 228968 173304 231122 173360
rect 231178 173304 231183 173360
rect 228968 173302 231183 173304
rect 214005 173299 214071 173302
rect 217182 172924 217242 173302
rect 231117 173299 231183 173302
rect 265893 173362 265959 173365
rect 265893 173360 268394 173362
rect 265893 173304 265898 173360
rect 265954 173304 268394 173360
rect 265893 173302 268394 173304
rect 265893 173299 265959 173302
rect 268334 173060 268394 173302
rect 282361 173226 282427 173229
rect 279956 173224 282427 173226
rect 279956 173168 282366 173224
rect 282422 173168 282427 173224
rect 279956 173166 282427 173168
rect 282361 173163 282427 173166
rect 231485 172818 231551 172821
rect 228968 172816 231551 172818
rect 228968 172760 231490 172816
rect 231546 172760 231551 172816
rect 228968 172758 231551 172760
rect 231485 172755 231551 172758
rect 265801 172818 265867 172821
rect 265801 172816 268210 172818
rect 265801 172760 265806 172816
rect 265862 172760 268210 172816
rect 265801 172758 268210 172760
rect 265801 172755 265867 172758
rect 268150 172652 268210 172758
rect 213913 172410 213979 172413
rect 231761 172410 231827 172413
rect 281533 172410 281599 172413
rect 213913 172408 217242 172410
rect 213913 172352 213918 172408
rect 213974 172352 217242 172408
rect 213913 172350 217242 172352
rect 228968 172408 231827 172410
rect 228968 172352 231766 172408
rect 231822 172352 231827 172408
rect 228968 172350 231827 172352
rect 279956 172408 281599 172410
rect 279956 172352 281538 172408
rect 281594 172352 281599 172408
rect 279956 172350 281599 172352
rect 213913 172347 213979 172350
rect 217182 172244 217242 172350
rect 231761 172347 231827 172350
rect 281533 172347 281599 172350
rect 214005 172002 214071 172005
rect 265249 172002 265315 172005
rect 268150 172002 268210 172244
rect 279366 172076 279372 172140
rect 279436 172076 279442 172140
rect 214005 172000 217242 172002
rect 214005 171944 214010 172000
rect 214066 171944 217242 172000
rect 214005 171942 217242 171944
rect 214005 171939 214071 171942
rect 169017 171594 169083 171597
rect 164694 171592 169083 171594
rect 164694 171536 169022 171592
rect 169078 171536 169083 171592
rect 217182 171564 217242 171942
rect 265249 172000 268210 172002
rect 265249 171944 265254 172000
rect 265310 171944 268210 172000
rect 265249 171942 268210 171944
rect 265249 171939 265315 171942
rect 231485 171866 231551 171869
rect 228968 171864 231551 171866
rect 228968 171808 231490 171864
rect 231546 171808 231551 171864
rect 228968 171806 231551 171808
rect 231485 171803 231551 171806
rect 265433 171594 265499 171597
rect 268150 171594 268210 171836
rect 279374 171700 279434 172076
rect 265433 171592 268210 171594
rect 164694 171534 169083 171536
rect 169017 171531 169083 171534
rect 265433 171536 265438 171592
rect 265494 171536 268210 171592
rect 265433 171534 268210 171536
rect 265433 171531 265499 171534
rect 231669 171458 231735 171461
rect 228968 171456 231735 171458
rect 228968 171400 231674 171456
rect 231730 171400 231735 171456
rect 228968 171398 231735 171400
rect 231669 171395 231735 171398
rect 265525 171186 265591 171189
rect 268150 171186 268210 171428
rect 216998 171126 217242 171186
rect 214649 171050 214715 171053
rect 216998 171050 217058 171126
rect 214649 171048 217058 171050
rect 214649 170992 214654 171048
rect 214710 170992 217058 171048
rect 217182 171020 217242 171126
rect 265525 171184 268210 171186
rect 265525 171128 265530 171184
rect 265586 171128 268210 171184
rect 265525 171126 268210 171128
rect 265525 171123 265591 171126
rect 214649 170990 217058 170992
rect 214649 170987 214715 170990
rect 231761 170914 231827 170917
rect 228968 170912 231827 170914
rect 228968 170856 231766 170912
rect 231822 170856 231827 170912
rect 228968 170854 231827 170856
rect 231761 170851 231827 170854
rect 213913 170778 213979 170781
rect 213913 170776 217242 170778
rect 213913 170720 213918 170776
rect 213974 170720 217242 170776
rect 213913 170718 217242 170720
rect 213913 170715 213979 170718
rect 217182 170340 217242 170718
rect 265525 170642 265591 170645
rect 268150 170642 268210 171020
rect 282177 170914 282243 170917
rect 279956 170912 282243 170914
rect 279956 170856 282182 170912
rect 282238 170856 282243 170912
rect 279956 170854 282243 170856
rect 282177 170851 282243 170854
rect 265525 170640 268210 170642
rect 265525 170584 265530 170640
rect 265586 170584 268210 170640
rect 265525 170582 268210 170584
rect 265525 170579 265591 170582
rect 231209 170506 231275 170509
rect 228968 170504 231275 170506
rect 228968 170448 231214 170504
rect 231270 170448 231275 170504
rect 228968 170446 231275 170448
rect 231209 170443 231275 170446
rect 265157 170234 265223 170237
rect 268150 170234 268210 170476
rect 265157 170232 268210 170234
rect 265157 170176 265162 170232
rect 265218 170176 268210 170232
rect 265157 170174 268210 170176
rect 265157 170171 265223 170174
rect 281625 170098 281691 170101
rect 279956 170096 281691 170098
rect 231301 169962 231367 169965
rect 228968 169960 231367 169962
rect 228968 169904 231306 169960
rect 231362 169904 231367 169960
rect 228968 169902 231367 169904
rect 231301 169899 231367 169902
rect 265801 169826 265867 169829
rect 268334 169826 268394 170068
rect 279956 170040 281630 170096
rect 281686 170040 281691 170096
rect 279956 170038 281691 170040
rect 281625 170035 281691 170038
rect 216998 169766 217242 169826
rect 213913 169690 213979 169693
rect 216998 169690 217058 169766
rect 213913 169688 217058 169690
rect 213913 169632 213918 169688
rect 213974 169632 217058 169688
rect 217182 169660 217242 169766
rect 265801 169824 268394 169826
rect 265801 169768 265806 169824
rect 265862 169768 268394 169824
rect 265801 169766 268394 169768
rect 265801 169763 265867 169766
rect 279550 169764 279556 169828
rect 279620 169764 279626 169828
rect 213913 169630 217058 169632
rect 213913 169627 213979 169630
rect 229185 169554 229251 169557
rect 228968 169552 229251 169554
rect 228968 169496 229190 169552
rect 229246 169496 229251 169552
rect 228968 169494 229251 169496
rect 229185 169491 229251 169494
rect 214005 169418 214071 169421
rect 265893 169418 265959 169421
rect 268150 169418 268210 169660
rect 214005 169416 217242 169418
rect 214005 169360 214010 169416
rect 214066 169360 217242 169416
rect 214005 169358 217242 169360
rect 214005 169355 214071 169358
rect 217182 168980 217242 169358
rect 265893 169416 268210 169418
rect 265893 169360 265898 169416
rect 265954 169360 268210 169416
rect 279558 169388 279618 169764
rect 265893 169358 268210 169360
rect 265893 169355 265959 169358
rect 229553 169010 229619 169013
rect 228968 169008 229619 169010
rect 228968 168952 229558 169008
rect 229614 168952 229619 169008
rect 228968 168950 229619 168952
rect 229553 168947 229619 168950
rect 265985 169010 266051 169013
rect 268150 169010 268210 169252
rect 265985 169008 268210 169010
rect 265985 168952 265990 169008
rect 266046 168952 268210 169008
rect 265985 168950 268210 168952
rect 265985 168947 266051 168950
rect 231761 168602 231827 168605
rect 228968 168600 231827 168602
rect 228968 168544 231766 168600
rect 231822 168544 231827 168600
rect 228968 168542 231827 168544
rect 231761 168539 231827 168542
rect 265801 168602 265867 168605
rect 268150 168602 268210 168844
rect 281717 168602 281783 168605
rect 265801 168600 268210 168602
rect 265801 168544 265806 168600
rect 265862 168544 268210 168600
rect 265801 168542 268210 168544
rect 279956 168600 281783 168602
rect 279956 168544 281722 168600
rect 281778 168544 281783 168600
rect 279956 168542 281783 168544
rect 265801 168539 265867 168542
rect 281717 168539 281783 168542
rect 265893 168466 265959 168469
rect 265893 168464 267842 168466
rect 265893 168408 265898 168464
rect 265954 168408 267842 168464
rect 265893 168406 267842 168408
rect 265893 168403 265959 168406
rect 213913 168058 213979 168061
rect 217182 168058 217242 168300
rect 267782 168194 267842 168406
rect 268334 168194 268394 168436
rect 267782 168134 268394 168194
rect 231761 168058 231827 168061
rect 213913 168056 217242 168058
rect 213913 168000 213918 168056
rect 213974 168000 217242 168056
rect 213913 167998 217242 168000
rect 228968 168056 231827 168058
rect 228968 168000 231766 168056
rect 231822 168000 231827 168056
rect 228968 167998 231827 168000
rect 213913 167995 213979 167998
rect 231761 167995 231827 167998
rect 214005 167922 214071 167925
rect 214005 167920 217242 167922
rect 214005 167864 214010 167920
rect 214066 167864 217242 167920
rect 214005 167862 217242 167864
rect 214005 167859 214071 167862
rect 217182 167620 217242 167862
rect 231485 167650 231551 167653
rect 228968 167648 231551 167650
rect 228968 167592 231490 167648
rect 231546 167592 231551 167648
rect 228968 167590 231551 167592
rect 231485 167587 231551 167590
rect 265341 167650 265407 167653
rect 268150 167650 268210 167892
rect 281809 167786 281875 167789
rect 279956 167784 281875 167786
rect 279956 167728 281814 167784
rect 281870 167728 281875 167784
rect 279956 167726 281875 167728
rect 281809 167723 281875 167726
rect 265341 167648 268210 167650
rect 265341 167592 265346 167648
rect 265402 167592 268210 167648
rect 265341 167590 268210 167592
rect 265341 167587 265407 167590
rect 265801 167242 265867 167245
rect 268150 167242 268210 167484
rect 265801 167240 268210 167242
rect 265801 167184 265806 167240
rect 265862 167184 268210 167240
rect 265801 167182 268210 167184
rect 265801 167179 265867 167182
rect 231393 167106 231459 167109
rect 228968 167104 231459 167106
rect 228968 167048 231398 167104
rect 231454 167048 231459 167104
rect 228968 167046 231459 167048
rect 231393 167043 231459 167046
rect 265157 167106 265223 167109
rect 282269 167106 282335 167109
rect 265157 167104 268026 167106
rect 265157 167048 265162 167104
rect 265218 167048 268026 167104
rect 279956 167104 282335 167106
rect 265157 167046 268026 167048
rect 265157 167043 265223 167046
rect 267966 167010 268026 167046
rect 268150 167010 268210 167076
rect 279956 167048 282274 167104
rect 282330 167048 282335 167104
rect 279956 167046 282335 167048
rect 282269 167043 282335 167046
rect 213913 166970 213979 166973
rect 216998 166970 217242 167010
rect 213913 166968 217242 166970
rect 213913 166912 213918 166968
rect 213974 166950 217242 166968
rect 267966 166950 268210 167010
rect 213974 166912 217058 166950
rect 217182 166940 217242 166950
rect 213913 166910 217058 166912
rect 213913 166907 213979 166910
rect 214005 166698 214071 166701
rect 231301 166698 231367 166701
rect 214005 166696 217242 166698
rect 214005 166640 214010 166696
rect 214066 166640 217242 166696
rect 214005 166638 217242 166640
rect 228968 166696 231367 166698
rect 228968 166640 231306 166696
rect 231362 166640 231367 166696
rect 228968 166638 231367 166640
rect 214005 166635 214071 166638
rect 217182 166396 217242 166638
rect 231301 166635 231367 166638
rect 265801 166426 265867 166429
rect 268150 166426 268210 166668
rect 265801 166424 268210 166426
rect 265801 166368 265806 166424
rect 265862 166368 268210 166424
rect 265801 166366 268210 166368
rect 265801 166363 265867 166366
rect 281758 166290 281764 166292
rect 214097 166154 214163 166157
rect 231761 166154 231827 166157
rect 214097 166152 217242 166154
rect 214097 166096 214102 166152
rect 214158 166096 217242 166152
rect 214097 166094 217242 166096
rect 228968 166152 231827 166154
rect 228968 166096 231766 166152
rect 231822 166096 231827 166152
rect 228968 166094 231827 166096
rect 214097 166091 214163 166094
rect 217182 165716 217242 166094
rect 231761 166091 231827 166094
rect 265433 166018 265499 166021
rect 268150 166018 268210 166260
rect 279956 166230 281764 166290
rect 281758 166228 281764 166230
rect 281828 166228 281834 166292
rect 265433 166016 268210 166018
rect 265433 165960 265438 166016
rect 265494 165960 268210 166016
rect 265433 165958 268210 165960
rect 265433 165955 265499 165958
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 231761 165746 231827 165749
rect 228968 165744 231827 165746
rect 228968 165688 231766 165744
rect 231822 165688 231827 165744
rect 228968 165686 231827 165688
rect 231761 165683 231827 165686
rect 264421 165746 264487 165749
rect 264421 165744 267842 165746
rect 264421 165688 264426 165744
rect 264482 165688 267842 165744
rect 264421 165686 267842 165688
rect 264421 165683 264487 165686
rect 267782 165610 267842 165686
rect 268334 165610 268394 165852
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 267782 165550 268394 165610
rect 213913 165474 213979 165477
rect 282821 165474 282887 165477
rect 213913 165472 217242 165474
rect 213913 165416 213918 165472
rect 213974 165416 217242 165472
rect 213913 165414 217242 165416
rect 279956 165472 282887 165474
rect 279956 165416 282826 165472
rect 282882 165416 282887 165472
rect 279956 165414 282887 165416
rect 213913 165411 213979 165414
rect 217182 165036 217242 165414
rect 282821 165411 282887 165414
rect 231761 165202 231827 165205
rect 228968 165200 231827 165202
rect 228968 165144 231766 165200
rect 231822 165144 231827 165200
rect 228968 165142 231827 165144
rect 231761 165139 231827 165142
rect 265433 165066 265499 165069
rect 268150 165066 268210 165308
rect 265433 165064 268210 165066
rect 265433 165008 265438 165064
rect 265494 165008 268210 165064
rect 265433 165006 268210 165008
rect 265433 165003 265499 165006
rect 214005 164794 214071 164797
rect 231393 164794 231459 164797
rect 214005 164792 217242 164794
rect 214005 164736 214010 164792
rect 214066 164736 217242 164792
rect 214005 164734 217242 164736
rect 228968 164792 231459 164794
rect 228968 164736 231398 164792
rect 231454 164736 231459 164792
rect 228968 164734 231459 164736
rect 214005 164731 214071 164734
rect 217182 164356 217242 164734
rect 231393 164731 231459 164734
rect 265893 164658 265959 164661
rect 268150 164658 268210 164900
rect 281993 164794 282059 164797
rect 279956 164792 282059 164794
rect 279956 164736 281998 164792
rect 282054 164736 282059 164792
rect 279956 164734 282059 164736
rect 281993 164731 282059 164734
rect 265893 164656 268210 164658
rect 265893 164600 265898 164656
rect 265954 164600 268210 164656
rect 265893 164598 268210 164600
rect 265893 164595 265959 164598
rect 231761 164386 231827 164389
rect 228968 164384 231827 164386
rect 228968 164328 231766 164384
rect 231822 164328 231827 164384
rect 228968 164326 231827 164328
rect 231761 164323 231827 164326
rect 265801 164250 265867 164253
rect 268334 164250 268394 164492
rect 265801 164248 268394 164250
rect 265801 164192 265806 164248
rect 265862 164192 268394 164248
rect 265801 164190 268394 164192
rect 265801 164187 265867 164190
rect 213913 163978 213979 163981
rect 213913 163976 217242 163978
rect 213913 163920 213918 163976
rect 213974 163920 217242 163976
rect 213913 163918 217242 163920
rect 213913 163915 213979 163918
rect 217182 163676 217242 163918
rect 231393 163842 231459 163845
rect 228968 163840 231459 163842
rect 228968 163784 231398 163840
rect 231454 163784 231459 163840
rect 228968 163782 231459 163784
rect 231393 163779 231459 163782
rect 265157 163842 265223 163845
rect 268150 163842 268210 164084
rect 282126 163978 282132 163980
rect 279956 163918 282132 163978
rect 282126 163916 282132 163918
rect 282196 163916 282202 163980
rect 265157 163840 268210 163842
rect 265157 163784 265162 163840
rect 265218 163784 268210 163840
rect 265157 163782 268210 163784
rect 265157 163779 265223 163782
rect 214005 163434 214071 163437
rect 231761 163434 231827 163437
rect 214005 163432 217242 163434
rect 214005 163376 214010 163432
rect 214066 163376 217242 163432
rect 214005 163374 217242 163376
rect 228968 163432 231827 163434
rect 228968 163376 231766 163432
rect 231822 163376 231827 163432
rect 228968 163374 231827 163376
rect 214005 163371 214071 163374
rect 217182 162996 217242 163374
rect 231761 163371 231827 163374
rect 264697 163434 264763 163437
rect 268150 163434 268210 163676
rect 264697 163432 268210 163434
rect 264697 163376 264702 163432
rect 264758 163376 268210 163432
rect 264697 163374 268210 163376
rect 264697 163371 264763 163374
rect 265801 163026 265867 163029
rect 268518 163028 268578 163268
rect 281574 163162 281580 163164
rect 279956 163102 281580 163162
rect 281574 163100 281580 163102
rect 281644 163100 281650 163164
rect 265801 163024 268210 163026
rect -960 162890 480 162980
rect 265801 162968 265806 163024
rect 265862 162968 268210 163024
rect 265801 162966 268210 162968
rect 265801 162963 265867 162966
rect 3233 162890 3299 162893
rect 231485 162890 231551 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect 228968 162888 231551 162890
rect 228968 162832 231490 162888
rect 231546 162832 231551 162888
rect 268150 162860 268210 162966
rect 268510 162964 268516 163028
rect 268580 162964 268586 163028
rect 228968 162830 231551 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 231485 162827 231551 162830
rect 213913 162618 213979 162621
rect 213913 162616 217242 162618
rect 213913 162560 213918 162616
rect 213974 162560 217242 162616
rect 213913 162558 217242 162560
rect 213913 162555 213979 162558
rect 217182 162316 217242 162558
rect 244038 162482 244044 162484
rect 228968 162422 244044 162482
rect 244038 162420 244044 162422
rect 244108 162420 244114 162484
rect 282085 162482 282151 162485
rect 279956 162480 282151 162482
rect 279956 162424 282090 162480
rect 282146 162424 282151 162480
rect 279956 162422 282151 162424
rect 282085 162419 282151 162422
rect 214005 162074 214071 162077
rect 265433 162074 265499 162077
rect 268150 162074 268210 162316
rect 214005 162072 217242 162074
rect 214005 162016 214010 162072
rect 214066 162016 217242 162072
rect 214005 162014 217242 162016
rect 214005 162011 214071 162014
rect 217182 161772 217242 162014
rect 265433 162072 268210 162074
rect 265433 162016 265438 162072
rect 265494 162016 268210 162072
rect 265433 162014 268210 162016
rect 265433 162011 265499 162014
rect 231025 161938 231091 161941
rect 228968 161936 231091 161938
rect 228968 161880 231030 161936
rect 231086 161880 231091 161936
rect 228968 161878 231091 161880
rect 231025 161875 231091 161878
rect 265801 161666 265867 161669
rect 268150 161666 268210 161908
rect 282821 161666 282887 161669
rect 265801 161664 268210 161666
rect 265801 161608 265806 161664
rect 265862 161608 268210 161664
rect 265801 161606 268210 161608
rect 279956 161664 282887 161666
rect 279956 161608 282826 161664
rect 282882 161608 282887 161664
rect 279956 161606 282887 161608
rect 265801 161603 265867 161606
rect 282821 161603 282887 161606
rect 229461 161530 229527 161533
rect 228968 161528 229527 161530
rect 228968 161472 229466 161528
rect 229522 161472 229527 161528
rect 228968 161470 229527 161472
rect 229461 161467 229527 161470
rect 266261 161530 266327 161533
rect 266261 161528 267842 161530
rect 266261 161472 266266 161528
rect 266322 161472 267842 161528
rect 266261 161470 267842 161472
rect 266261 161467 266327 161470
rect 213913 161394 213979 161397
rect 213913 161392 217242 161394
rect 213913 161336 213918 161392
rect 213974 161336 217242 161392
rect 213913 161334 217242 161336
rect 213913 161331 213979 161334
rect 217182 161092 217242 161334
rect 267782 161258 267842 161470
rect 268334 161258 268394 161500
rect 267782 161198 268394 161258
rect 231761 160986 231827 160989
rect 228968 160984 231827 160986
rect 228968 160928 231766 160984
rect 231822 160928 231827 160984
rect 228968 160926 231827 160928
rect 231761 160923 231827 160926
rect 214741 160850 214807 160853
rect 265985 160850 266051 160853
rect 268150 160850 268210 161092
rect 282177 160850 282243 160853
rect 214741 160848 217242 160850
rect 214741 160792 214746 160848
rect 214802 160792 217242 160848
rect 214741 160790 217242 160792
rect 214741 160787 214807 160790
rect 217182 160412 217242 160790
rect 265985 160848 268210 160850
rect 265985 160792 265990 160848
rect 266046 160792 268210 160848
rect 265985 160790 268210 160792
rect 279956 160848 282243 160850
rect 279956 160792 282182 160848
rect 282238 160792 282243 160848
rect 279956 160790 282243 160792
rect 265985 160787 266051 160790
rect 282177 160787 282243 160790
rect 231761 160578 231827 160581
rect 228968 160576 231827 160578
rect 228968 160520 231766 160576
rect 231822 160520 231827 160576
rect 228968 160518 231827 160520
rect 231761 160515 231827 160518
rect 265893 160442 265959 160445
rect 268150 160442 268210 160684
rect 265893 160440 268210 160442
rect 265893 160384 265898 160440
rect 265954 160384 268210 160440
rect 265893 160382 268210 160384
rect 265893 160379 265959 160382
rect 265525 160170 265591 160173
rect 265525 160168 267842 160170
rect 265525 160112 265530 160168
rect 265586 160112 267842 160168
rect 265525 160110 267842 160112
rect 265525 160107 265591 160110
rect 231761 160034 231827 160037
rect 228968 160032 231827 160034
rect 228968 159976 231766 160032
rect 231822 159976 231827 160032
rect 228968 159974 231827 159976
rect 267782 160034 267842 160110
rect 268334 160034 268394 160276
rect 280705 160170 280771 160173
rect 279956 160168 280771 160170
rect 279956 160112 280710 160168
rect 280766 160112 280771 160168
rect 279956 160110 280771 160112
rect 280705 160107 280771 160110
rect 267782 159974 268394 160034
rect 231761 159971 231827 159974
rect 213913 159898 213979 159901
rect 262949 159898 263015 159901
rect 268510 159898 268516 159900
rect 213913 159896 217242 159898
rect 213913 159840 213918 159896
rect 213974 159840 217242 159896
rect 213913 159838 217242 159840
rect 213913 159835 213979 159838
rect 217182 159732 217242 159838
rect 262949 159896 268516 159898
rect 262949 159840 262954 159896
rect 263010 159840 268516 159896
rect 262949 159838 268516 159840
rect 262949 159835 263015 159838
rect 268510 159836 268516 159838
rect 268580 159836 268586 159900
rect 230657 159626 230723 159629
rect 228968 159624 230723 159626
rect 228968 159568 230662 159624
rect 230718 159568 230723 159624
rect 228968 159566 230723 159568
rect 230657 159563 230723 159566
rect 214005 159490 214071 159493
rect 265893 159490 265959 159493
rect 268150 159490 268210 159732
rect 214005 159488 217242 159490
rect 214005 159432 214010 159488
rect 214066 159432 217242 159488
rect 214005 159430 217242 159432
rect 214005 159427 214071 159430
rect 217182 159052 217242 159430
rect 265893 159488 268210 159490
rect 265893 159432 265898 159488
rect 265954 159432 268210 159488
rect 265893 159430 268210 159432
rect 265893 159427 265959 159430
rect 282821 159354 282887 159357
rect 279956 159352 282887 159354
rect 231209 159082 231275 159085
rect 228968 159080 231275 159082
rect 228968 159024 231214 159080
rect 231270 159024 231275 159080
rect 228968 159022 231275 159024
rect 231209 159019 231275 159022
rect 265433 159082 265499 159085
rect 268150 159082 268210 159324
rect 279956 159296 282826 159352
rect 282882 159296 282887 159352
rect 279956 159294 282887 159296
rect 282821 159291 282887 159294
rect 265433 159080 268210 159082
rect 265433 159024 265438 159080
rect 265494 159024 268210 159080
rect 265433 159022 268210 159024
rect 265433 159019 265499 159022
rect 265341 158810 265407 158813
rect 265341 158808 267842 158810
rect 265341 158752 265346 158808
rect 265402 158752 267842 158808
rect 265341 158750 267842 158752
rect 265341 158747 265407 158750
rect 214465 158674 214531 158677
rect 230473 158674 230539 158677
rect 214465 158672 217242 158674
rect 214465 158616 214470 158672
rect 214526 158616 217242 158672
rect 214465 158614 217242 158616
rect 228968 158672 230539 158674
rect 228968 158616 230478 158672
rect 230534 158616 230539 158672
rect 228968 158614 230539 158616
rect 267782 158674 267842 158750
rect 268334 158674 268394 158916
rect 267782 158614 268394 158674
rect 214465 158611 214531 158614
rect 217182 158372 217242 158614
rect 230473 158611 230539 158614
rect 281901 158538 281967 158541
rect 279956 158536 281967 158538
rect 265893 158266 265959 158269
rect 268150 158266 268210 158508
rect 279956 158480 281906 158536
rect 281962 158480 281967 158536
rect 279956 158478 281967 158480
rect 281901 158475 281967 158478
rect 265893 158264 268210 158266
rect 265893 158208 265898 158264
rect 265954 158208 268210 158264
rect 265893 158206 268210 158208
rect 265893 158203 265959 158206
rect 213913 158130 213979 158133
rect 231761 158130 231827 158133
rect 213913 158128 217242 158130
rect 213913 158072 213918 158128
rect 213974 158072 217242 158128
rect 213913 158070 217242 158072
rect 228968 158128 231827 158130
rect 228968 158072 231766 158128
rect 231822 158072 231827 158128
rect 228968 158070 231827 158072
rect 213913 158067 213979 158070
rect 217182 157692 217242 158070
rect 231761 158067 231827 158070
rect 265157 157858 265223 157861
rect 268150 157858 268210 158100
rect 281993 157858 282059 157861
rect 265157 157856 268210 157858
rect 265157 157800 265162 157856
rect 265218 157800 268210 157856
rect 265157 157798 268210 157800
rect 279956 157856 282059 157858
rect 279956 157800 281998 157856
rect 282054 157800 282059 157856
rect 279956 157798 282059 157800
rect 265157 157795 265223 157798
rect 281993 157795 282059 157798
rect 231025 157722 231091 157725
rect 228968 157720 231091 157722
rect 228968 157664 231030 157720
rect 231086 157664 231091 157720
rect 228968 157662 231091 157664
rect 231025 157659 231091 157662
rect 265801 157450 265867 157453
rect 268150 157450 268210 157692
rect 265801 157448 268210 157450
rect 265801 157392 265806 157448
rect 265862 157392 268210 157448
rect 265801 157390 268210 157392
rect 265801 157387 265867 157390
rect 213913 157314 213979 157317
rect 213913 157312 217242 157314
rect 213913 157256 213918 157312
rect 213974 157256 217242 157312
rect 213913 157254 217242 157256
rect 213913 157251 213979 157254
rect 217182 157148 217242 157254
rect 231761 157178 231827 157181
rect 228968 157176 231827 157178
rect 228968 157120 231766 157176
rect 231822 157120 231827 157176
rect 228968 157118 231827 157120
rect 231761 157115 231827 157118
rect 214005 156906 214071 156909
rect 265893 156906 265959 156909
rect 268150 156906 268210 157148
rect 282821 157042 282887 157045
rect 279956 157040 282887 157042
rect 279956 156984 282826 157040
rect 282882 156984 282887 157040
rect 279956 156982 282887 156984
rect 282821 156979 282887 156982
rect 214005 156904 217242 156906
rect 214005 156848 214010 156904
rect 214066 156848 217242 156904
rect 214005 156846 217242 156848
rect 214005 156843 214071 156846
rect 217182 156468 217242 156846
rect 265893 156904 268210 156906
rect 265893 156848 265898 156904
rect 265954 156848 268210 156904
rect 265893 156846 268210 156848
rect 265893 156843 265959 156846
rect 231485 156770 231551 156773
rect 228968 156768 231551 156770
rect 228968 156712 231490 156768
rect 231546 156712 231551 156768
rect 228968 156710 231551 156712
rect 231485 156707 231551 156710
rect 265801 156498 265867 156501
rect 268150 156498 268210 156740
rect 265801 156496 268210 156498
rect 265801 156440 265806 156496
rect 265862 156440 268210 156496
rect 265801 156438 268210 156440
rect 265801 156435 265867 156438
rect 282453 156362 282519 156365
rect 279956 156360 282519 156362
rect 231117 156226 231183 156229
rect 228968 156224 231183 156226
rect 228968 156168 231122 156224
rect 231178 156168 231183 156224
rect 228968 156166 231183 156168
rect 231117 156163 231183 156166
rect 266077 156090 266143 156093
rect 268150 156090 268210 156332
rect 279956 156304 282458 156360
rect 282514 156304 282519 156360
rect 279956 156302 282519 156304
rect 282453 156299 282519 156302
rect 266077 156088 268210 156090
rect 266077 156032 266082 156088
rect 266138 156032 268210 156088
rect 266077 156030 268210 156032
rect 266077 156027 266143 156030
rect 213913 155954 213979 155957
rect 213913 155952 217242 155954
rect 213913 155896 213918 155952
rect 213974 155896 217242 155952
rect 213913 155894 217242 155896
rect 213913 155891 213979 155894
rect 217182 155788 217242 155894
rect 230473 155818 230539 155821
rect 228968 155816 230539 155818
rect 228968 155760 230478 155816
rect 230534 155760 230539 155816
rect 228968 155758 230539 155760
rect 230473 155755 230539 155758
rect 265433 155682 265499 155685
rect 268150 155682 268210 155924
rect 265433 155680 268210 155682
rect 265433 155624 265438 155680
rect 265494 155624 268210 155680
rect 265433 155622 268210 155624
rect 265433 155619 265499 155622
rect 282821 155546 282887 155549
rect 279956 155544 282887 155546
rect 214005 155410 214071 155413
rect 214005 155408 217242 155410
rect 214005 155352 214010 155408
rect 214066 155352 217242 155408
rect 214005 155350 217242 155352
rect 214005 155347 214071 155350
rect 217182 155108 217242 155350
rect 230473 155274 230539 155277
rect 228968 155272 230539 155274
rect 228968 155216 230478 155272
rect 230534 155216 230539 155272
rect 228968 155214 230539 155216
rect 230473 155211 230539 155214
rect 265525 155274 265591 155277
rect 268150 155274 268210 155516
rect 279956 155488 282826 155544
rect 282882 155488 282887 155544
rect 279956 155486 282887 155488
rect 282821 155483 282887 155486
rect 265525 155272 268210 155274
rect 265525 155216 265530 155272
rect 265586 155216 268210 155272
rect 265525 155214 268210 155216
rect 265525 155211 265591 155214
rect 230565 154866 230631 154869
rect 228968 154864 230631 154866
rect 228968 154808 230570 154864
rect 230626 154808 230631 154864
rect 228968 154806 230631 154808
rect 230565 154803 230631 154806
rect 265801 154866 265867 154869
rect 268150 154866 268210 155108
rect 265801 154864 268210 154866
rect 265801 154808 265806 154864
rect 265862 154808 268210 154864
rect 265801 154806 268210 154808
rect 265801 154803 265867 154806
rect 265985 154730 266051 154733
rect 281809 154730 281875 154733
rect 265985 154728 268210 154730
rect 265985 154672 265990 154728
rect 266046 154672 268210 154728
rect 265985 154670 268210 154672
rect 279956 154728 281875 154730
rect 279956 154672 281814 154728
rect 281870 154672 281875 154728
rect 279956 154670 281875 154672
rect 265985 154667 266051 154670
rect 268150 154564 268210 154670
rect 281809 154667 281875 154670
rect 214005 153914 214071 153917
rect 217182 153914 217242 154428
rect 229277 154322 229343 154325
rect 228968 154320 229343 154322
rect 228968 154264 229282 154320
rect 229338 154264 229343 154320
rect 228968 154262 229343 154264
rect 229277 154259 229343 154262
rect 230841 153914 230907 153917
rect 214005 153912 217242 153914
rect 214005 153856 214010 153912
rect 214066 153856 217242 153912
rect 214005 153854 217242 153856
rect 228968 153912 230907 153914
rect 228968 153856 230846 153912
rect 230902 153856 230907 153912
rect 228968 153854 230907 153856
rect 214005 153851 214071 153854
rect 230841 153851 230907 153854
rect 265525 153914 265591 153917
rect 268150 153914 268210 154156
rect 282085 154050 282151 154053
rect 279956 154048 282151 154050
rect 279956 153992 282090 154048
rect 282146 153992 282151 154048
rect 279956 153990 282151 153992
rect 282085 153987 282151 153990
rect 265525 153912 268210 153914
rect 265525 153856 265530 153912
rect 265586 153856 268210 153912
rect 265525 153854 268210 153856
rect 265525 153851 265591 153854
rect 213913 153506 213979 153509
rect 217182 153506 217242 153748
rect 213913 153504 217242 153506
rect 213913 153448 213918 153504
rect 213974 153448 217242 153504
rect 213913 153446 217242 153448
rect 265801 153506 265867 153509
rect 268518 153508 268578 153748
rect 265801 153504 268210 153506
rect 265801 153448 265806 153504
rect 265862 153448 268210 153504
rect 265801 153446 268210 153448
rect 213913 153443 213979 153446
rect 265801 153443 265867 153446
rect 229369 153370 229435 153373
rect 228968 153368 229435 153370
rect 228968 153312 229374 153368
rect 229430 153312 229435 153368
rect 268150 153340 268210 153446
rect 268510 153444 268516 153508
rect 268580 153444 268586 153508
rect 228968 153310 229435 153312
rect 229369 153307 229435 153310
rect 282269 153234 282335 153237
rect 279956 153232 282335 153234
rect 279956 153176 282274 153232
rect 282330 153176 282335 153232
rect 279956 153174 282335 153176
rect 282269 153171 282335 153174
rect 264513 153098 264579 153101
rect 268510 153098 268516 153100
rect 264513 153096 268516 153098
rect 213913 152690 213979 152693
rect 217182 152690 217242 153068
rect 264513 153040 264518 153096
rect 264574 153040 268516 153096
rect 264513 153038 268516 153040
rect 264513 153035 264579 153038
rect 268510 153036 268516 153038
rect 268580 153036 268586 153100
rect 231761 152962 231827 152965
rect 228968 152960 231827 152962
rect 228968 152904 231766 152960
rect 231822 152904 231827 152960
rect 228968 152902 231827 152904
rect 231761 152899 231827 152902
rect 213913 152688 217242 152690
rect 213913 152632 213918 152688
rect 213974 152632 217242 152688
rect 213913 152630 217242 152632
rect 265249 152690 265315 152693
rect 268150 152690 268210 152932
rect 583520 152690 584960 152780
rect 265249 152688 268210 152690
rect 265249 152632 265254 152688
rect 265310 152632 268210 152688
rect 265249 152630 268210 152632
rect 583342 152630 584960 152690
rect 213913 152627 213979 152630
rect 265249 152627 265315 152630
rect 231117 152554 231183 152557
rect 228968 152552 231183 152554
rect 214741 152146 214807 152149
rect 217182 152146 217242 152524
rect 228968 152496 231122 152552
rect 231178 152496 231183 152552
rect 583342 152554 583402 152630
rect 583520 152554 584960 152630
rect 583342 152540 584960 152554
rect 228968 152494 231183 152496
rect 231117 152491 231183 152494
rect 214741 152144 217242 152146
rect 214741 152088 214746 152144
rect 214802 152088 217242 152144
rect 214741 152086 217242 152088
rect 265893 152146 265959 152149
rect 268150 152146 268210 152524
rect 583342 152494 583586 152540
rect 282085 152418 282151 152421
rect 279956 152416 282151 152418
rect 279956 152360 282090 152416
rect 282146 152360 282151 152416
rect 279956 152358 282151 152360
rect 282085 152355 282151 152358
rect 265893 152144 268210 152146
rect 265893 152088 265898 152144
rect 265954 152088 268210 152144
rect 265893 152086 268210 152088
rect 214741 152083 214807 152086
rect 265893 152083 265959 152086
rect 214833 152010 214899 152013
rect 231301 152010 231367 152013
rect 214833 152008 217242 152010
rect 214833 151952 214838 152008
rect 214894 151952 217242 152008
rect 214833 151950 217242 151952
rect 228968 152008 231367 152010
rect 228968 151952 231306 152008
rect 231362 151952 231367 152008
rect 228968 151950 231367 151952
rect 214833 151947 214899 151950
rect 217182 151844 217242 151950
rect 231301 151947 231367 151950
rect 265801 151874 265867 151877
rect 265801 151872 267842 151874
rect 265801 151816 265806 151872
rect 265862 151816 267842 151872
rect 265801 151814 267842 151816
rect 265801 151811 265867 151814
rect 267782 151738 267842 151814
rect 268334 151738 268394 151980
rect 288934 151812 288940 151876
rect 289004 151874 289010 151876
rect 583526 151874 583586 152494
rect 289004 151814 583586 151874
rect 289004 151812 289010 151814
rect 282269 151738 282335 151741
rect 267782 151678 268394 151738
rect 279956 151736 282335 151738
rect 279956 151680 282274 151736
rect 282330 151680 282335 151736
rect 279956 151678 282335 151680
rect 282269 151675 282335 151678
rect 231577 151602 231643 151605
rect 228968 151600 231643 151602
rect 228968 151544 231582 151600
rect 231638 151544 231643 151600
rect 228968 151542 231643 151544
rect 231577 151539 231643 151542
rect 265801 151330 265867 151333
rect 268150 151330 268210 151572
rect 265801 151328 268210 151330
rect 265801 151272 265806 151328
rect 265862 151272 268210 151328
rect 265801 151270 268210 151272
rect 265801 151267 265867 151270
rect 214005 150922 214071 150925
rect 217182 150922 217242 151164
rect 230749 151058 230815 151061
rect 228968 151056 230815 151058
rect 228968 151000 230754 151056
rect 230810 151000 230815 151056
rect 228968 150998 230815 151000
rect 230749 150995 230815 150998
rect 214005 150920 217242 150922
rect 214005 150864 214010 150920
rect 214066 150864 217242 150920
rect 214005 150862 217242 150864
rect 265341 150922 265407 150925
rect 268150 150922 268210 151164
rect 281625 150922 281691 150925
rect 265341 150920 268210 150922
rect 265341 150864 265346 150920
rect 265402 150864 268210 150920
rect 265341 150862 268210 150864
rect 279956 150920 281691 150922
rect 279956 150864 281630 150920
rect 281686 150864 281691 150920
rect 279956 150862 281691 150864
rect 214005 150859 214071 150862
rect 265341 150859 265407 150862
rect 281625 150859 281691 150862
rect 214741 150786 214807 150789
rect 214741 150784 217426 150786
rect 214741 150728 214746 150784
rect 214802 150728 217426 150784
rect 214741 150726 217426 150728
rect 214741 150723 214807 150726
rect 217366 150484 217426 150726
rect 229093 150650 229159 150653
rect 228968 150648 229159 150650
rect 228968 150592 229098 150648
rect 229154 150592 229159 150648
rect 228968 150590 229159 150592
rect 229093 150587 229159 150590
rect 265065 150514 265131 150517
rect 268150 150514 268210 150756
rect 265065 150512 268210 150514
rect 265065 150456 265070 150512
rect 265126 150456 268210 150512
rect 265065 150454 268210 150456
rect 265065 150451 265131 150454
rect 280654 150452 280660 150516
rect 280724 150514 280730 150516
rect 281717 150514 281783 150517
rect 280724 150512 281783 150514
rect 280724 150456 281722 150512
rect 281778 150456 281783 150512
rect 280724 150454 281783 150456
rect 280724 150452 280730 150454
rect 281717 150451 281783 150454
rect 213177 150242 213243 150245
rect 213177 150240 217242 150242
rect 213177 150184 213182 150240
rect 213238 150184 217242 150240
rect 213177 150182 217242 150184
rect 213177 150179 213243 150182
rect -960 149834 480 149924
rect 3693 149834 3759 149837
rect -960 149832 3759 149834
rect -960 149776 3698 149832
rect 3754 149776 3759 149832
rect 217182 149804 217242 150182
rect 231761 150106 231827 150109
rect 228968 150104 231827 150106
rect 228968 150048 231766 150104
rect 231822 150048 231827 150104
rect 228968 150046 231827 150048
rect 231761 150043 231827 150046
rect 265341 150106 265407 150109
rect 268150 150106 268210 150348
rect 282821 150106 282887 150109
rect 265341 150104 268210 150106
rect 265341 150048 265346 150104
rect 265402 150048 268210 150104
rect 265341 150046 268210 150048
rect 279956 150104 282887 150106
rect 279956 150048 282826 150104
rect 282882 150048 282887 150104
rect 279956 150046 282887 150048
rect 265341 150043 265407 150046
rect 282821 150043 282887 150046
rect -960 149774 3759 149776
rect -960 149684 480 149774
rect 3693 149771 3759 149774
rect 230749 149698 230815 149701
rect 228968 149696 230815 149698
rect 228968 149640 230754 149696
rect 230810 149640 230815 149696
rect 228968 149638 230815 149640
rect 230749 149635 230815 149638
rect 265525 149698 265591 149701
rect 268150 149698 268210 149940
rect 279325 149834 279391 149837
rect 279325 149832 279434 149834
rect 279325 149776 279330 149832
rect 279386 149776 279434 149832
rect 279325 149771 279434 149776
rect 265525 149696 268210 149698
rect 265525 149640 265530 149696
rect 265586 149640 268210 149696
rect 265525 149638 268210 149640
rect 265525 149635 265591 149638
rect 213913 149562 213979 149565
rect 213913 149560 217242 149562
rect 213913 149504 213918 149560
rect 213974 149504 217242 149560
rect 213913 149502 217242 149504
rect 213913 149499 213979 149502
rect 217182 149124 217242 149502
rect 265801 149290 265867 149293
rect 268150 149290 268210 149532
rect 279374 149396 279434 149771
rect 265801 149288 268210 149290
rect 265801 149232 265806 149288
rect 265862 149232 268210 149288
rect 265801 149230 268210 149232
rect 265801 149227 265867 149230
rect 242934 149154 242940 149156
rect 228968 149094 242940 149154
rect 242934 149092 242940 149094
rect 243004 149092 243010 149156
rect 213913 148746 213979 148749
rect 231209 148746 231275 148749
rect 213913 148744 217242 148746
rect 213913 148688 213918 148744
rect 213974 148688 217242 148744
rect 213913 148686 217242 148688
rect 228968 148744 231275 148746
rect 228968 148688 231214 148744
rect 231270 148688 231275 148744
rect 228968 148686 231275 148688
rect 213913 148683 213979 148686
rect 217182 148444 217242 148686
rect 231209 148683 231275 148686
rect 266077 148746 266143 148749
rect 268150 148746 268210 148988
rect 266077 148744 268210 148746
rect 266077 148688 266082 148744
rect 266138 148688 268210 148744
rect 266077 148686 268210 148688
rect 266077 148683 266143 148686
rect 282821 148610 282887 148613
rect 279956 148608 282887 148610
rect 265893 148338 265959 148341
rect 268150 148338 268210 148580
rect 279956 148552 282826 148608
rect 282882 148552 282887 148608
rect 279956 148550 282887 148552
rect 282821 148547 282887 148550
rect 265893 148336 268210 148338
rect 265893 148280 265898 148336
rect 265954 148280 268210 148336
rect 265893 148278 268210 148280
rect 265893 148275 265959 148278
rect 231761 148202 231827 148205
rect 228968 148200 231827 148202
rect 228968 148144 231766 148200
rect 231822 148144 231827 148200
rect 228968 148142 231827 148144
rect 231761 148139 231827 148142
rect 213913 148066 213979 148069
rect 213913 148064 217242 148066
rect 213913 148008 213918 148064
rect 213974 148008 217242 148064
rect 213913 148006 217242 148008
rect 213913 148003 213979 148006
rect 217182 147900 217242 148006
rect 265249 147930 265315 147933
rect 268334 147932 268394 148172
rect 265249 147928 268210 147930
rect 265249 147872 265254 147928
rect 265310 147872 268210 147928
rect 265249 147870 268210 147872
rect 265249 147867 265315 147870
rect 231945 147794 232011 147797
rect 228968 147792 232011 147794
rect 228968 147736 231950 147792
rect 232006 147736 232011 147792
rect 268150 147764 268210 147870
rect 268326 147868 268332 147932
rect 268396 147868 268402 147932
rect 282085 147794 282151 147797
rect 279956 147792 282151 147794
rect 228968 147734 232011 147736
rect 279956 147736 282090 147792
rect 282146 147736 282151 147792
rect 279956 147734 282151 147736
rect 231945 147731 232011 147734
rect 282085 147731 282151 147734
rect 231761 147250 231827 147253
rect 228968 147248 231827 147250
rect 214005 146706 214071 146709
rect 217182 146706 217242 147220
rect 228968 147192 231766 147248
rect 231822 147192 231827 147248
rect 228968 147190 231827 147192
rect 231761 147187 231827 147190
rect 265525 147114 265591 147117
rect 268150 147114 268210 147356
rect 285622 147114 285628 147116
rect 265525 147112 268210 147114
rect 265525 147056 265530 147112
rect 265586 147056 268210 147112
rect 265525 147054 268210 147056
rect 279956 147054 285628 147114
rect 265525 147051 265591 147054
rect 285622 147052 285628 147054
rect 285692 147052 285698 147116
rect 230565 146842 230631 146845
rect 228968 146840 230631 146842
rect 228968 146784 230570 146840
rect 230626 146784 230631 146840
rect 228968 146782 230631 146784
rect 230565 146779 230631 146782
rect 214005 146704 217242 146706
rect 214005 146648 214010 146704
rect 214066 146648 217242 146704
rect 214005 146646 217242 146648
rect 265893 146706 265959 146709
rect 268150 146706 268210 146948
rect 265893 146704 268210 146706
rect 265893 146648 265898 146704
rect 265954 146648 268210 146704
rect 265893 146646 268210 146648
rect 214005 146643 214071 146646
rect 265893 146643 265959 146646
rect 265801 146570 265867 146573
rect 265801 146568 268210 146570
rect 213913 146434 213979 146437
rect 213913 146432 216874 146434
rect 213913 146376 213918 146432
rect 213974 146376 216874 146432
rect 213913 146374 216874 146376
rect 213913 146371 213979 146374
rect 216814 146298 216874 146374
rect 217366 146298 217426 146540
rect 265801 146512 265806 146568
rect 265862 146512 268210 146568
rect 265801 146510 268210 146512
rect 265801 146507 265867 146510
rect 268150 146404 268210 146510
rect 231669 146298 231735 146301
rect 282821 146298 282887 146301
rect 216814 146238 217426 146298
rect 228968 146296 231735 146298
rect 228968 146240 231674 146296
rect 231730 146240 231735 146296
rect 228968 146238 231735 146240
rect 279956 146296 282887 146298
rect 279956 146240 282826 146296
rect 282882 146240 282887 146296
rect 279956 146238 282887 146240
rect 231669 146235 231735 146238
rect 282821 146235 282887 146238
rect 265341 146162 265407 146165
rect 268326 146162 268332 146164
rect 265341 146160 268332 146162
rect 265341 146104 265346 146160
rect 265402 146104 268332 146160
rect 265341 146102 268332 146104
rect 265341 146099 265407 146102
rect 268326 146100 268332 146102
rect 268396 146100 268402 146164
rect 230841 145890 230907 145893
rect 228968 145888 230907 145890
rect 214005 145346 214071 145349
rect 217182 145346 217242 145860
rect 228968 145832 230846 145888
rect 230902 145832 230907 145888
rect 228968 145830 230907 145832
rect 230841 145827 230907 145830
rect 265893 145754 265959 145757
rect 268150 145754 268210 145996
rect 265893 145752 268210 145754
rect 265893 145696 265898 145752
rect 265954 145696 268210 145752
rect 265893 145694 268210 145696
rect 265893 145691 265959 145694
rect 231301 145346 231367 145349
rect 214005 145344 217242 145346
rect 214005 145288 214010 145344
rect 214066 145288 217242 145344
rect 214005 145286 217242 145288
rect 228968 145344 231367 145346
rect 228968 145288 231306 145344
rect 231362 145288 231367 145344
rect 228968 145286 231367 145288
rect 214005 145283 214071 145286
rect 231301 145283 231367 145286
rect 265157 145346 265223 145349
rect 268150 145346 268210 145588
rect 284886 145482 284892 145484
rect 279956 145422 284892 145482
rect 284886 145420 284892 145422
rect 284956 145420 284962 145484
rect 265157 145344 268210 145346
rect 265157 145288 265162 145344
rect 265218 145288 268210 145344
rect 265157 145286 268210 145288
rect 265157 145283 265223 145286
rect 213913 144938 213979 144941
rect 217366 144938 217426 145180
rect 231117 144938 231183 144941
rect 213913 144936 217426 144938
rect 213913 144880 213918 144936
rect 213974 144880 217426 144936
rect 213913 144878 217426 144880
rect 228968 144936 231183 144938
rect 228968 144880 231122 144936
rect 231178 144880 231183 144936
rect 228968 144878 231183 144880
rect 213913 144875 213979 144878
rect 231117 144875 231183 144878
rect 265801 144938 265867 144941
rect 268334 144938 268394 145180
rect 265801 144936 268394 144938
rect 265801 144880 265806 144936
rect 265862 144880 268394 144936
rect 265801 144878 268394 144880
rect 265801 144875 265867 144878
rect 284702 144802 284708 144804
rect 265341 144530 265407 144533
rect 268150 144530 268210 144772
rect 279956 144742 284708 144802
rect 284702 144740 284708 144742
rect 284772 144740 284778 144804
rect 265341 144528 268210 144530
rect 214465 143986 214531 143989
rect 217182 143986 217242 144500
rect 265341 144472 265346 144528
rect 265402 144472 268210 144528
rect 265341 144470 268210 144472
rect 265341 144467 265407 144470
rect 231301 144394 231367 144397
rect 228968 144392 231367 144394
rect 228968 144336 231306 144392
rect 231362 144336 231367 144392
rect 228968 144334 231367 144336
rect 231301 144331 231367 144334
rect 265801 144122 265867 144125
rect 268150 144122 268210 144364
rect 265801 144120 268210 144122
rect 265801 144064 265806 144120
rect 265862 144064 268210 144120
rect 265801 144062 268210 144064
rect 265801 144059 265867 144062
rect 231761 143986 231827 143989
rect 281901 143986 281967 143989
rect 214465 143984 217242 143986
rect 214465 143928 214470 143984
rect 214526 143928 217242 143984
rect 214465 143926 217242 143928
rect 228968 143984 231827 143986
rect 228968 143928 231766 143984
rect 231822 143928 231827 143984
rect 228968 143926 231827 143928
rect 279956 143984 281967 143986
rect 279956 143928 281906 143984
rect 281962 143928 281967 143984
rect 279956 143926 281967 143928
rect 214465 143923 214531 143926
rect 231761 143923 231827 143926
rect 281901 143923 281967 143926
rect 213913 143578 213979 143581
rect 217366 143578 217426 143820
rect 213913 143576 217426 143578
rect 213913 143520 213918 143576
rect 213974 143520 217426 143576
rect 213913 143518 217426 143520
rect 265525 143578 265591 143581
rect 268150 143578 268210 143820
rect 265525 143576 268210 143578
rect 265525 143520 265530 143576
rect 265586 143520 268210 143576
rect 265525 143518 268210 143520
rect 213913 143515 213979 143518
rect 265525 143515 265591 143518
rect 231761 143442 231827 143445
rect 228968 143440 231827 143442
rect 228968 143384 231766 143440
rect 231822 143384 231827 143440
rect 228968 143382 231827 143384
rect 231761 143379 231827 143382
rect 214005 142762 214071 142765
rect 217182 142762 217242 143276
rect 265157 143170 265223 143173
rect 268150 143170 268210 143412
rect 284518 143170 284524 143172
rect 265157 143168 268210 143170
rect 265157 143112 265162 143168
rect 265218 143112 268210 143168
rect 265157 143110 268210 143112
rect 279956 143110 284524 143170
rect 265157 143107 265223 143110
rect 284518 143108 284524 143110
rect 284588 143108 284594 143172
rect 231301 143034 231367 143037
rect 228968 143032 231367 143034
rect 228968 142976 231306 143032
rect 231362 142976 231367 143032
rect 228968 142974 231367 142976
rect 231301 142971 231367 142974
rect 214005 142760 217242 142762
rect 214005 142704 214010 142760
rect 214066 142704 217242 142760
rect 214005 142702 217242 142704
rect 266169 142762 266235 142765
rect 268150 142762 268210 143004
rect 266169 142760 268210 142762
rect 266169 142704 266174 142760
rect 266230 142704 268210 142760
rect 266169 142702 268210 142704
rect 214005 142699 214071 142702
rect 266169 142699 266235 142702
rect 213913 142354 213979 142357
rect 217182 142354 217242 142596
rect 231669 142490 231735 142493
rect 228968 142488 231735 142490
rect 228968 142432 231674 142488
rect 231730 142432 231735 142488
rect 228968 142430 231735 142432
rect 231669 142427 231735 142430
rect 213913 142352 217242 142354
rect 213913 142296 213918 142352
rect 213974 142296 217242 142352
rect 213913 142294 217242 142296
rect 266077 142354 266143 142357
rect 268518 142356 268578 142596
rect 282821 142490 282887 142493
rect 279956 142488 282887 142490
rect 279956 142432 282826 142488
rect 282882 142432 282887 142488
rect 279956 142430 282887 142432
rect 282821 142427 282887 142430
rect 266077 142352 268210 142354
rect 266077 142296 266082 142352
rect 266138 142296 268210 142352
rect 266077 142294 268210 142296
rect 213913 142291 213979 142294
rect 266077 142291 266143 142294
rect 268150 142188 268210 142294
rect 268510 142292 268516 142356
rect 268580 142292 268586 142356
rect 231761 142082 231827 142085
rect 228968 142080 231827 142082
rect 228968 142024 231766 142080
rect 231822 142024 231827 142080
rect 228968 142022 231827 142024
rect 231761 142019 231827 142022
rect 261569 141946 261635 141949
rect 268510 141946 268516 141948
rect 261569 141944 268516 141946
rect 214005 141402 214071 141405
rect 217182 141402 217242 141916
rect 261569 141888 261574 141944
rect 261630 141888 268516 141944
rect 261569 141886 268516 141888
rect 261569 141883 261635 141886
rect 268510 141884 268516 141886
rect 268580 141884 268586 141948
rect 231761 141674 231827 141677
rect 228968 141672 231827 141674
rect 228968 141616 231766 141672
rect 231822 141616 231827 141672
rect 228968 141614 231827 141616
rect 231761 141611 231827 141614
rect 214005 141400 217242 141402
rect 214005 141344 214010 141400
rect 214066 141344 217242 141400
rect 214005 141342 217242 141344
rect 265801 141402 265867 141405
rect 268150 141402 268210 141780
rect 280613 141674 280679 141677
rect 279956 141672 280679 141674
rect 279956 141616 280618 141672
rect 280674 141616 280679 141672
rect 279956 141614 280679 141616
rect 280613 141611 280679 141614
rect 265801 141400 268210 141402
rect 265801 141344 265806 141400
rect 265862 141344 268210 141400
rect 265801 141342 268210 141344
rect 214005 141339 214071 141342
rect 265801 141339 265867 141342
rect 213913 140994 213979 140997
rect 217182 140994 217242 141236
rect 231393 141130 231459 141133
rect 228968 141128 231459 141130
rect 228968 141072 231398 141128
rect 231454 141072 231459 141128
rect 228968 141070 231459 141072
rect 231393 141067 231459 141070
rect 213913 140992 217242 140994
rect 213913 140936 213918 140992
rect 213974 140936 217242 140992
rect 213913 140934 217242 140936
rect 265893 140994 265959 140997
rect 268150 140994 268210 141236
rect 265893 140992 268210 140994
rect 265893 140936 265898 140992
rect 265954 140936 268210 140992
rect 265893 140934 268210 140936
rect 213913 140931 213979 140934
rect 265893 140931 265959 140934
rect 265985 140858 266051 140861
rect 284334 140858 284340 140860
rect 265985 140856 267842 140858
rect 265985 140800 265990 140856
rect 266046 140800 267842 140856
rect 265985 140798 267842 140800
rect 265985 140795 266051 140798
rect 230422 140722 230428 140724
rect 228968 140662 230428 140722
rect 230422 140660 230428 140662
rect 230492 140660 230498 140724
rect 267782 140586 267842 140798
rect 268334 140586 268394 140828
rect 279956 140798 284340 140858
rect 284334 140796 284340 140798
rect 284404 140796 284410 140860
rect 214005 140042 214071 140045
rect 217182 140042 217242 140556
rect 267782 140526 268394 140586
rect 231209 140178 231275 140181
rect 228968 140176 231275 140178
rect 228968 140120 231214 140176
rect 231270 140120 231275 140176
rect 228968 140118 231275 140120
rect 231209 140115 231275 140118
rect 264237 140178 264303 140181
rect 268150 140178 268210 140420
rect 282821 140178 282887 140181
rect 264237 140176 268210 140178
rect 264237 140120 264242 140176
rect 264298 140120 268210 140176
rect 264237 140118 268210 140120
rect 279956 140176 282887 140178
rect 279956 140120 282826 140176
rect 282882 140120 282887 140176
rect 279956 140118 282887 140120
rect 264237 140115 264303 140118
rect 282821 140115 282887 140118
rect 214005 140040 217242 140042
rect 214005 139984 214010 140040
rect 214066 139984 217242 140040
rect 214005 139982 217242 139984
rect 214005 139979 214071 139982
rect 213913 139634 213979 139637
rect 217182 139634 217242 139876
rect 231761 139770 231827 139773
rect 228968 139768 231827 139770
rect 228968 139712 231766 139768
rect 231822 139712 231827 139768
rect 228968 139710 231827 139712
rect 231761 139707 231827 139710
rect 265893 139770 265959 139773
rect 268150 139770 268210 140012
rect 265893 139768 268210 139770
rect 265893 139712 265898 139768
rect 265954 139712 268210 139768
rect 265893 139710 268210 139712
rect 265893 139707 265959 139710
rect 213913 139632 217242 139634
rect 213913 139576 213918 139632
rect 213974 139576 217242 139632
rect 213913 139574 217242 139576
rect 213913 139571 213979 139574
rect 265801 139498 265867 139501
rect 265801 139496 267842 139498
rect 265801 139440 265806 139496
rect 265862 139440 267842 139496
rect 265801 139438 267842 139440
rect 265801 139435 265867 139438
rect 267782 139362 267842 139438
rect 268334 139362 268394 139604
rect 282729 139362 282795 139365
rect 267782 139302 268394 139362
rect 279956 139360 282795 139362
rect 279956 139304 282734 139360
rect 282790 139304 282795 139360
rect 279956 139302 282795 139304
rect 282729 139299 282795 139302
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 231761 139226 231827 139229
rect 228968 139224 231827 139226
rect 217182 138818 217242 139196
rect 228968 139168 231766 139224
rect 231822 139168 231827 139224
rect 583520 139212 584960 139302
rect 228968 139166 231827 139168
rect 231761 139163 231827 139166
rect 231301 138818 231367 138821
rect 200070 138758 217242 138818
rect 228968 138816 231367 138818
rect 228968 138760 231306 138816
rect 231362 138760 231367 138816
rect 228968 138758 231367 138760
rect 164918 138212 164924 138276
rect 164988 138274 164994 138276
rect 200070 138274 200130 138758
rect 231301 138755 231367 138758
rect 265985 138818 266051 138821
rect 268150 138818 268210 139196
rect 265985 138816 268210 138818
rect 265985 138760 265990 138816
rect 266046 138760 268210 138816
rect 265985 138758 268210 138760
rect 265985 138755 266051 138758
rect 164988 138214 200130 138274
rect 164988 138212 164994 138214
rect 214833 138138 214899 138141
rect 217182 138138 217242 138652
rect 265433 138410 265499 138413
rect 268150 138410 268210 138652
rect 282821 138546 282887 138549
rect 279956 138544 282887 138546
rect 279956 138488 282826 138544
rect 282882 138488 282887 138544
rect 279956 138486 282887 138488
rect 282821 138483 282887 138486
rect 265433 138408 268210 138410
rect 265433 138352 265438 138408
rect 265494 138352 268210 138408
rect 265433 138350 268210 138352
rect 265433 138347 265499 138350
rect 230933 138274 230999 138277
rect 228968 138272 230999 138274
rect 228968 138216 230938 138272
rect 230994 138216 230999 138272
rect 228968 138214 230999 138216
rect 230933 138211 230999 138214
rect 214833 138136 217242 138138
rect 214833 138080 214838 138136
rect 214894 138080 217242 138136
rect 214833 138078 217242 138080
rect 265525 138138 265591 138141
rect 265525 138136 267842 138138
rect 265525 138080 265530 138136
rect 265586 138080 267842 138136
rect 265525 138078 267842 138080
rect 214833 138075 214899 138078
rect 265525 138075 265591 138078
rect 267782 138002 267842 138078
rect 268334 138002 268394 138244
rect 217182 137458 217242 137972
rect 267782 137942 268394 138002
rect 231761 137866 231827 137869
rect 281625 137866 281691 137869
rect 228968 137864 231827 137866
rect 228968 137808 231766 137864
rect 231822 137808 231827 137864
rect 279956 137864 281691 137866
rect 228968 137806 231827 137808
rect 231761 137803 231827 137806
rect 265433 137594 265499 137597
rect 268150 137594 268210 137836
rect 279956 137808 281630 137864
rect 281686 137808 281691 137864
rect 279956 137806 281691 137808
rect 281625 137803 281691 137806
rect 265433 137592 268210 137594
rect 265433 137536 265438 137592
rect 265494 137536 268210 137592
rect 265433 137534 268210 137536
rect 265433 137531 265499 137534
rect 200070 137398 217242 137458
rect -960 136778 480 136868
rect 166206 136852 166212 136916
rect 166276 136914 166282 136916
rect 200070 136914 200130 137398
rect 231669 137322 231735 137325
rect 228968 137320 231735 137322
rect 166276 136854 200130 136914
rect 166276 136852 166282 136854
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 213913 136778 213979 136781
rect 217182 136778 217242 137292
rect 228968 137264 231674 137320
rect 231730 137264 231735 137320
rect 228968 137262 231735 137264
rect 231669 137259 231735 137262
rect 265525 137186 265591 137189
rect 268150 137186 268210 137428
rect 265525 137184 268210 137186
rect 265525 137128 265530 137184
rect 265586 137128 268210 137184
rect 265525 137126 268210 137128
rect 265525 137123 265591 137126
rect 282269 137050 282335 137053
rect 279956 137048 282335 137050
rect 229645 136914 229711 136917
rect 228968 136912 229711 136914
rect 228968 136856 229650 136912
rect 229706 136856 229711 136912
rect 228968 136854 229711 136856
rect 229645 136851 229711 136854
rect 213913 136776 217242 136778
rect 213913 136720 213918 136776
rect 213974 136720 217242 136776
rect 213913 136718 217242 136720
rect 265985 136778 266051 136781
rect 268150 136778 268210 137020
rect 279956 136992 282274 137048
rect 282330 136992 282335 137048
rect 279956 136990 282335 136992
rect 282269 136987 282335 136990
rect 265985 136776 268210 136778
rect 265985 136720 265990 136776
rect 266046 136720 268210 136776
rect 265985 136718 268210 136720
rect 213913 136715 213979 136718
rect 265985 136715 266051 136718
rect 214005 136098 214071 136101
rect 217182 136098 217242 136612
rect 233182 136370 233188 136372
rect 228968 136310 233188 136370
rect 233182 136308 233188 136310
rect 233252 136308 233258 136372
rect 265249 136370 265315 136373
rect 268150 136370 268210 136612
rect 265249 136368 268210 136370
rect 265249 136312 265254 136368
rect 265310 136312 268210 136368
rect 265249 136310 268210 136312
rect 265249 136307 265315 136310
rect 268326 136308 268332 136372
rect 268396 136308 268402 136372
rect 282821 136370 282887 136373
rect 279956 136368 282887 136370
rect 279956 136312 282826 136368
rect 282882 136312 282887 136368
rect 279956 136310 282887 136312
rect 268334 136204 268394 136308
rect 282821 136307 282887 136310
rect 214005 136096 217242 136098
rect 214005 136040 214010 136096
rect 214066 136040 217242 136096
rect 214005 136038 217242 136040
rect 214005 136035 214071 136038
rect 231393 135962 231459 135965
rect 228968 135960 231459 135962
rect 214097 135690 214163 135693
rect 217182 135690 217242 135932
rect 228968 135904 231398 135960
rect 231454 135904 231459 135960
rect 228968 135902 231459 135904
rect 231393 135899 231459 135902
rect 264513 135962 264579 135965
rect 264513 135960 268578 135962
rect 264513 135904 264518 135960
rect 264574 135904 268578 135960
rect 264513 135902 268578 135904
rect 264513 135899 264579 135902
rect 262581 135826 262647 135829
rect 268142 135826 268148 135828
rect 262581 135824 268148 135826
rect 262581 135768 262586 135824
rect 262642 135768 268148 135824
rect 262581 135766 268148 135768
rect 262581 135763 262647 135766
rect 268142 135764 268148 135766
rect 268212 135764 268218 135828
rect 214097 135688 217242 135690
rect 214097 135632 214102 135688
rect 214158 135632 217242 135688
rect 268518 135660 268578 135902
rect 214097 135630 217242 135632
rect 214097 135627 214163 135630
rect 282177 135554 282243 135557
rect 279956 135552 282243 135554
rect 279956 135496 282182 135552
rect 282238 135496 282243 135552
rect 279956 135494 282243 135496
rect 282177 135491 282243 135494
rect 213913 135418 213979 135421
rect 231761 135418 231827 135421
rect 213913 135416 217242 135418
rect 213913 135360 213918 135416
rect 213974 135360 217242 135416
rect 213913 135358 217242 135360
rect 228968 135416 231827 135418
rect 228968 135360 231766 135416
rect 231822 135360 231827 135416
rect 228968 135358 231827 135360
rect 213913 135355 213979 135358
rect 217182 135252 217242 135358
rect 231761 135355 231827 135358
rect 265985 135418 266051 135421
rect 265985 135416 268210 135418
rect 265985 135360 265990 135416
rect 266046 135360 268210 135416
rect 265985 135358 268210 135360
rect 265985 135355 266051 135358
rect 268150 135252 268210 135358
rect 231761 135010 231827 135013
rect 228968 135008 231827 135010
rect 228968 134952 231766 135008
rect 231822 134952 231827 135008
rect 228968 134950 231827 134952
rect 231761 134947 231827 134950
rect 265249 134602 265315 134605
rect 268150 134602 268210 134844
rect 282545 134738 282611 134741
rect 279956 134736 282611 134738
rect 279956 134680 282550 134736
rect 282606 134680 282611 134736
rect 279956 134678 282611 134680
rect 282545 134675 282611 134678
rect 265249 134600 268210 134602
rect 213913 134330 213979 134333
rect 217182 134330 217242 134572
rect 265249 134544 265254 134600
rect 265310 134544 268210 134600
rect 265249 134542 268210 134544
rect 265249 134539 265315 134542
rect 231669 134466 231735 134469
rect 228968 134464 231735 134466
rect 228968 134408 231674 134464
rect 231730 134408 231735 134464
rect 228968 134406 231735 134408
rect 231669 134403 231735 134406
rect 213913 134328 217242 134330
rect 213913 134272 213918 134328
rect 213974 134272 217242 134328
rect 213913 134270 217242 134272
rect 213913 134267 213979 134270
rect 215109 134194 215175 134197
rect 265985 134194 266051 134197
rect 268518 134196 268578 134436
rect 215109 134192 217426 134194
rect 215109 134136 215114 134192
rect 215170 134136 217426 134192
rect 215109 134134 217426 134136
rect 215109 134131 215175 134134
rect 217366 133892 217426 134134
rect 265985 134192 268210 134194
rect 265985 134136 265990 134192
rect 266046 134136 268210 134192
rect 265985 134134 268210 134136
rect 265985 134131 266051 134134
rect 231577 134058 231643 134061
rect 228968 134056 231643 134058
rect 228968 134000 231582 134056
rect 231638 134000 231643 134056
rect 268150 134028 268210 134134
rect 268510 134132 268516 134196
rect 268580 134132 268586 134196
rect 281809 134058 281875 134061
rect 279956 134056 281875 134058
rect 228968 133998 231643 134000
rect 279956 134000 281814 134056
rect 281870 134000 281875 134056
rect 279956 133998 281875 134000
rect 231577 133995 231643 133998
rect 281809 133995 281875 133998
rect 264513 133786 264579 133789
rect 268510 133786 268516 133788
rect 264513 133784 268516 133786
rect 264513 133728 264518 133784
rect 264574 133728 268516 133784
rect 264513 133726 268516 133728
rect 264513 133723 264579 133726
rect 268510 133724 268516 133726
rect 268580 133724 268586 133788
rect 230657 133514 230723 133517
rect 228968 133512 230723 133514
rect 228968 133456 230662 133512
rect 230718 133456 230723 133512
rect 228968 133454 230723 133456
rect 230657 133451 230723 133454
rect 214005 132834 214071 132837
rect 217182 132834 217242 133348
rect 266169 133242 266235 133245
rect 268150 133242 268210 133620
rect 282269 133242 282335 133245
rect 266169 133240 268210 133242
rect 266169 133184 266174 133240
rect 266230 133184 268210 133240
rect 266169 133182 268210 133184
rect 279956 133240 282335 133242
rect 279956 133184 282274 133240
rect 282330 133184 282335 133240
rect 279956 133182 282335 133184
rect 266169 133179 266235 133182
rect 282269 133179 282335 133182
rect 231761 133106 231827 133109
rect 228968 133104 231827 133106
rect 228968 133048 231766 133104
rect 231822 133048 231827 133104
rect 228968 133046 231827 133048
rect 231761 133043 231827 133046
rect 214005 132832 217242 132834
rect 214005 132776 214010 132832
rect 214066 132776 217242 132832
rect 214005 132774 217242 132776
rect 265157 132834 265223 132837
rect 268150 132834 268210 133076
rect 265157 132832 268210 132834
rect 265157 132776 265162 132832
rect 265218 132776 268210 132832
rect 265157 132774 268210 132776
rect 214005 132771 214071 132774
rect 265157 132771 265223 132774
rect 213913 132562 213979 132565
rect 213913 132560 216874 132562
rect 213913 132504 213918 132560
rect 213974 132510 216874 132560
rect 217366 132510 217426 132668
rect 231669 132562 231735 132565
rect 213974 132504 217426 132510
rect 213913 132502 217426 132504
rect 228968 132560 231735 132562
rect 228968 132504 231674 132560
rect 231730 132504 231735 132560
rect 228968 132502 231735 132504
rect 213913 132499 213979 132502
rect 216814 132450 217426 132502
rect 231669 132499 231735 132502
rect 265985 132562 266051 132565
rect 265985 132560 267842 132562
rect 265985 132504 265990 132560
rect 266046 132504 267842 132560
rect 265985 132502 267842 132504
rect 265985 132499 266051 132502
rect 267782 132426 267842 132502
rect 268334 132426 268394 132668
rect 282545 132426 282611 132429
rect 267782 132366 268394 132426
rect 279956 132424 282611 132426
rect 279956 132368 282550 132424
rect 282606 132368 282611 132424
rect 279956 132366 282611 132368
rect 282545 132363 282611 132366
rect 231761 132154 231827 132157
rect 228968 132152 231827 132154
rect 228968 132096 231766 132152
rect 231822 132096 231827 132152
rect 228968 132094 231827 132096
rect 231761 132091 231827 132094
rect 264513 132018 264579 132021
rect 268150 132018 268210 132260
rect 264513 132016 268210 132018
rect 214005 131474 214071 131477
rect 217182 131474 217242 131988
rect 264513 131960 264518 132016
rect 264574 131960 268210 132016
rect 264513 131958 268210 131960
rect 264513 131955 264579 131958
rect 231669 131610 231735 131613
rect 228968 131608 231735 131610
rect 228968 131552 231674 131608
rect 231730 131552 231735 131608
rect 228968 131550 231735 131552
rect 231669 131547 231735 131550
rect 265985 131610 266051 131613
rect 268150 131610 268210 131852
rect 282085 131746 282151 131749
rect 279956 131744 282151 131746
rect 279956 131688 282090 131744
rect 282146 131688 282151 131744
rect 279956 131686 282151 131688
rect 282085 131683 282151 131686
rect 265985 131608 268210 131610
rect 265985 131552 265990 131608
rect 266046 131552 268210 131608
rect 265985 131550 268210 131552
rect 265985 131547 266051 131550
rect 214005 131472 217242 131474
rect 214005 131416 214010 131472
rect 214066 131416 217242 131472
rect 214005 131414 217242 131416
rect 214005 131411 214071 131414
rect 213913 131202 213979 131205
rect 213913 131200 216874 131202
rect 213913 131144 213918 131200
rect 213974 131144 216874 131200
rect 213913 131142 216874 131144
rect 213913 131139 213979 131142
rect 216814 131066 216874 131142
rect 217366 131066 217426 131308
rect 231577 131202 231643 131205
rect 228968 131200 231643 131202
rect 228968 131144 231582 131200
rect 231638 131144 231643 131200
rect 228968 131142 231643 131144
rect 231577 131139 231643 131142
rect 266169 131202 266235 131205
rect 268334 131202 268394 131444
rect 266169 131200 268394 131202
rect 266169 131144 266174 131200
rect 266230 131144 268394 131200
rect 266169 131142 268394 131144
rect 266169 131139 266235 131142
rect 216814 131006 217426 131066
rect 231025 130658 231091 130661
rect 228968 130656 231091 130658
rect 214005 130114 214071 130117
rect 217182 130114 217242 130628
rect 228968 130600 231030 130656
rect 231086 130600 231091 130656
rect 228968 130598 231091 130600
rect 231025 130595 231091 130598
rect 266169 130658 266235 130661
rect 268150 130658 268210 131036
rect 281901 130930 281967 130933
rect 279956 130928 281967 130930
rect 279956 130872 281906 130928
rect 281962 130872 281967 130928
rect 279956 130870 281967 130872
rect 281901 130867 281967 130870
rect 266169 130656 268210 130658
rect 266169 130600 266174 130656
rect 266230 130600 268210 130656
rect 266169 130598 268210 130600
rect 266169 130595 266235 130598
rect 231485 130250 231551 130253
rect 228968 130248 231551 130250
rect 228968 130192 231490 130248
rect 231546 130192 231551 130248
rect 228968 130190 231551 130192
rect 231485 130187 231551 130190
rect 264329 130250 264395 130253
rect 268150 130250 268210 130492
rect 264329 130248 268210 130250
rect 264329 130192 264334 130248
rect 264390 130192 268210 130248
rect 264329 130190 268210 130192
rect 264329 130187 264395 130190
rect 282085 130114 282151 130117
rect 214005 130112 217242 130114
rect 214005 130056 214010 130112
rect 214066 130056 217242 130112
rect 279956 130112 282151 130114
rect 214005 130054 217242 130056
rect 214005 130051 214071 130054
rect 213913 129842 213979 129845
rect 213913 129840 216874 129842
rect 213913 129784 213918 129840
rect 213974 129784 216874 129840
rect 213913 129782 216874 129784
rect 213913 129779 213979 129782
rect 216814 129706 216874 129782
rect 217366 129706 217426 129948
rect 230933 129842 230999 129845
rect 228968 129840 230999 129842
rect 228968 129784 230938 129840
rect 230994 129784 230999 129840
rect 228968 129782 230999 129784
rect 230933 129779 230999 129782
rect 265985 129842 266051 129845
rect 268334 129842 268394 130084
rect 279956 130056 282090 130112
rect 282146 130056 282151 130112
rect 279956 130054 282151 130056
rect 282085 130051 282151 130054
rect 265985 129840 268394 129842
rect 265985 129784 265990 129840
rect 266046 129784 268394 129840
rect 265985 129782 268394 129784
rect 265985 129779 266051 129782
rect 216814 129646 217426 129706
rect 265525 129434 265591 129437
rect 268150 129434 268210 129676
rect 281901 129434 281967 129437
rect 265525 129432 268210 129434
rect 265525 129376 265530 129432
rect 265586 129376 268210 129432
rect 265525 129374 268210 129376
rect 279956 129432 281967 129434
rect 279956 129376 281906 129432
rect 281962 129376 281967 129432
rect 279956 129374 281967 129376
rect 265525 129371 265591 129374
rect 281901 129371 281967 129374
rect 66161 129298 66227 129301
rect 68142 129298 68816 129304
rect 231669 129298 231735 129301
rect 66161 129296 68816 129298
rect 66161 129240 66166 129296
rect 66222 129244 68816 129296
rect 228968 129296 231735 129298
rect 66222 129240 68202 129244
rect 66161 129238 68202 129240
rect 66161 129235 66227 129238
rect 214005 128890 214071 128893
rect 217182 128890 217242 129268
rect 228968 129240 231674 129296
rect 231730 129240 231735 129296
rect 228968 129238 231735 129240
rect 231669 129235 231735 129238
rect 265341 129026 265407 129029
rect 268150 129026 268210 129268
rect 265341 129024 268210 129026
rect 265341 128968 265346 129024
rect 265402 128968 268210 129024
rect 265341 128966 268210 128968
rect 265341 128963 265407 128966
rect 231761 128890 231827 128893
rect 214005 128888 217242 128890
rect 214005 128832 214010 128888
rect 214066 128832 217242 128888
rect 214005 128830 217242 128832
rect 228968 128888 231827 128890
rect 228968 128832 231766 128888
rect 231822 128832 231827 128888
rect 228968 128830 231827 128832
rect 214005 128827 214071 128830
rect 231761 128827 231827 128830
rect 213913 128482 213979 128485
rect 217182 128482 217242 128724
rect 265985 128618 266051 128621
rect 268150 128618 268210 128860
rect 282085 128618 282151 128621
rect 265985 128616 268210 128618
rect 265985 128560 265990 128616
rect 266046 128560 268210 128616
rect 265985 128558 268210 128560
rect 279956 128616 282151 128618
rect 279956 128560 282090 128616
rect 282146 128560 282151 128616
rect 279956 128558 282151 128560
rect 265985 128555 266051 128558
rect 282085 128555 282151 128558
rect 213913 128480 217242 128482
rect 213913 128424 213918 128480
rect 213974 128424 217242 128480
rect 213913 128422 217242 128424
rect 266169 128482 266235 128485
rect 266169 128480 268026 128482
rect 266169 128424 266174 128480
rect 266230 128424 268026 128480
rect 266169 128422 268026 128424
rect 213913 128419 213979 128422
rect 266169 128419 266235 128422
rect 231669 128346 231735 128349
rect 228968 128344 231735 128346
rect 228968 128288 231674 128344
rect 231730 128288 231735 128344
rect 228968 128286 231735 128288
rect 231669 128283 231735 128286
rect 267966 128210 268026 128422
rect 268150 128210 268210 128452
rect 267966 128150 268210 128210
rect 66069 128074 66135 128077
rect 68142 128074 68816 128080
rect 66069 128072 68816 128074
rect 66069 128016 66074 128072
rect 66130 128020 68816 128072
rect 66130 128016 68202 128020
rect 66069 128014 68202 128016
rect 66069 128011 66135 128014
rect 214005 127530 214071 127533
rect 217182 127530 217242 128044
rect 231761 127938 231827 127941
rect 228968 127936 231827 127938
rect 228968 127880 231766 127936
rect 231822 127880 231827 127936
rect 228968 127878 231827 127880
rect 231761 127875 231827 127878
rect 266169 127666 266235 127669
rect 268150 127666 268210 127908
rect 281901 127802 281967 127805
rect 279956 127800 281967 127802
rect 279956 127744 281906 127800
rect 281962 127744 281967 127800
rect 279956 127742 281967 127744
rect 281901 127739 281967 127742
rect 266169 127664 268210 127666
rect 266169 127608 266174 127664
rect 266230 127608 268210 127664
rect 266169 127606 268210 127608
rect 266169 127603 266235 127606
rect 214005 127528 217242 127530
rect 214005 127472 214010 127528
rect 214066 127472 217242 127528
rect 214005 127470 217242 127472
rect 214005 127467 214071 127470
rect 231577 127394 231643 127397
rect 228968 127392 231643 127394
rect 213913 127122 213979 127125
rect 217182 127122 217242 127364
rect 228968 127336 231582 127392
rect 231638 127336 231643 127392
rect 228968 127334 231643 127336
rect 231577 127331 231643 127334
rect 265525 127258 265591 127261
rect 268518 127260 268578 127500
rect 265525 127256 268210 127258
rect 265525 127200 265530 127256
rect 265586 127200 268210 127256
rect 265525 127198 268210 127200
rect 265525 127195 265591 127198
rect 213913 127120 217242 127122
rect 213913 127064 213918 127120
rect 213974 127064 217242 127120
rect 268150 127092 268210 127198
rect 268510 127196 268516 127260
rect 268580 127196 268586 127260
rect 281901 127122 281967 127125
rect 279956 127120 281967 127122
rect 213913 127062 217242 127064
rect 279956 127064 281906 127120
rect 281962 127064 281967 127120
rect 279956 127062 281967 127064
rect 213913 127059 213979 127062
rect 281901 127059 281967 127062
rect 231669 126986 231735 126989
rect 228968 126984 231735 126986
rect 228968 126928 231674 126984
rect 231730 126928 231735 126984
rect 228968 126926 231735 126928
rect 231669 126923 231735 126926
rect 264145 126850 264211 126853
rect 268510 126850 268516 126852
rect 264145 126848 268516 126850
rect 264145 126792 264150 126848
rect 264206 126792 268516 126848
rect 264145 126790 268516 126792
rect 264145 126787 264211 126790
rect 268510 126788 268516 126790
rect 268580 126788 268586 126852
rect 65977 126306 66043 126309
rect 68142 126306 68816 126312
rect 65977 126304 68816 126306
rect 65977 126248 65982 126304
rect 66038 126252 68816 126304
rect 66038 126248 68202 126252
rect 65977 126246 68202 126248
rect 65977 126243 66043 126246
rect 214005 126170 214071 126173
rect 217182 126170 217242 126684
rect 231761 126442 231827 126445
rect 228968 126440 231827 126442
rect 228968 126384 231766 126440
rect 231822 126384 231827 126440
rect 228968 126382 231827 126384
rect 231761 126379 231827 126382
rect 266169 126442 266235 126445
rect 268150 126442 268210 126684
rect 266169 126440 268210 126442
rect 266169 126384 266174 126440
rect 266230 126384 268210 126440
rect 266169 126382 268210 126384
rect 266169 126379 266235 126382
rect 282821 126306 282887 126309
rect 279956 126304 282887 126306
rect 214005 126168 217242 126170
rect 214005 126112 214010 126168
rect 214066 126112 217242 126168
rect 214005 126110 217242 126112
rect 214005 126107 214071 126110
rect 231577 126034 231643 126037
rect 228968 126032 231643 126034
rect 213913 125762 213979 125765
rect 217182 125762 217242 126004
rect 228968 125976 231582 126032
rect 231638 125976 231643 126032
rect 228968 125974 231643 125976
rect 231577 125971 231643 125974
rect 266261 126034 266327 126037
rect 268150 126034 268210 126276
rect 279956 126248 282826 126304
rect 282882 126248 282887 126304
rect 279956 126246 282887 126248
rect 282821 126243 282887 126246
rect 266261 126032 268210 126034
rect 266261 125976 266266 126032
rect 266322 125976 268210 126032
rect 266261 125974 268210 125976
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 266261 125971 266327 125974
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 213913 125760 217242 125762
rect 213913 125704 213918 125760
rect 213974 125704 217242 125760
rect 213913 125702 217242 125704
rect 213913 125699 213979 125702
rect 265525 125626 265591 125629
rect 268334 125626 268394 125868
rect 265525 125624 268394 125626
rect 265525 125568 265530 125624
rect 265586 125568 268394 125624
rect 265525 125566 268394 125568
rect 265525 125563 265591 125566
rect 231761 125490 231827 125493
rect 280153 125490 280219 125493
rect 228968 125488 231827 125490
rect 228968 125432 231766 125488
rect 231822 125432 231827 125488
rect 228968 125430 231827 125432
rect 279956 125488 280219 125490
rect 279956 125432 280158 125488
rect 280214 125432 280219 125488
rect 279956 125430 280219 125432
rect 231761 125427 231827 125430
rect 280153 125427 280219 125430
rect 67633 125218 67699 125221
rect 68142 125218 68816 125224
rect 67633 125216 68816 125218
rect 67633 125160 67638 125216
rect 67694 125164 68816 125216
rect 67694 125160 68202 125164
rect 67633 125158 68202 125160
rect 67633 125155 67699 125158
rect 214005 124810 214071 124813
rect 217182 124810 217242 125324
rect 231301 125082 231367 125085
rect 228968 125080 231367 125082
rect 228968 125024 231306 125080
rect 231362 125024 231367 125080
rect 228968 125022 231367 125024
rect 231301 125019 231367 125022
rect 266169 125082 266235 125085
rect 268150 125082 268210 125324
rect 266169 125080 268210 125082
rect 266169 125024 266174 125080
rect 266230 125024 268210 125080
rect 266169 125022 268210 125024
rect 266169 125019 266235 125022
rect 214005 124808 217242 124810
rect 214005 124752 214010 124808
rect 214066 124752 217242 124808
rect 214005 124750 217242 124752
rect 214005 124747 214071 124750
rect 265157 124674 265223 124677
rect 268150 124674 268210 124916
rect 282821 124810 282887 124813
rect 279956 124808 282887 124810
rect 279956 124752 282826 124808
rect 282882 124752 282887 124808
rect 279956 124750 282887 124752
rect 282821 124747 282887 124750
rect 265157 124672 268210 124674
rect 213913 124266 213979 124269
rect 217182 124266 217242 124644
rect 265157 124616 265162 124672
rect 265218 124616 268210 124672
rect 265157 124614 268210 124616
rect 265157 124611 265223 124614
rect 231117 124538 231183 124541
rect 228968 124536 231183 124538
rect 228968 124480 231122 124536
rect 231178 124480 231183 124536
rect 228968 124478 231183 124480
rect 231117 124475 231183 124478
rect 213913 124264 217242 124266
rect 213913 124208 213918 124264
rect 213974 124208 217242 124264
rect 213913 124206 217242 124208
rect 265341 124266 265407 124269
rect 268334 124266 268394 124508
rect 265341 124264 268394 124266
rect 265341 124208 265346 124264
rect 265402 124208 268394 124264
rect 265341 124206 268394 124208
rect 213913 124203 213979 124206
rect 265341 124203 265407 124206
rect 230841 124130 230907 124133
rect 228968 124128 230907 124130
rect -960 123572 480 123812
rect 65885 123586 65951 123589
rect 68142 123586 68816 123592
rect 65885 123584 68816 123586
rect 65885 123528 65890 123584
rect 65946 123532 68816 123584
rect 214005 123586 214071 123589
rect 217182 123586 217242 124100
rect 228968 124072 230846 124128
rect 230902 124072 230907 124128
rect 228968 124070 230907 124072
rect 230841 124067 230907 124070
rect 266169 123858 266235 123861
rect 268150 123858 268210 124100
rect 282821 123994 282887 123997
rect 279956 123992 282887 123994
rect 279956 123936 282826 123992
rect 282882 123936 282887 123992
rect 279956 123934 282887 123936
rect 282821 123931 282887 123934
rect 266169 123856 268210 123858
rect 266169 123800 266174 123856
rect 266230 123800 268210 123856
rect 266169 123798 268210 123800
rect 266169 123795 266235 123798
rect 231761 123586 231827 123589
rect 214005 123584 217242 123586
rect 65946 123528 68202 123532
rect 65885 123526 68202 123528
rect 214005 123528 214010 123584
rect 214066 123528 217242 123584
rect 214005 123526 217242 123528
rect 228968 123584 231827 123586
rect 228968 123528 231766 123584
rect 231822 123528 231827 123584
rect 228968 123526 231827 123528
rect 65885 123523 65951 123526
rect 214005 123523 214071 123526
rect 231761 123523 231827 123526
rect 265433 123450 265499 123453
rect 268150 123450 268210 123692
rect 265433 123448 268210 123450
rect 213913 123178 213979 123181
rect 217182 123178 217242 123420
rect 265433 123392 265438 123448
rect 265494 123392 268210 123448
rect 265433 123390 268210 123392
rect 265433 123387 265499 123390
rect 230749 123178 230815 123181
rect 213913 123176 217242 123178
rect 213913 123120 213918 123176
rect 213974 123120 217242 123176
rect 213913 123118 217242 123120
rect 228968 123176 230815 123178
rect 228968 123120 230754 123176
rect 230810 123120 230815 123176
rect 228968 123118 230815 123120
rect 213913 123115 213979 123118
rect 230749 123115 230815 123118
rect 265157 123042 265223 123045
rect 268518 123044 268578 123284
rect 281625 123178 281691 123181
rect 279956 123176 281691 123178
rect 279956 123120 281630 123176
rect 281686 123120 281691 123176
rect 279956 123118 281691 123120
rect 281625 123115 281691 123118
rect 265157 123040 268210 123042
rect 265157 122984 265162 123040
rect 265218 122984 268210 123040
rect 265157 122982 268210 122984
rect 265157 122979 265223 122982
rect 268150 122876 268210 122982
rect 268510 122980 268516 123044
rect 268580 122980 268586 123044
rect 65793 122634 65859 122637
rect 68142 122634 68816 122640
rect 65793 122632 68816 122634
rect 65793 122576 65798 122632
rect 65854 122580 68816 122632
rect 65854 122576 68202 122580
rect 65793 122574 68202 122576
rect 65793 122571 65859 122574
rect 214005 122226 214071 122229
rect 217182 122226 217242 122740
rect 231761 122634 231827 122637
rect 228968 122632 231827 122634
rect 228968 122576 231766 122632
rect 231822 122576 231827 122632
rect 228968 122574 231827 122576
rect 231761 122571 231827 122574
rect 264421 122634 264487 122637
rect 268510 122634 268516 122636
rect 264421 122632 268516 122634
rect 264421 122576 264426 122632
rect 264482 122576 268516 122632
rect 264421 122574 268516 122576
rect 264421 122571 264487 122574
rect 268510 122572 268516 122574
rect 268580 122572 268586 122636
rect 281533 122498 281599 122501
rect 279956 122496 281599 122498
rect 279956 122440 281538 122496
rect 281594 122440 281599 122496
rect 279956 122438 281599 122440
rect 281533 122435 281599 122438
rect 231117 122226 231183 122229
rect 214005 122224 217242 122226
rect 214005 122168 214010 122224
rect 214066 122168 217242 122224
rect 214005 122166 217242 122168
rect 228968 122224 231183 122226
rect 228968 122168 231122 122224
rect 231178 122168 231183 122224
rect 228968 122166 231183 122168
rect 214005 122163 214071 122166
rect 231117 122163 231183 122166
rect 264421 122090 264487 122093
rect 268150 122090 268210 122332
rect 264421 122088 268210 122090
rect 213913 121818 213979 121821
rect 217182 121818 217242 122060
rect 264421 122032 264426 122088
rect 264482 122032 268210 122088
rect 264421 122030 268210 122032
rect 264421 122027 264487 122030
rect 213913 121816 217242 121818
rect 213913 121760 213918 121816
rect 213974 121760 217242 121816
rect 213913 121758 217242 121760
rect 213913 121755 213979 121758
rect 231393 121682 231459 121685
rect 228968 121680 231459 121682
rect 228968 121624 231398 121680
rect 231454 121624 231459 121680
rect 228968 121622 231459 121624
rect 231393 121619 231459 121622
rect 265525 121682 265591 121685
rect 268518 121684 268578 121924
rect 265525 121680 268210 121682
rect 265525 121624 265530 121680
rect 265586 121624 268210 121680
rect 265525 121622 268210 121624
rect 265525 121619 265591 121622
rect 268150 121516 268210 121622
rect 268510 121620 268516 121684
rect 268580 121620 268586 121684
rect 280429 121682 280495 121685
rect 279956 121680 280495 121682
rect 279956 121624 280434 121680
rect 280490 121624 280495 121680
rect 279956 121622 280495 121624
rect 280429 121619 280495 121622
rect 67817 120866 67883 120869
rect 68142 120866 68816 120872
rect 67817 120864 68816 120866
rect 67817 120808 67822 120864
rect 67878 120812 68816 120864
rect 214005 120866 214071 120869
rect 217182 120866 217242 121380
rect 231485 121274 231551 121277
rect 228968 121272 231551 121274
rect 228968 121216 231490 121272
rect 231546 121216 231551 121272
rect 228968 121214 231551 121216
rect 231485 121211 231551 121214
rect 264697 121274 264763 121277
rect 268510 121274 268516 121276
rect 264697 121272 268516 121274
rect 264697 121216 264702 121272
rect 264758 121216 268516 121272
rect 264697 121214 268516 121216
rect 264697 121211 264763 121214
rect 268510 121212 268516 121214
rect 268580 121212 268586 121276
rect 214005 120864 217242 120866
rect 67878 120808 68202 120812
rect 67817 120806 68202 120808
rect 214005 120808 214010 120864
rect 214066 120808 217242 120864
rect 214005 120806 217242 120808
rect 265525 120866 265591 120869
rect 268150 120866 268210 121108
rect 280337 120866 280403 120869
rect 265525 120864 268210 120866
rect 265525 120808 265530 120864
rect 265586 120808 268210 120864
rect 265525 120806 268210 120808
rect 279956 120864 280403 120866
rect 279956 120808 280342 120864
rect 280398 120808 280403 120864
rect 279956 120806 280403 120808
rect 67817 120803 67883 120806
rect 214005 120803 214071 120806
rect 265525 120803 265591 120806
rect 280337 120803 280403 120806
rect 231761 120730 231827 120733
rect 228968 120728 231827 120730
rect 213913 120458 213979 120461
rect 217182 120458 217242 120700
rect 228968 120672 231766 120728
rect 231822 120672 231827 120728
rect 228968 120670 231827 120672
rect 231761 120667 231827 120670
rect 213913 120456 217242 120458
rect 213913 120400 213918 120456
rect 213974 120400 217242 120456
rect 213913 120398 217242 120400
rect 266169 120458 266235 120461
rect 268150 120458 268210 120700
rect 266169 120456 268210 120458
rect 266169 120400 266174 120456
rect 266230 120400 268210 120456
rect 266169 120398 268210 120400
rect 213913 120395 213979 120398
rect 266169 120395 266235 120398
rect 231393 120322 231459 120325
rect 228968 120320 231459 120322
rect 228968 120264 231398 120320
rect 231454 120264 231459 120320
rect 228968 120262 231459 120264
rect 231393 120259 231459 120262
rect 265433 120186 265499 120189
rect 265433 120184 267842 120186
rect 265433 120128 265438 120184
rect 265494 120128 267842 120184
rect 265433 120126 267842 120128
rect 265433 120123 265499 120126
rect 267782 120050 267842 120126
rect 268334 120050 268394 120292
rect 281717 120186 281783 120189
rect 279956 120184 281783 120186
rect 279956 120128 281722 120184
rect 281778 120128 281783 120184
rect 279956 120126 281783 120128
rect 281717 120123 281783 120126
rect 213913 119642 213979 119645
rect 217182 119642 217242 120020
rect 267782 119990 268394 120050
rect 231761 119778 231827 119781
rect 228968 119776 231827 119778
rect 228968 119720 231766 119776
rect 231822 119720 231827 119776
rect 228968 119718 231827 119720
rect 231761 119715 231827 119718
rect 213913 119640 217242 119642
rect 213913 119584 213918 119640
rect 213974 119584 217242 119640
rect 213913 119582 217242 119584
rect 213913 119579 213979 119582
rect 266169 119506 266235 119509
rect 268150 119506 268210 119748
rect 266169 119504 268210 119506
rect 214005 118962 214071 118965
rect 217182 118962 217242 119476
rect 266169 119448 266174 119504
rect 266230 119448 268210 119504
rect 266169 119446 268210 119448
rect 266169 119443 266235 119446
rect 231577 119370 231643 119373
rect 280521 119370 280587 119373
rect 228968 119368 231643 119370
rect 228968 119312 231582 119368
rect 231638 119312 231643 119368
rect 279956 119368 280587 119370
rect 228968 119310 231643 119312
rect 231577 119307 231643 119310
rect 265525 119098 265591 119101
rect 268150 119098 268210 119340
rect 279956 119312 280526 119368
rect 280582 119312 280587 119368
rect 279956 119310 280587 119312
rect 280521 119307 280587 119310
rect 265525 119096 268210 119098
rect 265525 119040 265530 119096
rect 265586 119040 268210 119096
rect 265525 119038 268210 119040
rect 265525 119035 265591 119038
rect 230565 118962 230631 118965
rect 214005 118960 217242 118962
rect 214005 118904 214010 118960
rect 214066 118904 217242 118960
rect 214005 118902 217242 118904
rect 228968 118960 230631 118962
rect 228968 118904 230570 118960
rect 230626 118904 230631 118960
rect 228968 118902 230631 118904
rect 214005 118899 214071 118902
rect 230565 118899 230631 118902
rect 213177 118826 213243 118829
rect 265433 118826 265499 118829
rect 213177 118824 216874 118826
rect 213177 118768 213182 118824
rect 213238 118768 216874 118824
rect 265433 118824 267842 118826
rect 213177 118766 216874 118768
rect 213177 118763 213243 118766
rect 216814 118554 216874 118766
rect 217366 118554 217426 118796
rect 265433 118768 265438 118824
rect 265494 118768 267842 118824
rect 265433 118766 267842 118768
rect 265433 118763 265499 118766
rect 267782 118690 267842 118766
rect 268334 118690 268394 118932
rect 267782 118630 268394 118690
rect 282729 118554 282795 118557
rect 216814 118494 217426 118554
rect 279956 118552 282795 118554
rect 230565 118418 230631 118421
rect 228968 118416 230631 118418
rect 228968 118360 230570 118416
rect 230626 118360 230631 118416
rect 228968 118358 230631 118360
rect 230565 118355 230631 118358
rect 265525 118282 265591 118285
rect 268150 118282 268210 118524
rect 279956 118496 282734 118552
rect 282790 118496 282795 118552
rect 279956 118494 282795 118496
rect 282729 118491 282795 118494
rect 265525 118280 268210 118282
rect 265525 118224 265530 118280
rect 265586 118224 268210 118280
rect 265525 118222 268210 118224
rect 265525 118219 265591 118222
rect 214833 117602 214899 117605
rect 217182 117602 217242 118116
rect 231761 118010 231827 118013
rect 228968 118008 231827 118010
rect 228968 117952 231766 118008
rect 231822 117952 231827 118008
rect 228968 117950 231827 117952
rect 231761 117947 231827 117950
rect 265893 117874 265959 117877
rect 268150 117874 268210 118116
rect 282821 117874 282887 117877
rect 265893 117872 268210 117874
rect 265893 117816 265898 117872
rect 265954 117816 268210 117872
rect 265893 117814 268210 117816
rect 279956 117872 282887 117874
rect 279956 117816 282826 117872
rect 282882 117816 282887 117872
rect 279956 117814 282887 117816
rect 265893 117811 265959 117814
rect 282821 117811 282887 117814
rect 214833 117600 217242 117602
rect 214833 117544 214838 117600
rect 214894 117544 217242 117600
rect 214833 117542 217242 117544
rect 214833 117539 214899 117542
rect 230749 117466 230815 117469
rect 228968 117464 230815 117466
rect 213913 117330 213979 117333
rect 213913 117328 216874 117330
rect 213913 117272 213918 117328
rect 213974 117272 216874 117328
rect 213913 117270 216874 117272
rect 213913 117267 213979 117270
rect 216814 117194 216874 117270
rect 217366 117194 217426 117436
rect 228968 117408 230754 117464
rect 230810 117408 230815 117464
rect 228968 117406 230815 117408
rect 230749 117403 230815 117406
rect 265801 117466 265867 117469
rect 268150 117466 268210 117708
rect 265801 117464 268210 117466
rect 265801 117408 265806 117464
rect 265862 117408 268210 117464
rect 265801 117406 268210 117408
rect 265801 117403 265867 117406
rect 216814 117134 217426 117194
rect 231761 117058 231827 117061
rect 228968 117056 231827 117058
rect 228968 117000 231766 117056
rect 231822 117000 231827 117056
rect 228968 116998 231827 117000
rect 231761 116995 231827 116998
rect 266077 116922 266143 116925
rect 268150 116922 268210 117164
rect 282821 117058 282887 117061
rect 279956 117056 282887 117058
rect 279956 117000 282826 117056
rect 282882 117000 282887 117056
rect 279956 116998 282887 117000
rect 282821 116995 282887 116998
rect 266077 116920 268210 116922
rect 266077 116864 266082 116920
rect 266138 116864 268210 116920
rect 266077 116862 268210 116864
rect 266077 116859 266143 116862
rect 214005 116242 214071 116245
rect 217182 116242 217242 116756
rect 231485 116514 231551 116517
rect 228968 116512 231551 116514
rect 228968 116456 231490 116512
rect 231546 116456 231551 116512
rect 228968 116454 231551 116456
rect 231485 116451 231551 116454
rect 265893 116514 265959 116517
rect 268150 116514 268210 116756
rect 265893 116512 268210 116514
rect 265893 116456 265898 116512
rect 265954 116456 268210 116512
rect 265893 116454 268210 116456
rect 265893 116451 265959 116454
rect 282821 116378 282887 116381
rect 279956 116376 282887 116378
rect 214005 116240 217242 116242
rect 214005 116184 214010 116240
rect 214066 116184 217242 116240
rect 214005 116182 217242 116184
rect 214005 116179 214071 116182
rect 231669 116106 231735 116109
rect 228968 116104 231735 116106
rect 213913 115970 213979 115973
rect 213913 115968 216874 115970
rect 213913 115912 213918 115968
rect 213974 115912 216874 115968
rect 213913 115910 216874 115912
rect 213913 115907 213979 115910
rect 216814 115834 216874 115910
rect 217366 115834 217426 116076
rect 228968 116048 231674 116104
rect 231730 116048 231735 116104
rect 228968 116046 231735 116048
rect 231669 116043 231735 116046
rect 265801 116106 265867 116109
rect 265801 116104 268210 116106
rect 265801 116048 265806 116104
rect 265862 116048 268210 116104
rect 265801 116046 268210 116048
rect 265801 116043 265867 116046
rect 264605 115970 264671 115973
rect 267774 115970 267780 115972
rect 264605 115968 267780 115970
rect 264605 115912 264610 115968
rect 264666 115912 267780 115968
rect 264605 115910 267780 115912
rect 264605 115907 264671 115910
rect 267774 115908 267780 115910
rect 267844 115908 267850 115972
rect 268150 115940 268210 116046
rect 268326 116044 268332 116108
rect 268396 116106 268402 116108
rect 268518 116106 268578 116348
rect 279956 116320 282826 116376
rect 282882 116320 282887 116376
rect 279956 116318 282887 116320
rect 282821 116315 282887 116318
rect 268396 116046 268578 116106
rect 268396 116044 268402 116046
rect 216814 115774 217426 115834
rect 231761 115562 231827 115565
rect 285806 115562 285812 115564
rect 228968 115560 231827 115562
rect 228968 115504 231766 115560
rect 231822 115504 231827 115560
rect 228968 115502 231827 115504
rect 231761 115499 231827 115502
rect 214005 115018 214071 115021
rect 217182 115018 217242 115396
rect 265893 115290 265959 115293
rect 268150 115290 268210 115532
rect 279956 115502 285812 115562
rect 285806 115500 285812 115502
rect 285876 115500 285882 115564
rect 265893 115288 268210 115290
rect 265893 115232 265898 115288
rect 265954 115232 268210 115288
rect 265893 115230 268210 115232
rect 265893 115227 265959 115230
rect 230933 115154 230999 115157
rect 228968 115152 230999 115154
rect 228968 115096 230938 115152
rect 230994 115096 230999 115152
rect 228968 115094 230999 115096
rect 230933 115091 230999 115094
rect 214005 115016 217242 115018
rect 214005 114960 214010 115016
rect 214066 114960 217242 115016
rect 214005 114958 217242 114960
rect 214005 114955 214071 114958
rect 266077 114882 266143 114885
rect 268150 114882 268210 115124
rect 266077 114880 268210 114882
rect 213913 114610 213979 114613
rect 217182 114610 217242 114852
rect 266077 114824 266082 114880
rect 266138 114824 268210 114880
rect 266077 114822 268210 114824
rect 266077 114819 266143 114822
rect 265801 114746 265867 114749
rect 282821 114746 282887 114749
rect 265801 114744 268210 114746
rect 265801 114688 265806 114744
rect 265862 114688 268210 114744
rect 265801 114686 268210 114688
rect 279956 114744 282887 114746
rect 279956 114688 282826 114744
rect 282882 114688 282887 114744
rect 279956 114686 282887 114688
rect 265801 114683 265867 114686
rect 231301 114610 231367 114613
rect 213913 114608 217242 114610
rect 213913 114552 213918 114608
rect 213974 114552 217242 114608
rect 213913 114550 217242 114552
rect 228968 114608 231367 114610
rect 228968 114552 231306 114608
rect 231362 114552 231367 114608
rect 268150 114580 268210 114686
rect 282821 114683 282887 114686
rect 228968 114550 231367 114552
rect 213913 114547 213979 114550
rect 231301 114547 231367 114550
rect 231025 114202 231091 114205
rect 228968 114200 231091 114202
rect 214005 113658 214071 113661
rect 217182 113658 217242 114172
rect 228968 114144 231030 114200
rect 231086 114144 231091 114200
rect 228968 114142 231091 114144
rect 231025 114139 231091 114142
rect 265893 113930 265959 113933
rect 268150 113930 268210 114172
rect 282729 114066 282795 114069
rect 279956 114064 282795 114066
rect 279956 114008 282734 114064
rect 282790 114008 282795 114064
rect 279956 114006 282795 114008
rect 282729 114003 282795 114006
rect 265893 113928 268210 113930
rect 265893 113872 265898 113928
rect 265954 113872 268210 113928
rect 265893 113870 268210 113872
rect 265893 113867 265959 113870
rect 231485 113658 231551 113661
rect 214005 113656 217242 113658
rect 214005 113600 214010 113656
rect 214066 113600 217242 113656
rect 214005 113598 217242 113600
rect 228968 113656 231551 113658
rect 228968 113600 231490 113656
rect 231546 113600 231551 113656
rect 228968 113598 231551 113600
rect 214005 113595 214071 113598
rect 231485 113595 231551 113598
rect 265801 113522 265867 113525
rect 268150 113522 268210 113764
rect 265801 113520 268210 113522
rect 213913 113250 213979 113253
rect 217182 113250 217242 113492
rect 265801 113464 265806 113520
rect 265862 113464 268210 113520
rect 265801 113462 268210 113464
rect 265801 113459 265867 113462
rect 231761 113250 231827 113253
rect 213913 113248 217242 113250
rect 213913 113192 213918 113248
rect 213974 113192 217242 113248
rect 213913 113190 217242 113192
rect 228968 113248 231827 113250
rect 228968 113192 231766 113248
rect 231822 113192 231827 113248
rect 228968 113190 231827 113192
rect 213913 113187 213979 113190
rect 231761 113187 231827 113190
rect 265801 113250 265867 113253
rect 265801 113248 267842 113250
rect 265801 113192 265806 113248
rect 265862 113192 267842 113248
rect 265801 113190 267842 113192
rect 265801 113187 265867 113190
rect 267782 113114 267842 113190
rect 268334 113114 268394 113356
rect 282821 113250 282887 113253
rect 279956 113248 282887 113250
rect 279956 113192 282826 113248
rect 282882 113192 282887 113248
rect 279956 113190 282887 113192
rect 282821 113187 282887 113190
rect 267782 113054 268394 113114
rect 214005 112298 214071 112301
rect 217182 112298 217242 112812
rect 231761 112706 231827 112709
rect 228968 112704 231827 112706
rect 228968 112648 231766 112704
rect 231822 112648 231827 112704
rect 228968 112646 231827 112648
rect 231761 112643 231827 112646
rect 265893 112706 265959 112709
rect 268150 112706 268210 112948
rect 583520 112842 584960 112932
rect 265893 112704 268210 112706
rect 265893 112648 265898 112704
rect 265954 112648 268210 112704
rect 265893 112646 268210 112648
rect 583342 112782 584960 112842
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 265893 112643 265959 112646
rect 231669 112298 231735 112301
rect 214005 112296 217242 112298
rect 214005 112240 214010 112296
rect 214066 112240 217242 112296
rect 214005 112238 217242 112240
rect 228968 112296 231735 112298
rect 228968 112240 231674 112296
rect 231730 112240 231735 112296
rect 228968 112238 231735 112240
rect 214005 112235 214071 112238
rect 231669 112235 231735 112238
rect 265525 112298 265591 112301
rect 268150 112298 268210 112540
rect 282821 112434 282887 112437
rect 279956 112432 282887 112434
rect 279956 112376 282826 112432
rect 282882 112376 282887 112432
rect 279956 112374 282887 112376
rect 282821 112371 282887 112374
rect 265525 112296 268210 112298
rect 265525 112240 265530 112296
rect 265586 112240 268210 112296
rect 265525 112238 268210 112240
rect 265525 112235 265591 112238
rect 265801 112162 265867 112165
rect 265801 112160 268210 112162
rect 213913 111890 213979 111893
rect 217366 111890 217426 112132
rect 265801 112104 265806 112160
rect 265862 112104 268210 112160
rect 265801 112102 268210 112104
rect 265801 112099 265867 112102
rect 268150 111996 268210 112102
rect 213913 111888 217426 111890
rect 213913 111832 213918 111888
rect 213974 111832 217426 111888
rect 213913 111830 217426 111832
rect 213913 111827 213979 111830
rect 287646 111828 287652 111892
rect 287716 111890 287722 111892
rect 583526 111890 583586 112646
rect 287716 111830 583586 111890
rect 287716 111828 287722 111830
rect 168281 111754 168347 111757
rect 231761 111754 231827 111757
rect 281993 111754 282059 111757
rect 164694 111752 168347 111754
rect 164694 111696 168286 111752
rect 168342 111696 168347 111752
rect 164694 111694 168347 111696
rect 228968 111752 231827 111754
rect 228968 111696 231766 111752
rect 231822 111696 231827 111752
rect 228968 111694 231827 111696
rect 279956 111752 282059 111754
rect 279956 111696 281998 111752
rect 282054 111696 282059 111752
rect 279956 111694 282059 111696
rect 168281 111691 168347 111694
rect 231761 111691 231827 111694
rect 281993 111691 282059 111694
rect 215017 110938 215083 110941
rect 217182 110938 217242 111452
rect 231577 111346 231643 111349
rect 228968 111344 231643 111346
rect 228968 111288 231582 111344
rect 231638 111288 231643 111344
rect 228968 111286 231643 111288
rect 231577 111283 231643 111286
rect 265893 111346 265959 111349
rect 268150 111346 268210 111588
rect 265893 111344 268210 111346
rect 265893 111288 265898 111344
rect 265954 111288 268210 111344
rect 265893 111286 268210 111288
rect 265893 111283 265959 111286
rect 215017 110936 217242 110938
rect 215017 110880 215022 110936
rect 215078 110880 217242 110936
rect 215017 110878 217242 110880
rect 265157 110938 265223 110941
rect 268150 110938 268210 111180
rect 282821 110938 282887 110941
rect 265157 110936 268210 110938
rect 265157 110880 265162 110936
rect 265218 110880 268210 110936
rect 265157 110878 268210 110880
rect 279956 110936 282887 110938
rect 279956 110880 282826 110936
rect 282882 110880 282887 110936
rect 279956 110878 282887 110880
rect 215017 110875 215083 110878
rect 265157 110875 265223 110878
rect 282821 110875 282887 110878
rect 231485 110802 231551 110805
rect 228968 110800 231551 110802
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 213913 110530 213979 110533
rect 217182 110530 217242 110772
rect 228968 110744 231490 110800
rect 231546 110744 231551 110800
rect 228968 110742 231551 110744
rect 231485 110739 231551 110742
rect 213913 110528 217242 110530
rect 213913 110472 213918 110528
rect 213974 110472 217242 110528
rect 213913 110470 217242 110472
rect 265801 110530 265867 110533
rect 268334 110530 268394 110772
rect 265801 110528 268394 110530
rect 265801 110472 265806 110528
rect 265862 110472 268394 110528
rect 265801 110470 268394 110472
rect 213913 110467 213979 110470
rect 265801 110467 265867 110470
rect 231761 110394 231827 110397
rect 228968 110392 231827 110394
rect 228968 110336 231766 110392
rect 231822 110336 231827 110392
rect 228968 110334 231827 110336
rect 231761 110331 231827 110334
rect 167545 110122 167611 110125
rect 164694 110120 167611 110122
rect 164694 110064 167550 110120
rect 167606 110064 167611 110120
rect 164694 110062 167611 110064
rect 167545 110059 167611 110062
rect 214005 109714 214071 109717
rect 217182 109714 217242 110228
rect 265893 110122 265959 110125
rect 268150 110122 268210 110364
rect 282269 110122 282335 110125
rect 265893 110120 268210 110122
rect 265893 110064 265898 110120
rect 265954 110064 268210 110120
rect 265893 110062 268210 110064
rect 279956 110120 282335 110122
rect 279956 110064 282274 110120
rect 282330 110064 282335 110120
rect 279956 110062 282335 110064
rect 265893 110059 265959 110062
rect 282269 110059 282335 110062
rect 230933 109850 230999 109853
rect 228968 109848 230999 109850
rect 228968 109792 230938 109848
rect 230994 109792 230999 109848
rect 228968 109790 230999 109792
rect 230933 109787 230999 109790
rect 214005 109712 217242 109714
rect 214005 109656 214010 109712
rect 214066 109656 217242 109712
rect 214005 109654 217242 109656
rect 265801 109714 265867 109717
rect 268150 109714 268210 109956
rect 265801 109712 268210 109714
rect 265801 109656 265806 109712
rect 265862 109656 268210 109712
rect 265801 109654 268210 109656
rect 214005 109651 214071 109654
rect 265801 109651 265867 109654
rect 213913 109170 213979 109173
rect 217182 109170 217242 109548
rect 231761 109442 231827 109445
rect 228968 109440 231827 109442
rect 228968 109384 231766 109440
rect 231822 109384 231827 109440
rect 228968 109382 231827 109384
rect 231761 109379 231827 109382
rect 265341 109306 265407 109309
rect 268150 109306 268210 109548
rect 282821 109442 282887 109445
rect 279956 109440 282887 109442
rect 279956 109384 282826 109440
rect 282882 109384 282887 109440
rect 279956 109382 282887 109384
rect 282821 109379 282887 109382
rect 265341 109304 268210 109306
rect 265341 109248 265346 109304
rect 265402 109248 268210 109304
rect 265341 109246 268210 109248
rect 265341 109243 265407 109246
rect 213913 109168 217242 109170
rect 213913 109112 213918 109168
rect 213974 109112 217242 109168
rect 213913 109110 217242 109112
rect 213913 109107 213979 109110
rect 231669 108898 231735 108901
rect 228968 108896 231735 108898
rect 167545 108762 167611 108765
rect 164694 108760 167611 108762
rect 164694 108704 167550 108760
rect 167606 108704 167611 108760
rect 164694 108702 167611 108704
rect 167545 108699 167611 108702
rect 213913 108354 213979 108357
rect 217182 108354 217242 108868
rect 228968 108840 231674 108896
rect 231730 108840 231735 108896
rect 228968 108838 231735 108840
rect 231669 108835 231735 108838
rect 264605 108762 264671 108765
rect 268150 108762 268210 109004
rect 264605 108760 268210 108762
rect 264605 108704 264610 108760
rect 264666 108704 268210 108760
rect 264605 108702 268210 108704
rect 264605 108699 264671 108702
rect 281533 108626 281599 108629
rect 279956 108624 281599 108626
rect 231761 108490 231827 108493
rect 228968 108488 231827 108490
rect 228968 108432 231766 108488
rect 231822 108432 231827 108488
rect 228968 108430 231827 108432
rect 231761 108427 231827 108430
rect 213913 108352 217242 108354
rect 213913 108296 213918 108352
rect 213974 108296 217242 108352
rect 213913 108294 217242 108296
rect 265525 108354 265591 108357
rect 268150 108354 268210 108596
rect 279956 108568 281538 108624
rect 281594 108568 281599 108624
rect 279956 108566 281599 108568
rect 281533 108563 281599 108566
rect 265525 108352 268210 108354
rect 265525 108296 265530 108352
rect 265586 108296 268210 108352
rect 265525 108294 268210 108296
rect 213913 108291 213979 108294
rect 265525 108291 265591 108294
rect 214925 107674 214991 107677
rect 217182 107674 217242 108188
rect 231025 107946 231091 107949
rect 228968 107944 231091 107946
rect 228968 107888 231030 107944
rect 231086 107888 231091 107944
rect 228968 107886 231091 107888
rect 231025 107883 231091 107886
rect 265801 107946 265867 107949
rect 268150 107946 268210 108188
rect 265801 107944 268210 107946
rect 265801 107888 265806 107944
rect 265862 107888 268210 107944
rect 265801 107886 268210 107888
rect 265801 107883 265867 107886
rect 282361 107810 282427 107813
rect 279956 107808 282427 107810
rect 214925 107672 217242 107674
rect 214925 107616 214930 107672
rect 214986 107616 217242 107672
rect 214925 107614 217242 107616
rect 265801 107674 265867 107677
rect 265801 107672 267842 107674
rect 265801 107616 265806 107672
rect 265862 107616 267842 107672
rect 265801 107614 267842 107616
rect 214925 107611 214991 107614
rect 265801 107611 265867 107614
rect 231761 107538 231827 107541
rect 228968 107536 231827 107538
rect 214005 106994 214071 106997
rect 217182 106994 217242 107508
rect 228968 107480 231766 107536
rect 231822 107480 231827 107536
rect 228968 107478 231827 107480
rect 267782 107538 267842 107614
rect 268334 107538 268394 107780
rect 279956 107752 282366 107808
rect 282422 107752 282427 107808
rect 279956 107750 282427 107752
rect 282361 107747 282427 107750
rect 267782 107478 268394 107538
rect 231761 107475 231827 107478
rect 231485 107130 231551 107133
rect 228968 107128 231551 107130
rect 228968 107072 231490 107128
rect 231546 107072 231551 107128
rect 228968 107070 231551 107072
rect 231485 107067 231551 107070
rect 265433 107130 265499 107133
rect 268150 107130 268210 107372
rect 281717 107130 281783 107133
rect 265433 107128 268210 107130
rect 265433 107072 265438 107128
rect 265494 107072 268210 107128
rect 265433 107070 268210 107072
rect 279956 107128 281783 107130
rect 279956 107072 281722 107128
rect 281778 107072 281783 107128
rect 279956 107070 281783 107072
rect 265433 107067 265499 107070
rect 281717 107067 281783 107070
rect 214005 106992 217242 106994
rect 214005 106936 214010 106992
rect 214066 106936 217242 106992
rect 214005 106934 217242 106936
rect 214005 106931 214071 106934
rect 213913 106586 213979 106589
rect 217182 106586 217242 106828
rect 265801 106722 265867 106725
rect 268150 106722 268210 106964
rect 265801 106720 268210 106722
rect 265801 106664 265806 106720
rect 265862 106664 268210 106720
rect 265801 106662 268210 106664
rect 265801 106659 265867 106662
rect 231209 106586 231275 106589
rect 213913 106584 217242 106586
rect 213913 106528 213918 106584
rect 213974 106528 217242 106584
rect 213913 106526 217242 106528
rect 228968 106584 231275 106586
rect 228968 106528 231214 106584
rect 231270 106528 231275 106584
rect 228968 106526 231275 106528
rect 213913 106523 213979 106526
rect 231209 106523 231275 106526
rect 265893 106586 265959 106589
rect 265893 106584 268210 106586
rect 265893 106528 265898 106584
rect 265954 106528 268210 106584
rect 265893 106526 268210 106528
rect 265893 106523 265959 106526
rect 268150 106420 268210 106526
rect 280245 106314 280311 106317
rect 279956 106312 280311 106314
rect 279956 106256 280250 106312
rect 280306 106256 280311 106312
rect 279956 106254 280311 106256
rect 280245 106251 280311 106254
rect 231761 106178 231827 106181
rect 228968 106176 231827 106178
rect 214097 105770 214163 105773
rect 217182 105770 217242 106148
rect 228968 106120 231766 106176
rect 231822 106120 231827 106176
rect 228968 106118 231827 106120
rect 231761 106115 231827 106118
rect 214097 105768 217242 105770
rect 214097 105712 214102 105768
rect 214158 105712 217242 105768
rect 214097 105710 217242 105712
rect 265801 105770 265867 105773
rect 268150 105770 268210 106012
rect 265801 105768 268210 105770
rect 265801 105712 265806 105768
rect 265862 105712 268210 105768
rect 265801 105710 268210 105712
rect 214097 105707 214163 105710
rect 265801 105707 265867 105710
rect 230749 105634 230815 105637
rect 228968 105632 230815 105634
rect 214005 105362 214071 105365
rect 217182 105362 217242 105604
rect 228968 105576 230754 105632
rect 230810 105576 230815 105632
rect 228968 105574 230815 105576
rect 230749 105571 230815 105574
rect 214005 105360 217242 105362
rect 214005 105304 214010 105360
rect 214066 105304 217242 105360
rect 214005 105302 217242 105304
rect 265433 105362 265499 105365
rect 268150 105362 268210 105604
rect 282821 105498 282887 105501
rect 279956 105496 282887 105498
rect 279956 105440 282826 105496
rect 282882 105440 282887 105496
rect 279956 105438 282887 105440
rect 282821 105435 282887 105438
rect 265433 105360 268210 105362
rect 265433 105304 265438 105360
rect 265494 105304 268210 105360
rect 265433 105302 268210 105304
rect 214005 105299 214071 105302
rect 265433 105299 265499 105302
rect 231669 105226 231735 105229
rect 228968 105224 231735 105226
rect 228968 105168 231674 105224
rect 231730 105168 231735 105224
rect 228968 105166 231735 105168
rect 231669 105163 231735 105166
rect 213913 105090 213979 105093
rect 213913 105088 217242 105090
rect 213913 105032 213918 105088
rect 213974 105032 217242 105088
rect 213913 105030 217242 105032
rect 213913 105027 213979 105030
rect 217182 104924 217242 105030
rect 264789 104954 264855 104957
rect 268150 104954 268210 105196
rect 264789 104952 268210 104954
rect 264789 104896 264794 104952
rect 264850 104896 268210 104952
rect 264789 104894 268210 104896
rect 264789 104891 264855 104894
rect 281533 104818 281599 104821
rect 279956 104816 281599 104818
rect 230749 104682 230815 104685
rect 228968 104680 230815 104682
rect 228968 104624 230754 104680
rect 230810 104624 230815 104680
rect 228968 104622 230815 104624
rect 230749 104619 230815 104622
rect 265341 104546 265407 104549
rect 268150 104546 268210 104788
rect 279956 104760 281538 104816
rect 281594 104760 281599 104816
rect 279956 104758 281599 104760
rect 281533 104755 281599 104758
rect 265341 104544 268210 104546
rect 265341 104488 265346 104544
rect 265402 104488 268210 104544
rect 265341 104486 268210 104488
rect 265341 104483 265407 104486
rect 230933 104274 230999 104277
rect 228968 104272 230999 104274
rect 213913 103730 213979 103733
rect 217182 103730 217242 104244
rect 228968 104216 230938 104272
rect 230994 104216 230999 104272
rect 228968 104214 230999 104216
rect 230933 104211 230999 104214
rect 265157 104002 265223 104005
rect 268150 104002 268210 104380
rect 281533 104002 281599 104005
rect 265157 104000 268210 104002
rect 265157 103944 265162 104000
rect 265218 103944 268210 104000
rect 265157 103942 268210 103944
rect 279956 104000 281599 104002
rect 279956 103944 281538 104000
rect 281594 103944 281599 104000
rect 279956 103942 281599 103944
rect 265157 103939 265223 103942
rect 281533 103939 281599 103942
rect 231761 103730 231827 103733
rect 213913 103728 217242 103730
rect 213913 103672 213918 103728
rect 213974 103672 217242 103728
rect 213913 103670 217242 103672
rect 228968 103728 231827 103730
rect 228968 103672 231766 103728
rect 231822 103672 231827 103728
rect 228968 103670 231827 103672
rect 213913 103667 213979 103670
rect 231761 103667 231827 103670
rect 214414 103532 214420 103596
rect 214484 103594 214490 103596
rect 265801 103594 265867 103597
rect 268334 103594 268394 103836
rect 214484 103534 217058 103594
rect 265801 103592 268394 103594
rect 214484 103532 214490 103534
rect 216998 103530 217058 103534
rect 217182 103530 217242 103564
rect 265801 103536 265806 103592
rect 265862 103536 268394 103592
rect 265801 103534 268394 103536
rect 265801 103531 265867 103534
rect 216998 103470 217242 103530
rect 231761 103322 231827 103325
rect 228968 103320 231827 103322
rect 228968 103264 231766 103320
rect 231822 103264 231827 103320
rect 228968 103262 231827 103264
rect 231761 103259 231827 103262
rect 264697 103186 264763 103189
rect 268150 103186 268210 103428
rect 282821 103186 282887 103189
rect 264697 103184 268210 103186
rect 264697 103128 264702 103184
rect 264758 103128 268210 103184
rect 264697 103126 268210 103128
rect 279956 103184 282887 103186
rect 279956 103128 282826 103184
rect 282882 103128 282887 103184
rect 279956 103126 282887 103128
rect 264697 103123 264763 103126
rect 282821 103123 282887 103126
rect 214005 102642 214071 102645
rect 217182 102642 217242 102884
rect 230565 102778 230631 102781
rect 228968 102776 230631 102778
rect 228968 102720 230570 102776
rect 230626 102720 230631 102776
rect 228968 102718 230631 102720
rect 230565 102715 230631 102718
rect 265433 102778 265499 102781
rect 268150 102778 268210 103020
rect 265433 102776 268210 102778
rect 265433 102720 265438 102776
rect 265494 102720 268210 102776
rect 265433 102718 268210 102720
rect 265433 102715 265499 102718
rect 214005 102640 217242 102642
rect 214005 102584 214010 102640
rect 214066 102584 217242 102640
rect 214005 102582 217242 102584
rect 214005 102579 214071 102582
rect 65977 102370 66043 102373
rect 68142 102370 68816 102376
rect 65977 102368 68816 102370
rect 65977 102312 65982 102368
rect 66038 102316 68816 102368
rect 213913 102370 213979 102373
rect 231485 102370 231551 102373
rect 213913 102368 217242 102370
rect 66038 102312 68202 102316
rect 65977 102310 68202 102312
rect 213913 102312 213918 102368
rect 213974 102312 217242 102368
rect 213913 102310 217242 102312
rect 228968 102368 231551 102370
rect 228968 102312 231490 102368
rect 231546 102312 231551 102368
rect 228968 102310 231551 102312
rect 65977 102307 66043 102310
rect 213913 102307 213979 102310
rect 217182 102204 217242 102310
rect 231485 102307 231551 102310
rect 265801 102370 265867 102373
rect 268518 102372 268578 102612
rect 281993 102506 282059 102509
rect 279956 102504 282059 102506
rect 279956 102448 281998 102504
rect 282054 102448 282059 102504
rect 279956 102446 282059 102448
rect 281993 102443 282059 102446
rect 265801 102368 268210 102370
rect 265801 102312 265806 102368
rect 265862 102312 268210 102368
rect 265801 102310 268210 102312
rect 265801 102307 265867 102310
rect 268150 102204 268210 102310
rect 268510 102308 268516 102372
rect 268580 102308 268586 102372
rect 230657 101826 230723 101829
rect 228968 101824 230723 101826
rect 228968 101768 230662 101824
rect 230718 101768 230723 101824
rect 228968 101766 230723 101768
rect 230657 101763 230723 101766
rect 213862 101084 213868 101148
rect 213932 101146 213938 101148
rect 217182 101146 217242 101524
rect 231761 101418 231827 101421
rect 228968 101416 231827 101418
rect 228968 101360 231766 101416
rect 231822 101360 231827 101416
rect 228968 101358 231827 101360
rect 231761 101355 231827 101358
rect 265893 101418 265959 101421
rect 268150 101418 268210 101796
rect 281625 101690 281691 101693
rect 279956 101688 281691 101690
rect 279956 101632 281630 101688
rect 281686 101632 281691 101688
rect 279956 101630 281691 101632
rect 281625 101627 281691 101630
rect 265893 101416 268210 101418
rect 265893 101360 265898 101416
rect 265954 101360 268210 101416
rect 265893 101358 268210 101360
rect 265893 101355 265959 101358
rect 213932 101086 217242 101146
rect 213932 101084 213938 101086
rect 265525 101010 265591 101013
rect 268150 101010 268210 101252
rect 265525 101008 268210 101010
rect 214373 100874 214439 100877
rect 214373 100872 216874 100874
rect 214373 100816 214378 100872
rect 214434 100816 216874 100872
rect 214373 100814 216874 100816
rect 214373 100811 214439 100814
rect 66161 100738 66227 100741
rect 68142 100738 68816 100744
rect 66161 100736 68816 100738
rect 66161 100680 66166 100736
rect 66222 100684 68816 100736
rect 216814 100738 216874 100814
rect 217366 100738 217426 100980
rect 265525 100952 265530 101008
rect 265586 100952 268210 101008
rect 265525 100950 268210 100952
rect 265525 100947 265591 100950
rect 231117 100874 231183 100877
rect 228968 100872 231183 100874
rect 228968 100816 231122 100872
rect 231178 100816 231183 100872
rect 228968 100814 231183 100816
rect 231117 100811 231183 100814
rect 265801 100874 265867 100877
rect 280286 100874 280292 100876
rect 265801 100872 268026 100874
rect 265801 100816 265806 100872
rect 265862 100840 268026 100872
rect 268150 100840 268210 100844
rect 265862 100816 268210 100840
rect 265801 100814 268210 100816
rect 279956 100814 280292 100874
rect 265801 100811 265867 100814
rect 267966 100780 268210 100814
rect 280286 100812 280292 100814
rect 280356 100812 280362 100876
rect 66222 100680 68202 100684
rect 66161 100678 68202 100680
rect 216814 100678 217426 100738
rect 66161 100675 66227 100678
rect 261661 100602 261727 100605
rect 268510 100602 268516 100604
rect 261661 100600 268516 100602
rect 261661 100544 261666 100600
rect 261722 100544 268516 100600
rect 261661 100542 268516 100544
rect 261661 100539 261727 100542
rect 268510 100540 268516 100542
rect 268580 100540 268586 100604
rect 231669 100466 231735 100469
rect 228968 100464 231735 100466
rect 228968 100408 231674 100464
rect 231730 100408 231735 100464
rect 228968 100406 231735 100408
rect 231669 100403 231735 100406
rect 214189 99786 214255 99789
rect 217182 99786 217242 100300
rect 265893 100194 265959 100197
rect 268150 100194 268210 100436
rect 282269 100194 282335 100197
rect 265893 100192 268210 100194
rect 265893 100136 265898 100192
rect 265954 100136 268210 100192
rect 265893 100134 268210 100136
rect 279956 100192 282335 100194
rect 279956 100136 282274 100192
rect 282330 100136 282335 100192
rect 279956 100134 282335 100136
rect 265893 100131 265959 100134
rect 282269 100131 282335 100134
rect 231761 99922 231827 99925
rect 228968 99920 231827 99922
rect 228968 99864 231766 99920
rect 231822 99864 231827 99920
rect 228968 99862 231827 99864
rect 231761 99859 231827 99862
rect 214189 99784 217242 99786
rect 214189 99728 214194 99784
rect 214250 99728 217242 99784
rect 214189 99726 217242 99728
rect 265801 99786 265867 99789
rect 268150 99786 268210 100028
rect 265801 99784 268210 99786
rect 265801 99728 265806 99784
rect 265862 99728 268210 99784
rect 265801 99726 268210 99728
rect 214189 99723 214255 99726
rect 265801 99723 265867 99726
rect 214097 99514 214163 99517
rect 214097 99512 216874 99514
rect 214097 99456 214102 99512
rect 214158 99456 216874 99512
rect 214097 99454 216874 99456
rect 214097 99451 214163 99454
rect 216814 99378 216874 99454
rect 217366 99378 217426 99620
rect 230841 99514 230907 99517
rect 228968 99512 230907 99514
rect 228968 99456 230846 99512
rect 230902 99456 230907 99512
rect 228968 99454 230907 99456
rect 230841 99451 230907 99454
rect 265525 99514 265591 99517
rect 265525 99512 267842 99514
rect 265525 99456 265530 99512
rect 265586 99456 267842 99512
rect 265525 99454 267842 99456
rect 265525 99451 265591 99454
rect 216814 99318 217426 99378
rect 267782 99378 267842 99454
rect 268334 99378 268394 99620
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 281533 99378 281599 99381
rect 267782 99318 268394 99378
rect 279956 99376 281599 99378
rect 279956 99320 281538 99376
rect 281594 99320 281599 99376
rect 583520 99364 584960 99454
rect 279956 99318 281599 99320
rect 281533 99315 281599 99318
rect 231025 98970 231091 98973
rect 228968 98968 231091 98970
rect 213913 98426 213979 98429
rect 217182 98426 217242 98940
rect 228968 98912 231030 98968
rect 231086 98912 231091 98968
rect 228968 98910 231091 98912
rect 231025 98907 231091 98910
rect 265709 98834 265775 98837
rect 268150 98834 268210 99212
rect 265709 98832 268210 98834
rect 265709 98776 265714 98832
rect 265770 98776 268210 98832
rect 265709 98774 268210 98776
rect 265709 98771 265775 98774
rect 231301 98562 231367 98565
rect 228968 98560 231367 98562
rect 228968 98504 231306 98560
rect 231362 98504 231367 98560
rect 228968 98502 231367 98504
rect 231301 98499 231367 98502
rect 213913 98424 217242 98426
rect 213913 98368 213918 98424
rect 213974 98368 217242 98424
rect 213913 98366 217242 98368
rect 265985 98426 266051 98429
rect 268150 98426 268210 98668
rect 265985 98424 268210 98426
rect 265985 98368 265990 98424
rect 266046 98368 268210 98424
rect 265985 98366 268210 98368
rect 213913 98363 213979 98366
rect 265985 98363 266051 98366
rect 214005 98018 214071 98021
rect 217182 98018 217242 98260
rect 230749 98018 230815 98021
rect 214005 98016 217242 98018
rect 214005 97960 214010 98016
rect 214066 97960 217242 98016
rect 214005 97958 217242 97960
rect 228968 98016 230815 98018
rect 228968 97960 230754 98016
rect 230810 97960 230815 98016
rect 228968 97958 230815 97960
rect 214005 97955 214071 97958
rect 230749 97955 230815 97958
rect 265801 98018 265867 98021
rect 268334 98018 268394 98260
rect 279374 98157 279434 98532
rect 279374 98152 279483 98157
rect 279374 98096 279422 98152
rect 279478 98096 279483 98152
rect 279374 98094 279483 98096
rect 279417 98091 279483 98094
rect 265801 98016 268394 98018
rect 265801 97960 265806 98016
rect 265862 97960 268394 98016
rect 265801 97958 268394 97960
rect 265801 97955 265867 97958
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect 231577 97610 231643 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect 228968 97608 231643 97610
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 213913 97066 213979 97069
rect 217182 97066 217242 97580
rect 228968 97552 231582 97608
rect 231638 97552 231643 97608
rect 228968 97550 231643 97552
rect 231577 97547 231643 97550
rect 265893 97610 265959 97613
rect 268150 97610 268210 97852
rect 265893 97608 268210 97610
rect 265893 97552 265898 97608
rect 265954 97552 268210 97608
rect 265893 97550 268210 97552
rect 265893 97547 265959 97550
rect 265617 97202 265683 97205
rect 268150 97202 268210 97444
rect 279558 97341 279618 97852
rect 279509 97336 279618 97341
rect 279509 97280 279514 97336
rect 279570 97280 279618 97336
rect 279509 97278 279618 97280
rect 279509 97275 279575 97278
rect 265617 97200 268210 97202
rect 265617 97144 265622 97200
rect 265678 97144 268210 97200
rect 265617 97142 268210 97144
rect 265617 97139 265683 97142
rect 268326 97140 268332 97204
rect 268396 97140 268402 97204
rect 230749 97066 230815 97069
rect 231761 97066 231827 97069
rect 213913 97064 217242 97066
rect 213913 97008 213918 97064
rect 213974 97008 217242 97064
rect 213913 97006 217242 97008
rect 228968 97064 231827 97066
rect 228968 97008 230754 97064
rect 230810 97008 231766 97064
rect 231822 97008 231827 97064
rect 268334 97036 268394 97140
rect 228968 97006 231827 97008
rect 213913 97003 213979 97006
rect 230749 97003 230815 97006
rect 231761 97003 231827 97006
rect 265801 96930 265867 96933
rect 267774 96930 267780 96932
rect 265801 96928 267780 96930
rect 166390 96596 166396 96660
rect 166460 96658 166466 96660
rect 217182 96658 217242 96900
rect 265801 96872 265806 96928
rect 265862 96872 267780 96928
rect 265801 96870 267780 96872
rect 265801 96867 265867 96870
rect 267774 96868 267780 96870
rect 267844 96868 267850 96932
rect 265525 96794 265591 96797
rect 265525 96792 268210 96794
rect 265525 96736 265530 96792
rect 265586 96736 268210 96792
rect 265525 96734 268210 96736
rect 265525 96731 265591 96734
rect 230657 96658 230723 96661
rect 231301 96658 231367 96661
rect 166460 96598 217242 96658
rect 228968 96656 231367 96658
rect 228968 96600 230662 96656
rect 230718 96600 231306 96656
rect 231362 96600 231367 96656
rect 268150 96628 268210 96734
rect 279374 96661 279434 97036
rect 279325 96656 279434 96661
rect 228968 96598 231367 96600
rect 166460 96596 166466 96598
rect 230657 96595 230723 96598
rect 231301 96595 231367 96598
rect 279325 96600 279330 96656
rect 279386 96600 279434 96656
rect 279325 96598 279434 96600
rect 279325 96595 279391 96598
rect 213913 95842 213979 95845
rect 217182 95842 217242 96356
rect 213913 95840 217242 95842
rect 213913 95784 213918 95840
rect 213974 95784 217242 95840
rect 213913 95782 217242 95784
rect 228774 95842 228834 96220
rect 230565 95842 230631 95845
rect 228774 95840 230631 95842
rect 228774 95784 230570 95840
rect 230626 95784 230631 95840
rect 228774 95782 230631 95784
rect 213913 95779 213979 95782
rect 230565 95779 230631 95782
rect 265709 95706 265775 95709
rect 268150 95706 268210 96220
rect 279233 96114 279299 96117
rect 279374 96114 279434 96356
rect 279233 96112 279434 96114
rect 279233 96056 279238 96112
rect 279294 96056 279434 96112
rect 279233 96054 279434 96056
rect 279233 96051 279299 96054
rect 265709 95704 268210 95706
rect 265709 95648 265714 95704
rect 265770 95648 268210 95704
rect 265709 95646 268210 95648
rect 265709 95643 265775 95646
rect 67817 94890 67883 94893
rect 213862 94890 213868 94892
rect 67817 94888 213868 94890
rect 67817 94832 67822 94888
rect 67878 94832 213868 94888
rect 67817 94830 213868 94832
rect 67817 94827 67883 94830
rect 213862 94828 213868 94830
rect 213932 94828 213938 94892
rect 67633 94754 67699 94757
rect 214414 94754 214420 94756
rect 67633 94752 214420 94754
rect 67633 94696 67638 94752
rect 67694 94696 214420 94752
rect 67633 94694 214420 94696
rect 67633 94691 67699 94694
rect 214414 94692 214420 94694
rect 214484 94692 214490 94756
rect 66161 94618 66227 94621
rect 166390 94618 166396 94620
rect 66161 94616 166396 94618
rect 66161 94560 66166 94616
rect 66222 94560 166396 94616
rect 66161 94558 166396 94560
rect 66161 94555 66227 94558
rect 166390 94556 166396 94558
rect 166460 94556 166466 94620
rect 65977 94482 66043 94485
rect 165521 94482 165587 94485
rect 65977 94480 165587 94482
rect 65977 94424 65982 94480
rect 66038 94424 165526 94480
rect 165582 94424 165587 94480
rect 65977 94422 165587 94424
rect 65977 94419 66043 94422
rect 165521 94419 165587 94422
rect 151629 94348 151695 94349
rect 151624 94346 151630 94348
rect 151538 94286 151630 94346
rect 151624 94284 151630 94286
rect 151694 94284 151700 94348
rect 151629 94283 151695 94284
rect 124121 94212 124187 94213
rect 124070 94148 124076 94212
rect 124140 94210 124187 94212
rect 124140 94208 124232 94210
rect 124182 94152 124232 94208
rect 124140 94150 124232 94152
rect 124140 94148 124187 94150
rect 124121 94147 124187 94148
rect 117129 94076 117195 94077
rect 122097 94076 122163 94077
rect 151721 94076 151787 94077
rect 117078 94012 117084 94076
rect 117148 94074 117195 94076
rect 117148 94072 117240 94074
rect 117190 94016 117240 94072
rect 117148 94014 117240 94016
rect 117148 94012 117195 94014
rect 122046 94012 122052 94076
rect 122116 94074 122163 94076
rect 122116 94072 122208 94074
rect 122158 94016 122208 94072
rect 122116 94014 122208 94016
rect 122116 94012 122163 94014
rect 151670 94012 151676 94076
rect 151740 94074 151787 94076
rect 151740 94072 151832 94074
rect 151782 94016 151832 94072
rect 151740 94014 151832 94016
rect 151740 94012 151787 94014
rect 117129 94011 117195 94012
rect 122097 94011 122163 94012
rect 151721 94011 151787 94012
rect 118233 93940 118299 93941
rect 151537 93940 151603 93941
rect 118182 93876 118188 93940
rect 118252 93938 118299 93940
rect 118252 93936 118344 93938
rect 118294 93880 118344 93936
rect 118252 93878 118344 93880
rect 118252 93876 118299 93878
rect 151486 93876 151492 93940
rect 151556 93938 151603 93940
rect 151556 93936 151648 93938
rect 151598 93880 151648 93936
rect 151556 93878 151648 93880
rect 151556 93876 151603 93878
rect 118233 93875 118299 93876
rect 151537 93875 151603 93876
rect 100886 93740 100892 93804
rect 100956 93802 100962 93804
rect 169017 93802 169083 93805
rect 100956 93800 169083 93802
rect 100956 93744 169022 93800
rect 169078 93744 169083 93800
rect 100956 93742 169083 93744
rect 100956 93740 100962 93742
rect 169017 93739 169083 93742
rect 102961 93668 103027 93669
rect 104249 93668 104315 93669
rect 105537 93668 105603 93669
rect 106457 93668 106523 93669
rect 107745 93668 107811 93669
rect 109217 93668 109283 93669
rect 119705 93668 119771 93669
rect 102910 93666 102916 93668
rect 102870 93606 102916 93666
rect 102980 93664 103027 93668
rect 104198 93666 104204 93668
rect 103022 93608 103027 93664
rect 102910 93604 102916 93606
rect 102980 93604 103027 93608
rect 104158 93606 104204 93666
rect 104268 93664 104315 93668
rect 105486 93666 105492 93668
rect 104310 93608 104315 93664
rect 104198 93604 104204 93606
rect 104268 93604 104315 93608
rect 105446 93606 105492 93666
rect 105556 93664 105603 93668
rect 106406 93666 106412 93668
rect 105598 93608 105603 93664
rect 105486 93604 105492 93606
rect 105556 93604 105603 93608
rect 106366 93606 106412 93666
rect 106476 93664 106523 93668
rect 107694 93666 107700 93668
rect 106518 93608 106523 93664
rect 106406 93604 106412 93606
rect 106476 93604 106523 93608
rect 107654 93606 107700 93666
rect 107764 93664 107811 93668
rect 109166 93666 109172 93668
rect 107806 93608 107811 93664
rect 107694 93604 107700 93606
rect 107764 93604 107811 93608
rect 109126 93606 109172 93666
rect 109236 93664 109283 93668
rect 119654 93666 119660 93668
rect 109278 93608 109283 93664
rect 109166 93604 109172 93606
rect 109236 93604 109283 93608
rect 119614 93606 119660 93666
rect 119724 93664 119771 93668
rect 164918 93666 164924 93668
rect 119766 93608 119771 93664
rect 119654 93604 119660 93606
rect 119724 93604 119771 93608
rect 102961 93603 103027 93604
rect 104249 93603 104315 93604
rect 105537 93603 105603 93604
rect 106457 93603 106523 93604
rect 107745 93603 107811 93604
rect 109217 93603 109283 93604
rect 119705 93603 119771 93604
rect 122790 93606 164924 93666
rect 90265 93532 90331 93533
rect 101857 93532 101923 93533
rect 90214 93530 90220 93532
rect 90174 93470 90220 93530
rect 90284 93528 90331 93532
rect 101806 93530 101812 93532
rect 90326 93472 90331 93528
rect 90214 93468 90220 93470
rect 90284 93468 90331 93472
rect 101766 93470 101812 93530
rect 101876 93528 101923 93532
rect 101918 93472 101923 93528
rect 101806 93468 101812 93470
rect 101876 93468 101923 93472
rect 111374 93468 111380 93532
rect 111444 93530 111450 93532
rect 111793 93530 111859 93533
rect 111444 93528 111859 93530
rect 111444 93472 111798 93528
rect 111854 93472 111859 93528
rect 111444 93470 111859 93472
rect 111444 93468 111450 93470
rect 90265 93467 90331 93468
rect 101857 93467 101923 93468
rect 111793 93467 111859 93470
rect 119286 93468 119292 93532
rect 119356 93530 119362 93532
rect 122790 93530 122850 93606
rect 164918 93604 164924 93606
rect 164988 93604 164994 93668
rect 125409 93532 125475 93533
rect 125358 93530 125364 93532
rect 119356 93470 122850 93530
rect 125318 93470 125364 93530
rect 125428 93528 125475 93532
rect 125470 93472 125475 93528
rect 119356 93468 119362 93470
rect 125358 93468 125364 93470
rect 125428 93468 125475 93472
rect 125409 93467 125475 93468
rect 135713 93396 135779 93397
rect 135662 93394 135668 93396
rect 135622 93334 135668 93394
rect 135732 93392 135779 93396
rect 135774 93336 135779 93392
rect 135662 93332 135668 93334
rect 135732 93332 135779 93336
rect 135713 93331 135779 93332
rect 110137 93260 110203 93261
rect 128169 93260 128235 93261
rect 110086 93258 110092 93260
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 128118 93258 128124 93260
rect 110198 93200 110203 93256
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 128078 93198 128124 93258
rect 128188 93256 128235 93260
rect 128230 93200 128235 93256
rect 128118 93196 128124 93198
rect 128188 93196 128235 93200
rect 110137 93195 110203 93196
rect 128169 93195 128235 93196
rect 126053 93122 126119 93125
rect 214741 93122 214807 93125
rect 126053 93120 214807 93122
rect 126053 93064 126058 93120
rect 126114 93064 214746 93120
rect 214802 93064 214807 93120
rect 126053 93062 214807 93064
rect 126053 93059 126119 93062
rect 214741 93059 214807 93062
rect 113030 92516 113036 92580
rect 113100 92578 113106 92580
rect 113173 92578 113239 92581
rect 113100 92576 113239 92578
rect 113100 92520 113178 92576
rect 113234 92520 113239 92576
rect 113100 92518 113239 92520
rect 113100 92516 113106 92518
rect 113173 92515 113239 92518
rect 84377 92444 84443 92445
rect 84326 92442 84332 92444
rect 84286 92382 84332 92442
rect 84396 92440 84443 92444
rect 84438 92384 84443 92440
rect 84326 92380 84332 92382
rect 84396 92380 84443 92384
rect 85798 92380 85804 92444
rect 85868 92442 85874 92444
rect 86677 92442 86743 92445
rect 88057 92444 88123 92445
rect 88006 92442 88012 92444
rect 85868 92440 86743 92442
rect 85868 92384 86682 92440
rect 86738 92384 86743 92440
rect 85868 92382 86743 92384
rect 87966 92382 88012 92442
rect 88076 92440 88123 92444
rect 88118 92384 88123 92440
rect 85868 92380 85874 92382
rect 84377 92379 84443 92380
rect 86677 92379 86743 92382
rect 88006 92380 88012 92382
rect 88076 92380 88123 92384
rect 88926 92380 88932 92444
rect 88996 92442 89002 92444
rect 89069 92442 89135 92445
rect 88996 92440 89135 92442
rect 88996 92384 89074 92440
rect 89130 92384 89135 92440
rect 88996 92382 89135 92384
rect 88996 92380 89002 92382
rect 88057 92379 88123 92380
rect 89069 92379 89135 92382
rect 91318 92380 91324 92444
rect 91388 92442 91394 92444
rect 91461 92442 91527 92445
rect 91388 92440 91527 92442
rect 91388 92384 91466 92440
rect 91522 92384 91527 92440
rect 91388 92382 91527 92384
rect 91388 92380 91394 92382
rect 91461 92379 91527 92382
rect 93894 92380 93900 92444
rect 93964 92442 93970 92444
rect 94957 92442 95023 92445
rect 100017 92444 100083 92445
rect 105721 92444 105787 92445
rect 108113 92444 108179 92445
rect 99966 92442 99972 92444
rect 93964 92440 95023 92442
rect 93964 92384 94962 92440
rect 95018 92384 95023 92440
rect 93964 92382 95023 92384
rect 99926 92382 99972 92442
rect 100036 92440 100083 92444
rect 105670 92442 105676 92444
rect 100078 92384 100083 92440
rect 93964 92380 93970 92382
rect 94957 92379 95023 92382
rect 99966 92380 99972 92382
rect 100036 92380 100083 92384
rect 105630 92382 105676 92442
rect 105740 92440 105787 92444
rect 108062 92442 108068 92444
rect 105782 92384 105787 92440
rect 105670 92380 105676 92382
rect 105740 92380 105787 92384
rect 108022 92382 108068 92442
rect 108132 92440 108179 92444
rect 108174 92384 108179 92440
rect 108062 92380 108068 92382
rect 108132 92380 108179 92384
rect 109534 92380 109540 92444
rect 109604 92442 109610 92444
rect 109953 92442 110019 92445
rect 109604 92440 110019 92442
rect 109604 92384 109958 92440
rect 110014 92384 110019 92440
rect 109604 92382 110019 92384
rect 109604 92380 109610 92382
rect 100017 92379 100083 92380
rect 105721 92379 105787 92380
rect 108113 92379 108179 92380
rect 109953 92379 110019 92382
rect 110638 92380 110644 92444
rect 110708 92442 110714 92444
rect 110965 92442 111031 92445
rect 111977 92444 112043 92445
rect 112345 92444 112411 92445
rect 111926 92442 111932 92444
rect 110708 92440 111031 92442
rect 110708 92384 110970 92440
rect 111026 92384 111031 92440
rect 110708 92382 111031 92384
rect 111886 92382 111932 92442
rect 111996 92440 112043 92444
rect 112294 92442 112300 92444
rect 112038 92384 112043 92440
rect 110708 92380 110714 92382
rect 110965 92379 111031 92382
rect 111926 92380 111932 92382
rect 111996 92380 112043 92384
rect 112254 92382 112300 92442
rect 112364 92440 112411 92444
rect 112406 92384 112411 92440
rect 112294 92380 112300 92382
rect 112364 92380 112411 92384
rect 113214 92380 113220 92444
rect 113284 92442 113290 92444
rect 113357 92442 113423 92445
rect 114369 92444 114435 92445
rect 114318 92442 114324 92444
rect 113284 92440 113423 92442
rect 113284 92384 113362 92440
rect 113418 92384 113423 92440
rect 113284 92382 113423 92384
rect 114278 92382 114324 92442
rect 114388 92440 114435 92444
rect 114430 92384 114435 92440
rect 113284 92380 113290 92382
rect 111977 92379 112043 92380
rect 112345 92379 112411 92380
rect 113357 92379 113423 92382
rect 114318 92380 114324 92382
rect 114388 92380 114435 92384
rect 114870 92380 114876 92444
rect 114940 92442 114946 92444
rect 115197 92442 115263 92445
rect 115841 92444 115907 92445
rect 118049 92444 118115 92445
rect 120257 92444 120323 92445
rect 115790 92442 115796 92444
rect 114940 92440 115263 92442
rect 114940 92384 115202 92440
rect 115258 92384 115263 92440
rect 114940 92382 115263 92384
rect 115750 92382 115796 92442
rect 115860 92440 115907 92444
rect 117998 92442 118004 92444
rect 115902 92384 115907 92440
rect 114940 92380 114946 92382
rect 114369 92379 114435 92380
rect 115197 92379 115263 92382
rect 115790 92380 115796 92382
rect 115860 92380 115907 92384
rect 117958 92382 118004 92442
rect 118068 92440 118115 92444
rect 120206 92442 120212 92444
rect 118110 92384 118115 92440
rect 117998 92380 118004 92382
rect 118068 92380 118115 92384
rect 120166 92382 120212 92442
rect 120276 92440 120323 92444
rect 120318 92384 120323 92440
rect 120206 92380 120212 92382
rect 120276 92380 120323 92384
rect 120574 92380 120580 92444
rect 120644 92442 120650 92444
rect 121177 92442 121243 92445
rect 125777 92444 125843 92445
rect 129457 92444 129523 92445
rect 132401 92444 132467 92445
rect 134425 92444 134491 92445
rect 125726 92442 125732 92444
rect 120644 92440 121243 92442
rect 120644 92384 121182 92440
rect 121238 92384 121243 92440
rect 120644 92382 121243 92384
rect 125686 92382 125732 92442
rect 125796 92440 125843 92444
rect 129406 92442 129412 92444
rect 125838 92384 125843 92440
rect 120644 92380 120650 92382
rect 115841 92379 115907 92380
rect 118049 92379 118115 92380
rect 120257 92379 120323 92380
rect 121177 92379 121243 92382
rect 125726 92380 125732 92382
rect 125796 92380 125843 92384
rect 129366 92382 129412 92442
rect 129476 92440 129523 92444
rect 132350 92442 132356 92444
rect 129518 92384 129523 92440
rect 129406 92380 129412 92382
rect 129476 92380 129523 92384
rect 132310 92382 132356 92442
rect 132420 92440 132467 92444
rect 134374 92442 134380 92444
rect 132462 92384 132467 92440
rect 132350 92380 132356 92382
rect 132420 92380 132467 92384
rect 134334 92382 134380 92442
rect 134444 92440 134491 92444
rect 134486 92384 134491 92440
rect 134374 92380 134380 92382
rect 134444 92380 134491 92384
rect 152038 92380 152044 92444
rect 152108 92442 152114 92444
rect 153101 92442 153167 92445
rect 152108 92440 153167 92442
rect 152108 92384 153106 92440
rect 153162 92384 153167 92440
rect 152108 92382 153167 92384
rect 152108 92380 152114 92382
rect 125777 92379 125843 92380
rect 129457 92379 129523 92380
rect 132401 92379 132467 92380
rect 134425 92379 134491 92380
rect 153101 92379 153167 92382
rect 98126 92244 98132 92308
rect 98196 92306 98202 92308
rect 167821 92306 167887 92309
rect 98196 92304 167887 92306
rect 98196 92248 167826 92304
rect 167882 92248 167887 92304
rect 98196 92246 167887 92248
rect 98196 92244 98202 92246
rect 167821 92243 167887 92246
rect 103830 92108 103836 92172
rect 103900 92170 103906 92172
rect 171777 92170 171843 92173
rect 103900 92168 171843 92170
rect 103900 92112 171782 92168
rect 171838 92112 171843 92168
rect 103900 92110 171843 92112
rect 103900 92108 103906 92110
rect 171777 92107 171843 92110
rect 106774 91972 106780 92036
rect 106844 92034 106850 92036
rect 169201 92034 169267 92037
rect 106844 92032 169267 92034
rect 106844 91976 169206 92032
rect 169262 91976 169267 92032
rect 106844 91974 169267 91976
rect 106844 91972 106850 91974
rect 169201 91971 169267 91974
rect 121678 91836 121684 91900
rect 121748 91898 121754 91900
rect 121913 91898 121979 91901
rect 121748 91896 121979 91898
rect 121748 91840 121918 91896
rect 121974 91840 121979 91896
rect 121748 91838 121979 91840
rect 121748 91836 121754 91838
rect 121913 91835 121979 91838
rect 126462 91836 126468 91900
rect 126532 91898 126538 91900
rect 126605 91898 126671 91901
rect 126532 91896 126671 91898
rect 126532 91840 126610 91896
rect 126666 91840 126671 91896
rect 126532 91838 126671 91840
rect 126532 91836 126538 91838
rect 126605 91835 126671 91838
rect 74758 91700 74764 91764
rect 74828 91762 74834 91764
rect 75729 91762 75795 91765
rect 95049 91764 95115 91765
rect 94998 91762 95004 91764
rect 74828 91760 75795 91762
rect 74828 91704 75734 91760
rect 75790 91704 75795 91760
rect 74828 91702 75795 91704
rect 94958 91702 95004 91762
rect 95068 91760 95115 91764
rect 95110 91704 95115 91760
rect 74828 91700 74834 91702
rect 75729 91699 75795 91702
rect 94998 91700 95004 91702
rect 95068 91700 95115 91704
rect 96654 91700 96660 91764
rect 96724 91762 96730 91764
rect 97809 91762 97875 91765
rect 100569 91764 100635 91765
rect 100518 91762 100524 91764
rect 96724 91760 97875 91762
rect 96724 91704 97814 91760
rect 97870 91704 97875 91760
rect 96724 91702 97875 91704
rect 100478 91702 100524 91762
rect 100588 91760 100635 91764
rect 100630 91704 100635 91760
rect 96724 91700 96730 91702
rect 95049 91699 95115 91700
rect 97809 91699 97875 91702
rect 100518 91700 100524 91702
rect 100588 91700 100635 91704
rect 100569 91699 100635 91700
rect 92606 91564 92612 91628
rect 92676 91626 92682 91628
rect 93209 91626 93275 91629
rect 96337 91628 96403 91629
rect 96286 91626 96292 91628
rect 92676 91624 93275 91626
rect 92676 91568 93214 91624
rect 93270 91568 93275 91624
rect 92676 91566 93275 91568
rect 96246 91566 96292 91626
rect 96356 91624 96403 91628
rect 96398 91568 96403 91624
rect 92676 91564 92682 91566
rect 93209 91563 93275 91566
rect 96286 91564 96292 91566
rect 96356 91564 96403 91568
rect 97206 91564 97212 91628
rect 97276 91626 97282 91628
rect 97533 91626 97599 91629
rect 97276 91624 97599 91626
rect 97276 91568 97538 91624
rect 97594 91568 97599 91624
rect 97276 91566 97599 91568
rect 97276 91564 97282 91566
rect 96337 91563 96403 91564
rect 97533 91563 97599 91566
rect 98494 91564 98500 91628
rect 98564 91626 98570 91628
rect 99281 91626 99347 91629
rect 98564 91624 99347 91626
rect 98564 91568 99286 91624
rect 99342 91568 99347 91624
rect 98564 91566 99347 91568
rect 98564 91564 98570 91566
rect 99281 91563 99347 91566
rect 115473 91492 115539 91493
rect 122833 91492 122899 91493
rect 115422 91490 115428 91492
rect 115382 91430 115428 91490
rect 115492 91488 115539 91492
rect 115534 91432 115539 91488
rect 115422 91428 115428 91430
rect 115492 91428 115539 91432
rect 122782 91428 122788 91492
rect 122852 91490 122899 91492
rect 122852 91488 122944 91490
rect 122894 91432 122944 91488
rect 122852 91430 122944 91432
rect 122852 91428 122899 91430
rect 124438 91428 124444 91492
rect 124508 91490 124514 91492
rect 125317 91490 125383 91493
rect 124508 91488 125383 91490
rect 124508 91432 125322 91488
rect 125378 91432 125383 91488
rect 124508 91430 125383 91432
rect 124508 91428 124514 91430
rect 115473 91427 115539 91428
rect 122833 91427 122899 91428
rect 125317 91427 125383 91430
rect 101990 91292 101996 91356
rect 102060 91354 102066 91356
rect 180149 91354 180215 91357
rect 102060 91352 180215 91354
rect 102060 91296 180154 91352
rect 180210 91296 180215 91352
rect 102060 91294 180215 91296
rect 102060 91292 102066 91294
rect 180149 91291 180215 91294
rect 86769 91220 86835 91221
rect 99097 91220 99163 91221
rect 104617 91220 104683 91221
rect 86718 91218 86724 91220
rect 86678 91158 86724 91218
rect 86788 91216 86835 91220
rect 99046 91218 99052 91220
rect 86830 91160 86835 91216
rect 86718 91156 86724 91158
rect 86788 91156 86835 91160
rect 99006 91158 99052 91218
rect 99116 91216 99163 91220
rect 104566 91218 104572 91220
rect 99158 91160 99163 91216
rect 99046 91156 99052 91158
rect 99116 91156 99163 91160
rect 104526 91158 104572 91218
rect 104636 91216 104683 91220
rect 104678 91160 104683 91216
rect 104566 91156 104572 91158
rect 104636 91156 104683 91160
rect 116710 91156 116716 91220
rect 116780 91156 116786 91220
rect 123150 91156 123156 91220
rect 123220 91218 123226 91220
rect 123569 91218 123635 91221
rect 126697 91220 126763 91221
rect 130745 91220 130811 91221
rect 126646 91218 126652 91220
rect 123220 91216 123635 91218
rect 123220 91160 123574 91216
rect 123630 91160 123635 91216
rect 123220 91158 123635 91160
rect 126606 91158 126652 91218
rect 126716 91216 126763 91220
rect 130694 91218 130700 91220
rect 126758 91160 126763 91216
rect 123220 91156 123226 91158
rect 86769 91155 86835 91156
rect 99097 91155 99163 91156
rect 104617 91155 104683 91156
rect 116718 91082 116778 91156
rect 123569 91155 123635 91158
rect 126646 91156 126652 91158
rect 126716 91156 126763 91160
rect 130654 91158 130700 91218
rect 130764 91216 130811 91220
rect 130806 91160 130811 91216
rect 130694 91156 130700 91158
rect 130764 91156 130811 91160
rect 133086 91156 133092 91220
rect 133156 91218 133162 91220
rect 133321 91218 133387 91221
rect 133156 91216 133387 91218
rect 133156 91160 133326 91216
rect 133382 91160 133387 91216
rect 133156 91158 133387 91160
rect 133156 91156 133162 91158
rect 126697 91155 126763 91156
rect 130745 91155 130811 91156
rect 133321 91155 133387 91158
rect 166206 91082 166212 91084
rect 116718 91022 166212 91082
rect 166206 91020 166212 91022
rect 166276 91020 166282 91084
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580257 46338 580323 46341
rect 583520 46338 584960 46428
rect 580257 46336 584960 46338
rect 580257 46280 580262 46336
rect 580318 46280 584960 46336
rect 580257 46278 584960 46280
rect 580257 46275 580323 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 280660 286044 280724 286108
rect 285628 285908 285692 285972
rect 284340 285636 284404 285700
rect 287652 284684 287716 284748
rect 278820 284412 278884 284476
rect 243308 284064 243372 284068
rect 243308 284008 243358 284064
rect 243358 284008 243372 284064
rect 243308 284004 243372 284008
rect 288940 277476 289004 277540
rect 199516 260884 199580 260948
rect 244044 252452 244108 252516
rect 200620 250276 200684 250340
rect 200804 246196 200868 246260
rect 243492 244836 243556 244900
rect 200804 244564 200868 244628
rect 243676 241844 243740 241908
rect 279004 237900 279068 237964
rect 284708 233820 284772 233884
rect 284524 232596 284588 232660
rect 284892 232460 284956 232524
rect 199516 231100 199580 231164
rect 281580 231100 281644 231164
rect 281764 186900 281828 186964
rect 230428 182956 230492 183020
rect 282132 182820 282196 182884
rect 200988 181460 201052 181524
rect 281948 181324 282012 181388
rect 285812 180100 285876 180164
rect 200620 177652 200684 177716
rect 233188 177516 233252 177580
rect 279740 177516 279804 177580
rect 200804 177380 200868 177444
rect 280292 177244 280356 177308
rect 97028 176700 97092 176764
rect 106964 176760 107028 176764
rect 106964 176704 107014 176760
rect 107014 176704 107028 176760
rect 106964 176700 107028 176704
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 109540 176700 109604 176764
rect 110644 176760 110708 176764
rect 110644 176704 110694 176760
rect 110694 176704 110708 176760
rect 110644 176700 110708 176704
rect 112116 176700 112180 176764
rect 113220 176700 113284 176764
rect 114324 176760 114388 176764
rect 114324 176704 114374 176760
rect 114374 176704 114388 176760
rect 114324 176700 114388 176704
rect 115796 176760 115860 176764
rect 115796 176704 115846 176760
rect 115846 176704 115860 176760
rect 115796 176700 115860 176704
rect 116900 176760 116964 176764
rect 116900 176704 116950 176760
rect 116950 176704 116964 176760
rect 116900 176700 116964 176704
rect 118372 176760 118436 176764
rect 118372 176704 118422 176760
rect 118422 176704 118436 176760
rect 118372 176700 118436 176704
rect 120764 176760 120828 176764
rect 120764 176704 120814 176760
rect 120814 176704 120828 176760
rect 120764 176700 120828 176704
rect 121868 176700 121932 176764
rect 124444 176760 124508 176764
rect 124444 176704 124494 176760
rect 124494 176704 124508 176760
rect 124444 176700 124508 176704
rect 127020 176700 127084 176764
rect 129412 176760 129476 176764
rect 129412 176704 129462 176760
rect 129462 176704 129476 176760
rect 129412 176700 129476 176704
rect 130700 176700 130764 176764
rect 133092 176760 133156 176764
rect 133092 176704 133142 176760
rect 133142 176704 133156 176760
rect 133092 176700 133156 176704
rect 134380 176700 134444 176764
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 103284 176428 103348 176492
rect 135668 175536 135732 175540
rect 135668 175480 135718 175536
rect 135718 175480 135732 175536
rect 135668 175476 135732 175480
rect 98316 175400 98380 175404
rect 98316 175344 98366 175400
rect 98366 175344 98380 175400
rect 98316 175340 98380 175344
rect 99420 175400 99484 175404
rect 99420 175344 99470 175400
rect 99470 175344 99484 175400
rect 99420 175340 99484 175344
rect 100708 175400 100772 175404
rect 100708 175344 100758 175400
rect 100758 175344 100772 175400
rect 100708 175340 100772 175344
rect 101996 175400 102060 175404
rect 101996 175344 102046 175400
rect 102046 175344 102060 175400
rect 101996 175340 102060 175344
rect 104572 175400 104636 175404
rect 104572 175344 104622 175400
rect 104622 175344 104636 175400
rect 104572 175340 104636 175344
rect 105676 175400 105740 175404
rect 105676 175344 105726 175400
rect 105726 175344 105740 175400
rect 105676 175340 105740 175344
rect 128124 175400 128188 175404
rect 128124 175344 128174 175400
rect 128174 175344 128188 175400
rect 128124 175340 128188 175344
rect 131988 175400 132052 175404
rect 131988 175344 132038 175400
rect 132038 175344 132052 175400
rect 131988 175340 132052 175344
rect 158852 175400 158916 175404
rect 158852 175344 158902 175400
rect 158902 175344 158916 175400
rect 158852 175340 158916 175344
rect 119398 174992 119462 174996
rect 119398 174936 119434 174992
rect 119434 174936 119462 174992
rect 119398 174932 119462 174936
rect 123070 174992 123134 174996
rect 123070 174936 123114 174992
rect 123114 174936 123134 174992
rect 123070 174932 123134 174936
rect 125654 174992 125718 174996
rect 125654 174936 125690 174992
rect 125690 174936 125718 174992
rect 279740 175204 279804 175268
rect 125654 174932 125718 174936
rect 268332 174524 268396 174588
rect 267780 174388 267844 174452
rect 281948 173980 282012 174044
rect 279372 172076 279436 172140
rect 279556 169764 279620 169828
rect 281764 166228 281828 166292
rect 282132 163916 282196 163980
rect 281580 163100 281644 163164
rect 268516 162964 268580 163028
rect 244044 162420 244108 162484
rect 268516 159836 268580 159900
rect 268516 153444 268580 153508
rect 268516 153036 268580 153100
rect 288940 151812 289004 151876
rect 280660 150452 280724 150516
rect 242940 149092 243004 149156
rect 268332 147868 268396 147932
rect 285628 147052 285692 147116
rect 268332 146100 268396 146164
rect 284892 145420 284956 145484
rect 284708 144740 284772 144804
rect 284524 143108 284588 143172
rect 268516 142292 268580 142356
rect 268516 141884 268580 141948
rect 230428 140660 230492 140724
rect 284340 140796 284404 140860
rect 164924 138212 164988 138276
rect 166212 136852 166276 136916
rect 233188 136308 233252 136372
rect 268332 136308 268396 136372
rect 268148 135764 268212 135828
rect 268516 134132 268580 134196
rect 268516 133724 268580 133788
rect 268516 127196 268580 127260
rect 268516 126788 268580 126852
rect 268516 122980 268580 123044
rect 268516 122572 268580 122636
rect 268516 121620 268580 121684
rect 268516 121212 268580 121276
rect 267780 115908 267844 115972
rect 268332 116044 268396 116108
rect 285812 115500 285876 115564
rect 287652 111828 287716 111892
rect 214420 103532 214484 103596
rect 268516 102308 268580 102372
rect 213868 101084 213932 101148
rect 280292 100812 280356 100876
rect 268516 100540 268580 100604
rect 268332 97140 268396 97204
rect 166396 96596 166460 96660
rect 267780 96868 267844 96932
rect 213868 94828 213932 94892
rect 214420 94692 214484 94756
rect 166396 94556 166460 94620
rect 151630 94344 151694 94348
rect 151630 94288 151634 94344
rect 151634 94288 151690 94344
rect 151690 94288 151694 94344
rect 151630 94284 151694 94288
rect 124076 94208 124140 94212
rect 124076 94152 124126 94208
rect 124126 94152 124140 94208
rect 124076 94148 124140 94152
rect 117084 94072 117148 94076
rect 117084 94016 117134 94072
rect 117134 94016 117148 94072
rect 117084 94012 117148 94016
rect 122052 94072 122116 94076
rect 122052 94016 122102 94072
rect 122102 94016 122116 94072
rect 122052 94012 122116 94016
rect 151676 94072 151740 94076
rect 151676 94016 151726 94072
rect 151726 94016 151740 94072
rect 151676 94012 151740 94016
rect 118188 93936 118252 93940
rect 118188 93880 118238 93936
rect 118238 93880 118252 93936
rect 118188 93876 118252 93880
rect 151492 93936 151556 93940
rect 151492 93880 151542 93936
rect 151542 93880 151556 93936
rect 151492 93876 151556 93880
rect 100892 93740 100956 93804
rect 102916 93664 102980 93668
rect 102916 93608 102966 93664
rect 102966 93608 102980 93664
rect 102916 93604 102980 93608
rect 104204 93664 104268 93668
rect 104204 93608 104254 93664
rect 104254 93608 104268 93664
rect 104204 93604 104268 93608
rect 105492 93664 105556 93668
rect 105492 93608 105542 93664
rect 105542 93608 105556 93664
rect 105492 93604 105556 93608
rect 106412 93664 106476 93668
rect 106412 93608 106462 93664
rect 106462 93608 106476 93664
rect 106412 93604 106476 93608
rect 107700 93664 107764 93668
rect 107700 93608 107750 93664
rect 107750 93608 107764 93664
rect 107700 93604 107764 93608
rect 109172 93664 109236 93668
rect 109172 93608 109222 93664
rect 109222 93608 109236 93664
rect 109172 93604 109236 93608
rect 119660 93664 119724 93668
rect 119660 93608 119710 93664
rect 119710 93608 119724 93664
rect 119660 93604 119724 93608
rect 90220 93528 90284 93532
rect 90220 93472 90270 93528
rect 90270 93472 90284 93528
rect 90220 93468 90284 93472
rect 101812 93528 101876 93532
rect 101812 93472 101862 93528
rect 101862 93472 101876 93528
rect 101812 93468 101876 93472
rect 111380 93468 111444 93532
rect 119292 93468 119356 93532
rect 164924 93604 164988 93668
rect 125364 93528 125428 93532
rect 125364 93472 125414 93528
rect 125414 93472 125428 93528
rect 125364 93468 125428 93472
rect 135668 93392 135732 93396
rect 135668 93336 135718 93392
rect 135718 93336 135732 93392
rect 135668 93332 135732 93336
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 128124 93256 128188 93260
rect 128124 93200 128174 93256
rect 128174 93200 128188 93256
rect 128124 93196 128188 93200
rect 113036 92516 113100 92580
rect 84332 92440 84396 92444
rect 84332 92384 84382 92440
rect 84382 92384 84396 92440
rect 84332 92380 84396 92384
rect 85804 92380 85868 92444
rect 88012 92440 88076 92444
rect 88012 92384 88062 92440
rect 88062 92384 88076 92440
rect 88012 92380 88076 92384
rect 88932 92380 88996 92444
rect 91324 92380 91388 92444
rect 93900 92380 93964 92444
rect 99972 92440 100036 92444
rect 99972 92384 100022 92440
rect 100022 92384 100036 92440
rect 99972 92380 100036 92384
rect 105676 92440 105740 92444
rect 105676 92384 105726 92440
rect 105726 92384 105740 92440
rect 105676 92380 105740 92384
rect 108068 92440 108132 92444
rect 108068 92384 108118 92440
rect 108118 92384 108132 92440
rect 108068 92380 108132 92384
rect 109540 92380 109604 92444
rect 110644 92380 110708 92444
rect 111932 92440 111996 92444
rect 111932 92384 111982 92440
rect 111982 92384 111996 92440
rect 111932 92380 111996 92384
rect 112300 92440 112364 92444
rect 112300 92384 112350 92440
rect 112350 92384 112364 92440
rect 112300 92380 112364 92384
rect 113220 92380 113284 92444
rect 114324 92440 114388 92444
rect 114324 92384 114374 92440
rect 114374 92384 114388 92440
rect 114324 92380 114388 92384
rect 114876 92380 114940 92444
rect 115796 92440 115860 92444
rect 115796 92384 115846 92440
rect 115846 92384 115860 92440
rect 115796 92380 115860 92384
rect 118004 92440 118068 92444
rect 118004 92384 118054 92440
rect 118054 92384 118068 92440
rect 118004 92380 118068 92384
rect 120212 92440 120276 92444
rect 120212 92384 120262 92440
rect 120262 92384 120276 92440
rect 120212 92380 120276 92384
rect 120580 92380 120644 92444
rect 125732 92440 125796 92444
rect 125732 92384 125782 92440
rect 125782 92384 125796 92440
rect 125732 92380 125796 92384
rect 129412 92440 129476 92444
rect 129412 92384 129462 92440
rect 129462 92384 129476 92440
rect 129412 92380 129476 92384
rect 132356 92440 132420 92444
rect 132356 92384 132406 92440
rect 132406 92384 132420 92440
rect 132356 92380 132420 92384
rect 134380 92440 134444 92444
rect 134380 92384 134430 92440
rect 134430 92384 134444 92440
rect 134380 92380 134444 92384
rect 152044 92380 152108 92444
rect 98132 92244 98196 92308
rect 103836 92108 103900 92172
rect 106780 91972 106844 92036
rect 121684 91836 121748 91900
rect 126468 91836 126532 91900
rect 74764 91700 74828 91764
rect 95004 91760 95068 91764
rect 95004 91704 95054 91760
rect 95054 91704 95068 91760
rect 95004 91700 95068 91704
rect 96660 91700 96724 91764
rect 100524 91760 100588 91764
rect 100524 91704 100574 91760
rect 100574 91704 100588 91760
rect 100524 91700 100588 91704
rect 92612 91564 92676 91628
rect 96292 91624 96356 91628
rect 96292 91568 96342 91624
rect 96342 91568 96356 91624
rect 96292 91564 96356 91568
rect 97212 91564 97276 91628
rect 98500 91564 98564 91628
rect 115428 91488 115492 91492
rect 115428 91432 115478 91488
rect 115478 91432 115492 91488
rect 115428 91428 115492 91432
rect 122788 91488 122852 91492
rect 122788 91432 122838 91488
rect 122838 91432 122852 91488
rect 122788 91428 122852 91432
rect 124444 91428 124508 91492
rect 101996 91292 102060 91356
rect 86724 91216 86788 91220
rect 86724 91160 86774 91216
rect 86774 91160 86788 91216
rect 86724 91156 86788 91160
rect 99052 91216 99116 91220
rect 99052 91160 99102 91216
rect 99102 91160 99116 91216
rect 99052 91156 99116 91160
rect 104572 91216 104636 91220
rect 104572 91160 104622 91216
rect 104622 91160 104636 91216
rect 104572 91156 104636 91160
rect 116716 91156 116780 91220
rect 123156 91156 123220 91220
rect 126652 91216 126716 91220
rect 126652 91160 126702 91216
rect 126702 91160 126716 91216
rect 126652 91156 126716 91160
rect 130700 91216 130764 91220
rect 130700 91160 130750 91216
rect 130750 91160 130764 91216
rect 130700 91156 130764 91160
rect 133092 91156 133156 91220
rect 166212 91020 166276 91084
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176600 67574 212058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 176764 97093 176765
rect 97027 176700 97028 176764
rect 97092 176700 97093 176764
rect 97027 176699 97093 176700
rect 97030 175130 97090 176699
rect 99234 176600 99854 208338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176600 103574 212058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 106963 176764 107029 176765
rect 106963 176700 106964 176764
rect 107028 176700 107029 176764
rect 106963 176699 107029 176700
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 98315 175404 98381 175405
rect 98315 175340 98316 175404
rect 98380 175340 98381 175404
rect 98315 175339 98381 175340
rect 99419 175404 99485 175405
rect 99419 175340 99420 175404
rect 99484 175340 99485 175404
rect 99419 175339 99485 175340
rect 100707 175404 100773 175405
rect 100707 175340 100708 175404
rect 100772 175340 100773 175404
rect 100707 175339 100773 175340
rect 101995 175404 102061 175405
rect 101995 175340 101996 175404
rect 102060 175340 102061 175404
rect 101995 175339 102061 175340
rect 96960 175070 97090 175130
rect 98318 175130 98378 175339
rect 99422 175130 99482 175339
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 175339
rect 101998 175130 102058 175339
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104571 175404 104637 175405
rect 104571 175340 104572 175404
rect 104636 175340 104637 175404
rect 104571 175339 104637 175340
rect 105675 175404 105741 175405
rect 105675 175340 105676 175404
rect 105740 175340 105741 175404
rect 105675 175339 105741 175340
rect 104574 175130 104634 175339
rect 105678 175130 105738 175339
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 176699
rect 108070 175130 108130 176699
rect 109542 175130 109602 176699
rect 109794 176600 110414 182898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 110643 176764 110709 176765
rect 110643 176700 110644 176764
rect 110708 176700 110709 176764
rect 110643 176699 110709 176700
rect 112115 176764 112181 176765
rect 112115 176700 112116 176764
rect 112180 176700 112181 176764
rect 112115 176699 112181 176700
rect 113219 176764 113285 176765
rect 113219 176700 113220 176764
rect 113284 176700 113285 176764
rect 113219 176699 113285 176700
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 176699
rect 112118 175130 112178 176699
rect 113222 175130 113282 176699
rect 113514 176600 114134 186618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 114323 176764 114389 176765
rect 114323 176700 114324 176764
rect 114388 176700 114389 176764
rect 114323 176699 114389 176700
rect 115795 176764 115861 176765
rect 115795 176700 115796 176764
rect 115860 176700 115861 176764
rect 115795 176699 115861 176700
rect 116899 176764 116965 176765
rect 116899 176700 116900 176764
rect 116964 176700 116965 176764
rect 116899 176699 116965 176700
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 176699
rect 115798 175130 115858 176699
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 176699
rect 117234 176600 117854 190338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 118371 176764 118437 176765
rect 118371 176700 118372 176764
rect 118436 176700 118437 176764
rect 118371 176699 118437 176700
rect 120763 176764 120829 176765
rect 120763 176700 120764 176764
rect 120828 176700 120829 176764
rect 120763 176699 120829 176700
rect 118374 175130 118434 176699
rect 120766 175130 120826 176699
rect 120954 176600 121574 194058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 121867 176764 121933 176765
rect 121867 176700 121868 176764
rect 121932 176700 121933 176764
rect 121867 176699 121933 176700
rect 124443 176764 124509 176765
rect 124443 176700 124444 176764
rect 124508 176700 124509 176764
rect 124443 176699 124509 176700
rect 127019 176764 127085 176765
rect 127019 176700 127020 176764
rect 127084 176700 127085 176764
rect 127019 176699 127085 176700
rect 121870 175130 121930 176699
rect 124446 175130 124506 176699
rect 127022 175130 127082 176699
rect 127794 176600 128414 200898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 129411 176764 129477 176765
rect 129411 176700 129412 176764
rect 129476 176700 129477 176764
rect 129411 176699 129477 176700
rect 130699 176764 130765 176765
rect 130699 176700 130700 176764
rect 130764 176700 130765 176764
rect 130699 176699 130765 176700
rect 128123 175404 128189 175405
rect 128123 175340 128124 175404
rect 128188 175340 128189 175404
rect 128123 175339 128189 175340
rect 128126 175130 128186 175339
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 124432 175070 124506 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 176699
rect 130702 175130 130762 176699
rect 131514 176600 132134 204618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 133091 176764 133157 176765
rect 133091 176700 133092 176764
rect 133156 176700 133157 176764
rect 133091 176699 133157 176700
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 131987 175404 132053 175405
rect 131987 175340 131988 175404
rect 132052 175340 132053 175404
rect 131987 175339 132053 175340
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119397 174996 119463 174997
rect 119397 174932 119398 174996
rect 119462 174932 119463 174996
rect 119397 174931 119463 174932
rect 119400 174494 119460 174931
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123069 174996 123135 174997
rect 123069 174932 123070 174996
rect 123134 174932 123135 174996
rect 123069 174931 123135 174932
rect 123072 174494 123132 174931
rect 124432 174494 124492 175070
rect 125653 174996 125719 174997
rect 125653 174932 125654 174996
rect 125718 174932 125719 174996
rect 125653 174931 125719 174932
rect 125656 174494 125716 174931
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 131990 175130 132050 175339
rect 133094 175130 133154 176699
rect 134382 175130 134442 176699
rect 135234 176600 135854 208338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176600 139574 212058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 135667 175540 135733 175541
rect 135667 175476 135668 175540
rect 135732 175476 135733 175540
rect 135667 175475 135733 175476
rect 131990 175070 132108 175130
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135670 175130 135730 175475
rect 148182 175130 148242 176699
rect 149514 176600 150134 186618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 176600 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 158851 175404 158917 175405
rect 158851 175340 158852 175404
rect 158916 175340 158917 175404
rect 158851 175339 158917 175340
rect 158854 175130 158914 175339
rect 135670 175070 135780 175130
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 164923 138276 164989 138277
rect 164923 138212 164924 138276
rect 164988 138212 164989 138276
rect 164923 138211 164989 138212
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85866 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 93100
rect 74766 91765 74826 94830
rect 74763 91764 74829 91765
rect 74763 91700 74764 91764
rect 74828 91700 74829 91764
rect 74763 91699 74829 91700
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 92445 84394 94830
rect 84331 92444 84397 92445
rect 84331 92380 84332 92444
rect 84396 92380 84397 92444
rect 84331 92379 84397 92380
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 85806 92445 85866 94830
rect 85803 92444 85869 92445
rect 85803 92380 85804 92444
rect 85868 92380 85869 92444
rect 85803 92379 85869 92380
rect 86726 91221 86786 94830
rect 88014 92445 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 92445 88994 94830
rect 90222 93533 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 90219 93532 90285 93533
rect 90219 93468 90220 93532
rect 90284 93468 90285 93532
rect 90219 93467 90285 93468
rect 91326 92445 91386 94830
rect 88011 92444 88077 92445
rect 88011 92380 88012 92444
rect 88076 92380 88077 92444
rect 88011 92379 88077 92380
rect 88931 92444 88997 92445
rect 88931 92380 88932 92444
rect 88996 92380 88997 92444
rect 88931 92379 88997 92380
rect 91323 92444 91389 92445
rect 91323 92380 91324 92444
rect 91388 92380 91389 92444
rect 91323 92379 91389 92380
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91629 92674 94830
rect 93902 92445 93962 94830
rect 93899 92444 93965 92445
rect 93899 92380 93900 92444
rect 93964 92380 93965 92444
rect 93899 92379 93965 92380
rect 95006 91765 95066 94830
rect 95003 91764 95069 91765
rect 95003 91700 95004 91764
rect 95068 91700 95069 91764
rect 95003 91699 95069 91700
rect 92611 91628 92677 91629
rect 92611 91564 92612 91628
rect 92676 91564 92677 91628
rect 92611 91563 92677 91564
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91629 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91765 96722 94830
rect 96659 91764 96725 91765
rect 96659 91700 96660 91764
rect 96724 91700 96725 91764
rect 96659 91699 96725 91700
rect 97214 91629 97274 94830
rect 98134 92309 98194 94830
rect 98131 92308 98197 92309
rect 98131 92244 98132 92308
rect 98196 92244 98197 92308
rect 98131 92243 98197 92244
rect 98502 91629 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 99544 94830 100034 94890
rect 96291 91628 96357 91629
rect 96291 91564 96292 91628
rect 96356 91564 96357 91628
rect 96291 91563 96357 91564
rect 97211 91628 97277 91629
rect 97211 91564 97212 91628
rect 97276 91564 97277 91628
rect 97211 91563 97277 91564
rect 98499 91628 98565 91629
rect 98499 91564 98500 91628
rect 98564 91564 98565 91628
rect 98499 91563 98565 91564
rect 99054 91221 99114 94830
rect 99051 91220 99117 91221
rect 99051 91156 99052 91220
rect 99116 91156 99117 91220
rect 99051 91155 99117 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 92445 100034 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 99971 92444 100037 92445
rect 99971 92380 99972 92444
rect 100036 92380 100037 92444
rect 99971 92379 100037 92380
rect 100526 91765 100586 94830
rect 100894 93805 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 100891 93804 100957 93805
rect 100891 93740 100892 93804
rect 100956 93740 100957 93804
rect 100891 93739 100957 93740
rect 101814 93533 101874 94830
rect 101811 93532 101877 93533
rect 101811 93468 101812 93532
rect 101876 93468 101877 93532
rect 101811 93467 101877 93468
rect 100523 91764 100589 91765
rect 100523 91700 100524 91764
rect 100588 91700 100589 91764
rect 100523 91699 100589 91700
rect 101998 91357 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 102918 93669 102978 94830
rect 102915 93668 102981 93669
rect 102915 93604 102916 93668
rect 102980 93604 102981 93668
rect 102915 93603 102981 93604
rect 103286 93530 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 104206 93669 104266 94830
rect 104203 93668 104269 93669
rect 104203 93604 104204 93668
rect 104268 93604 104269 93668
rect 104203 93603 104269 93604
rect 103286 93470 103714 93530
rect 101995 91356 102061 91357
rect 101995 91292 101996 91356
rect 102060 91292 102061 91356
rect 101995 91291 102061 91292
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 103654 92170 103714 93470
rect 103835 92172 103901 92173
rect 103835 92170 103836 92172
rect 103654 92110 103836 92170
rect 103835 92108 103836 92110
rect 103900 92108 103901 92172
rect 103835 92107 103901 92108
rect 104574 91221 104634 94830
rect 105494 93669 105554 94830
rect 105491 93668 105557 93669
rect 105491 93604 105492 93668
rect 105556 93604 105557 93668
rect 105491 93603 105557 93604
rect 105678 92445 105738 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106616 94830 106842 94890
rect 106414 93669 106474 94830
rect 106411 93668 106477 93669
rect 106411 93604 106412 93668
rect 106476 93604 106477 93668
rect 106411 93603 106477 93604
rect 105675 92444 105741 92445
rect 105675 92380 105676 92444
rect 105740 92380 105741 92444
rect 105675 92379 105741 92380
rect 106782 92037 106842 94830
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 107702 93669 107762 94830
rect 107699 93668 107765 93669
rect 107699 93604 107700 93668
rect 107764 93604 107765 93668
rect 107699 93603 107765 93604
rect 108070 92445 108130 94830
rect 109174 93669 109234 94830
rect 109171 93668 109237 93669
rect 109171 93604 109172 93668
rect 109236 93604 109237 93668
rect 109171 93603 109237 93604
rect 109542 92445 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111240 94890 111300 95200
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 111240 94830 111442 94890
rect 111920 94830 111994 94890
rect 110094 93261 110154 94830
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 108067 92444 108133 92445
rect 108067 92380 108068 92444
rect 108132 92380 108133 92444
rect 108067 92379 108133 92380
rect 109539 92444 109605 92445
rect 109539 92380 109540 92444
rect 109604 92380 109605 92444
rect 109539 92379 109605 92380
rect 106779 92036 106845 92037
rect 106779 91972 106780 92036
rect 106844 91972 106845 92036
rect 106779 91971 106845 91972
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 92445 110706 94830
rect 111382 93533 111442 94830
rect 111379 93532 111445 93533
rect 111379 93468 111380 93532
rect 111444 93468 111445 93532
rect 111379 93467 111445 93468
rect 111934 92445 111994 94830
rect 112302 94830 112388 94890
rect 113038 94830 113204 94890
rect 113406 94830 113748 94890
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 112302 92445 112362 94830
rect 113038 92581 113098 94830
rect 113406 93870 113466 94830
rect 113222 93810 113466 93870
rect 113035 92580 113101 92581
rect 113035 92516 113036 92580
rect 113100 92516 113101 92580
rect 113035 92515 113101 92516
rect 113222 92445 113282 93810
rect 110643 92444 110709 92445
rect 110643 92380 110644 92444
rect 110708 92380 110709 92444
rect 110643 92379 110709 92380
rect 111931 92444 111997 92445
rect 111931 92380 111932 92444
rect 111996 92380 111997 92444
rect 111931 92379 111997 92380
rect 112299 92444 112365 92445
rect 112299 92380 112300 92444
rect 112364 92380 112365 92444
rect 112299 92379 112365 92380
rect 113219 92444 113285 92445
rect 113219 92380 113220 92444
rect 113284 92380 113285 92444
rect 113219 92379 113285 92380
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 92445 114386 94830
rect 114878 92445 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 114323 92444 114389 92445
rect 114323 92380 114324 92444
rect 114388 92380 114389 92444
rect 114323 92379 114389 92380
rect 114875 92444 114941 92445
rect 114875 92380 114876 92444
rect 114940 92380 114941 92444
rect 114875 92379 114941 92380
rect 115430 91493 115490 94830
rect 115798 92445 115858 94830
rect 115795 92444 115861 92445
rect 115795 92380 115796 92444
rect 115860 92380 115861 92444
rect 115795 92379 115861 92380
rect 115427 91492 115493 91493
rect 115427 91428 115428 91492
rect 115492 91428 115493 91492
rect 115427 91427 115493 91428
rect 116718 91221 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 117086 94077 117146 94830
rect 117083 94076 117149 94077
rect 117083 94012 117084 94076
rect 117148 94012 117149 94076
rect 117083 94011 117149 94012
rect 116715 91220 116781 91221
rect 116715 91156 116716 91220
rect 116780 91156 116781 91220
rect 116715 91155 116781 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 92445 118066 94830
rect 118190 93941 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 118187 93940 118253 93941
rect 118187 93876 118188 93940
rect 118252 93876 118253 93940
rect 118187 93875 118253 93876
rect 119294 93533 119354 94830
rect 119662 93669 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 119659 93668 119725 93669
rect 119659 93604 119660 93668
rect 119724 93604 119725 93668
rect 119659 93603 119725 93604
rect 119291 93532 119357 93533
rect 119291 93468 119292 93532
rect 119356 93468 119357 93532
rect 119291 93467 119357 93468
rect 120214 92445 120274 94830
rect 120582 92445 120642 94830
rect 118003 92444 118069 92445
rect 118003 92380 118004 92444
rect 118068 92380 118069 92444
rect 118003 92379 118069 92380
rect 120211 92444 120277 92445
rect 120211 92380 120212 92444
rect 120276 92380 120277 92444
rect 120211 92379 120277 92380
rect 120579 92444 120645 92445
rect 120579 92380 120580 92444
rect 120644 92380 120645 92444
rect 120579 92379 120645 92380
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 121686 91901 121746 94830
rect 122054 94077 122114 94830
rect 122051 94076 122117 94077
rect 122051 94012 122052 94076
rect 122116 94012 122117 94076
rect 122051 94011 122117 94012
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 121683 91900 121749 91901
rect 121683 91836 121684 91900
rect 121748 91836 121749 91900
rect 121683 91835 121749 91836
rect 122606 91490 122666 93810
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 123158 91221 123218 94830
rect 124078 94213 124138 94830
rect 124075 94212 124141 94213
rect 124075 94148 124076 94212
rect 124140 94148 124141 94212
rect 124075 94147 124141 94148
rect 124446 91493 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 125366 93533 125426 94830
rect 125363 93532 125429 93533
rect 125363 93468 125364 93532
rect 125428 93468 125429 93532
rect 125363 93467 125429 93468
rect 125734 92445 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 126608 94830 126714 94890
rect 128104 94830 128186 94890
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 125731 92444 125797 92445
rect 125731 92380 125732 92444
rect 125796 92380 125797 92444
rect 125731 92379 125797 92380
rect 126470 91901 126530 94830
rect 126467 91900 126533 91901
rect 126467 91836 126468 91900
rect 126532 91836 126533 91900
rect 126467 91835 126533 91836
rect 124443 91492 124509 91493
rect 124443 91428 124444 91492
rect 124508 91428 124509 91492
rect 124443 91427 124509 91428
rect 126654 91221 126714 94830
rect 128126 93261 128186 94830
rect 128123 93260 128189 93261
rect 128123 93196 128124 93260
rect 128188 93196 128189 93260
rect 128123 93195 128189 93196
rect 123155 91220 123221 91221
rect 123155 91156 123156 91220
rect 123220 91156 123221 91220
rect 123155 91155 123221 91156
rect 126651 91220 126717 91221
rect 126651 91156 126652 91220
rect 126716 91156 126717 91220
rect 126651 91155 126717 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 129414 92445 129474 94830
rect 129411 92444 129477 92445
rect 129411 92380 129412 92444
rect 129476 92380 129477 92444
rect 129411 92379 129477 92380
rect 130702 91221 130762 94830
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 92445 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 135730 94890
rect 132355 92444 132421 92445
rect 132355 92380 132356 92444
rect 132420 92380 132421 92444
rect 132355 92379 132421 92380
rect 133094 91221 133154 94830
rect 134382 92445 134442 94830
rect 135670 93397 135730 94830
rect 151494 94830 151556 94890
rect 151494 93941 151554 94830
rect 151632 94349 151692 95200
rect 151629 94348 151695 94349
rect 151629 94284 151630 94348
rect 151694 94284 151695 94348
rect 151629 94283 151695 94284
rect 151768 94210 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151678 94150 151828 94210
rect 151678 94077 151738 94150
rect 151675 94076 151741 94077
rect 151675 94012 151676 94076
rect 151740 94012 151741 94076
rect 151675 94011 151741 94012
rect 151491 93940 151557 93941
rect 151491 93876 151492 93940
rect 151556 93876 151557 93940
rect 151491 93875 151557 93876
rect 135667 93396 135733 93397
rect 135667 93332 135668 93396
rect 135732 93332 135733 93396
rect 135667 93331 135733 93332
rect 134379 92444 134445 92445
rect 134379 92380 134380 92444
rect 134444 92380 134445 92444
rect 134379 92379 134445 92380
rect 133091 91220 133157 91221
rect 133091 91156 133092 91220
rect 133156 91156 133157 91220
rect 133091 91155 133157 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 152046 92445 152106 94830
rect 164926 93669 164986 138211
rect 166211 136916 166277 136917
rect 166211 136852 166212 136916
rect 166276 136852 166277 136916
rect 166211 136851 166277 136852
rect 164923 93668 164989 93669
rect 164923 93604 164924 93668
rect 164988 93604 164989 93668
rect 164923 93603 164989 93604
rect 152043 92444 152109 92445
rect 152043 92380 152044 92444
rect 152108 92380 152109 92444
rect 152043 92379 152109 92380
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 91085 166274 136851
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 166395 96660 166461 96661
rect 166395 96596 166396 96660
rect 166460 96596 166461 96660
rect 166395 96595 166461 96596
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166398 94621 166458 96595
rect 166395 94620 166461 94621
rect 166395 94556 166396 94620
rect 166460 94556 166461 94620
rect 166395 94555 166461 94556
rect 166211 91084 166277 91085
rect 166211 91020 166212 91084
rect 166276 91020 166277 91084
rect 166211 91019 166277 91020
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 286182 200414 308898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 286182 204134 312618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 286182 207854 316338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 286182 211574 320058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 286182 218414 290898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 286182 222134 294618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 286182 225854 298338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 286182 229574 302058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 286182 236414 308898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 286182 240134 312618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 286182 243854 316338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 243307 284068 243373 284069
rect 243307 284004 243308 284068
rect 243372 284004 243373 284068
rect 243307 284003 243373 284004
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 243310 277410 243370 284003
rect 243310 277350 243554 277410
rect 219768 273454 220088 273486
rect 219768 273218 219810 273454
rect 220046 273218 220088 273454
rect 219768 273134 220088 273218
rect 219768 272898 219810 273134
rect 220046 272898 220088 273134
rect 219768 272866 220088 272898
rect 243494 267750 243554 277350
rect 243494 267690 243738 267750
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 199515 260948 199581 260949
rect 199515 260884 199516 260948
rect 199580 260884 199581 260948
rect 199515 260883 199581 260884
rect 199518 231165 199578 260883
rect 204408 255454 204728 255486
rect 204408 255218 204450 255454
rect 204686 255218 204728 255454
rect 204408 255134 204728 255218
rect 204408 254898 204450 255134
rect 204686 254898 204728 255134
rect 204408 254866 204728 254898
rect 235128 255454 235448 255486
rect 235128 255218 235170 255454
rect 235406 255218 235448 255454
rect 235128 255134 235448 255218
rect 235128 254898 235170 255134
rect 235406 254898 235448 255134
rect 235128 254866 235448 254898
rect 200619 250340 200685 250341
rect 200619 250276 200620 250340
rect 200684 250276 200685 250340
rect 200619 250275 200685 250276
rect 199794 237454 200414 238182
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199515 231164 199581 231165
rect 199515 231100 199516 231164
rect 199580 231100 199581 231164
rect 199515 231099 199581 231100
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 200622 177717 200682 250275
rect 200803 246260 200869 246261
rect 200803 246196 200804 246260
rect 200868 246196 200869 246260
rect 200803 246195 200869 246196
rect 200806 245170 200866 246195
rect 200806 245110 201050 245170
rect 200803 244628 200869 244629
rect 200803 244564 200804 244628
rect 200868 244564 200869 244628
rect 200803 244563 200869 244564
rect 200619 177716 200685 177717
rect 200619 177652 200620 177716
rect 200684 177652 200685 177716
rect 200619 177651 200685 177652
rect 200806 177445 200866 244563
rect 200990 181525 201050 245110
rect 243491 244900 243557 244901
rect 243491 244836 243492 244900
rect 243556 244836 243557 244900
rect 243491 244835 243557 244836
rect 243494 238770 243554 244835
rect 243678 241909 243738 267690
rect 244043 252516 244109 252517
rect 244043 252452 244044 252516
rect 244108 252452 244109 252516
rect 244043 252451 244109 252452
rect 243675 241908 243741 241909
rect 243675 241844 243676 241908
rect 243740 241844 243741 241908
rect 243675 241843 243741 241844
rect 242942 238710 243554 238770
rect 203514 205174 204134 238182
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 200987 181524 201053 181525
rect 200987 181460 200988 181524
rect 201052 181460 201053 181524
rect 200987 181459 201053 181460
rect 200803 177444 200869 177445
rect 200803 177380 200804 177444
rect 200868 177380 200869 177444
rect 200803 177379 200869 177380
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 208894 207854 238182
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 212614 211574 238182
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 217794 219454 218414 238182
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 223174 222134 238182
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 225234 226894 225854 238182
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 228954 230614 229574 238182
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 178000 229574 194058
rect 235794 237454 236414 238182
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 230427 183020 230493 183021
rect 230427 182956 230428 183020
rect 230492 182956 230493 183020
rect 230427 182955 230493 182956
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 221207 165454 221527 165486
rect 221207 165218 221249 165454
rect 221485 165218 221527 165454
rect 221207 165134 221527 165218
rect 221207 164898 221249 165134
rect 221485 164898 221527 165134
rect 221207 164866 221527 164898
rect 224471 165454 224791 165486
rect 224471 165218 224513 165454
rect 224749 165218 224791 165454
rect 224471 165134 224791 165218
rect 224471 164898 224513 165134
rect 224749 164898 224791 165134
rect 224471 164866 224791 164898
rect 219575 147454 219895 147486
rect 219575 147218 219617 147454
rect 219853 147218 219895 147454
rect 219575 147134 219895 147218
rect 219575 146898 219617 147134
rect 219853 146898 219895 147134
rect 219575 146866 219895 146898
rect 222839 147454 223159 147486
rect 222839 147218 222881 147454
rect 223117 147218 223159 147454
rect 222839 147134 223159 147218
rect 222839 146898 222881 147134
rect 223117 146898 223159 147134
rect 222839 146866 223159 146898
rect 226103 147454 226423 147486
rect 226103 147218 226145 147454
rect 226381 147218 226423 147454
rect 226103 147134 226423 147218
rect 226103 146898 226145 147134
rect 226381 146898 226423 147134
rect 226103 146866 226423 146898
rect 230430 140725 230490 182955
rect 233187 177580 233253 177581
rect 233187 177516 233188 177580
rect 233252 177516 233253 177580
rect 233187 177515 233253 177516
rect 230427 140724 230493 140725
rect 230427 140660 230428 140724
rect 230492 140660 230493 140724
rect 230427 140659 230493 140660
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 233190 136373 233250 177515
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 233187 136372 233253 136373
rect 233187 136308 233188 136372
rect 233252 136308 233253 136372
rect 233187 136307 233253 136308
rect 221207 129454 221527 129486
rect 221207 129218 221249 129454
rect 221485 129218 221527 129454
rect 221207 129134 221527 129218
rect 221207 128898 221249 129134
rect 221485 128898 221527 129134
rect 221207 128866 221527 128898
rect 224471 129454 224791 129486
rect 224471 129218 224513 129454
rect 224749 129218 224791 129454
rect 224471 129134 224791 129218
rect 224471 128898 224513 129134
rect 224749 128898 224791 129134
rect 224471 128866 224791 128898
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 219575 111454 219895 111486
rect 219575 111218 219617 111454
rect 219853 111218 219895 111454
rect 219575 111134 219895 111218
rect 219575 110898 219617 111134
rect 219853 110898 219895 111134
rect 219575 110866 219895 110898
rect 222839 111454 223159 111486
rect 222839 111218 222881 111454
rect 223117 111218 223159 111454
rect 222839 111134 223159 111218
rect 222839 110898 222881 111134
rect 223117 110898 223159 111134
rect 222839 110866 223159 110898
rect 226103 111454 226423 111486
rect 226103 111218 226145 111454
rect 226381 111218 226423 111454
rect 226103 111134 226423 111218
rect 226103 110898 226145 111134
rect 226381 110898 226423 111134
rect 226103 110866 226423 110898
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 214419 103596 214485 103597
rect 214419 103532 214420 103596
rect 214484 103532 214485 103596
rect 214419 103531 214485 103532
rect 213867 101148 213933 101149
rect 213867 101084 213868 101148
rect 213932 101084 213933 101148
rect 213867 101083 213933 101084
rect 213870 94893 213930 101083
rect 213867 94892 213933 94893
rect 213867 94828 213868 94892
rect 213932 94828 213933 94892
rect 213867 94827 213933 94828
rect 214422 94757 214482 103531
rect 214419 94756 214485 94757
rect 214419 94692 214420 94756
rect 214484 94692 214485 94756
rect 214419 94691 214485 94692
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 205174 240134 238182
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 242942 149157 243002 238710
rect 243234 208894 243854 238182
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 242939 149156 243005 149157
rect 242939 149092 242940 149156
rect 243004 149092 243005 149156
rect 242939 149091 243005 149092
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 136894 243854 172338
rect 244046 162485 244106 252451
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 244043 162484 244109 162485
rect 244043 162420 244044 162484
rect 244108 162420 244109 162484
rect 244043 162419 244109 162420
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 178000 272414 200898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 278819 284476 278885 284477
rect 278819 284412 278820 284476
rect 278884 284412 278885 284476
rect 278819 284411 278885 284412
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 178000 276134 204618
rect 278822 176490 278882 284411
rect 279234 280894 279854 316338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 280659 286108 280725 286109
rect 280659 286044 280660 286108
rect 280724 286044 280725 286108
rect 280659 286043 280725 286044
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279003 237964 279069 237965
rect 279003 237900 279004 237964
rect 279068 237900 279069 237964
rect 279003 237899 279069 237900
rect 279006 177170 279066 237899
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 178000 279854 208338
rect 279739 177580 279805 177581
rect 279739 177516 279740 177580
rect 279804 177516 279805 177580
rect 279739 177515 279805 177516
rect 279006 177110 279618 177170
rect 278822 176430 279434 176490
rect 268331 174588 268397 174589
rect 268331 174524 268332 174588
rect 268396 174524 268397 174588
rect 268331 174523 268397 174524
rect 267779 174452 267845 174453
rect 267779 174388 267780 174452
rect 267844 174450 267845 174452
rect 268334 174450 268394 174523
rect 267844 174390 268394 174450
rect 267844 174388 267845 174390
rect 267779 174387 267845 174388
rect 279374 172141 279434 176430
rect 279371 172140 279437 172141
rect 279371 172076 279372 172140
rect 279436 172076 279437 172140
rect 279371 172075 279437 172076
rect 279558 169829 279618 177110
rect 279742 175269 279802 177515
rect 280291 177308 280357 177309
rect 280291 177244 280292 177308
rect 280356 177244 280357 177308
rect 280291 177243 280357 177244
rect 279739 175268 279805 175269
rect 279739 175204 279740 175268
rect 279804 175204 279805 175268
rect 279739 175203 279805 175204
rect 279555 169828 279621 169829
rect 279555 169764 279556 169828
rect 279620 169764 279621 169828
rect 279555 169763 279621 169764
rect 272207 165454 272527 165486
rect 272207 165218 272249 165454
rect 272485 165218 272527 165454
rect 272207 165134 272527 165218
rect 272207 164898 272249 165134
rect 272485 164898 272527 165134
rect 272207 164866 272527 164898
rect 275471 165454 275791 165486
rect 275471 165218 275513 165454
rect 275749 165218 275791 165454
rect 275471 165134 275791 165218
rect 275471 164898 275513 165134
rect 275749 164898 275791 165134
rect 275471 164866 275791 164898
rect 268515 163028 268581 163029
rect 268515 162964 268516 163028
rect 268580 162964 268581 163028
rect 268515 162963 268581 162964
rect 268518 159901 268578 162963
rect 268515 159900 268581 159901
rect 268515 159836 268516 159900
rect 268580 159836 268581 159900
rect 268515 159835 268581 159836
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 268515 153508 268581 153509
rect 268515 153444 268516 153508
rect 268580 153444 268581 153508
rect 268515 153443 268581 153444
rect 268518 153101 268578 153443
rect 268515 153100 268581 153101
rect 268515 153036 268516 153100
rect 268580 153036 268581 153100
rect 268515 153035 268581 153036
rect 268331 147932 268397 147933
rect 268331 147868 268332 147932
rect 268396 147868 268397 147932
rect 268331 147867 268397 147868
rect 268334 146165 268394 147867
rect 270575 147454 270895 147486
rect 270575 147218 270617 147454
rect 270853 147218 270895 147454
rect 270575 147134 270895 147218
rect 270575 146898 270617 147134
rect 270853 146898 270895 147134
rect 270575 146866 270895 146898
rect 273839 147454 274159 147486
rect 273839 147218 273881 147454
rect 274117 147218 274159 147454
rect 273839 147134 274159 147218
rect 273839 146898 273881 147134
rect 274117 146898 274159 147134
rect 273839 146866 274159 146898
rect 277103 147454 277423 147486
rect 277103 147218 277145 147454
rect 277381 147218 277423 147454
rect 277103 147134 277423 147218
rect 277103 146898 277145 147134
rect 277381 146898 277423 147134
rect 277103 146866 277423 146898
rect 268331 146164 268397 146165
rect 268331 146100 268332 146164
rect 268396 146100 268397 146164
rect 268331 146099 268397 146100
rect 268515 142356 268581 142357
rect 268515 142292 268516 142356
rect 268580 142292 268581 142356
rect 268515 142291 268581 142292
rect 268518 141949 268578 142291
rect 268515 141948 268581 141949
rect 268515 141884 268516 141948
rect 268580 141884 268581 141948
rect 268515 141883 268581 141884
rect 268331 136372 268397 136373
rect 268331 136370 268332 136372
rect 268150 136310 268332 136370
rect 268150 135829 268210 136310
rect 268331 136308 268332 136310
rect 268396 136308 268397 136372
rect 268331 136307 268397 136308
rect 268147 135828 268213 135829
rect 268147 135764 268148 135828
rect 268212 135764 268213 135828
rect 268147 135763 268213 135764
rect 268515 134196 268581 134197
rect 268515 134132 268516 134196
rect 268580 134132 268581 134196
rect 268515 134131 268581 134132
rect 268518 133789 268578 134131
rect 268515 133788 268581 133789
rect 268515 133724 268516 133788
rect 268580 133724 268581 133788
rect 268515 133723 268581 133724
rect 272207 129454 272527 129486
rect 272207 129218 272249 129454
rect 272485 129218 272527 129454
rect 272207 129134 272527 129218
rect 272207 128898 272249 129134
rect 272485 128898 272527 129134
rect 272207 128866 272527 128898
rect 275471 129454 275791 129486
rect 275471 129218 275513 129454
rect 275749 129218 275791 129454
rect 275471 129134 275791 129218
rect 275471 128898 275513 129134
rect 275749 128898 275791 129134
rect 275471 128866 275791 128898
rect 268515 127260 268581 127261
rect 268515 127196 268516 127260
rect 268580 127196 268581 127260
rect 268515 127195 268581 127196
rect 268518 126853 268578 127195
rect 268515 126852 268581 126853
rect 268515 126788 268516 126852
rect 268580 126788 268581 126852
rect 268515 126787 268581 126788
rect 268515 123044 268581 123045
rect 268515 122980 268516 123044
rect 268580 122980 268581 123044
rect 268515 122979 268581 122980
rect 268518 122637 268578 122979
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 268515 122636 268581 122637
rect 268515 122572 268516 122636
rect 268580 122572 268581 122636
rect 268515 122571 268581 122572
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 268515 121684 268581 121685
rect 268515 121620 268516 121684
rect 268580 121620 268581 121684
rect 268515 121619 268581 121620
rect 268518 121277 268578 121619
rect 268515 121276 268581 121277
rect 268515 121212 268516 121276
rect 268580 121212 268581 121276
rect 268515 121211 268581 121212
rect 268331 116108 268397 116109
rect 268331 116044 268332 116108
rect 268396 116044 268397 116108
rect 268331 116043 268397 116044
rect 267779 115972 267845 115973
rect 267779 115908 267780 115972
rect 267844 115970 267845 115972
rect 268334 115970 268394 116043
rect 267844 115910 268394 115970
rect 267844 115908 267845 115910
rect 267779 115907 267845 115908
rect 270575 111454 270895 111486
rect 270575 111218 270617 111454
rect 270853 111218 270895 111454
rect 270575 111134 270895 111218
rect 270575 110898 270617 111134
rect 270853 110898 270895 111134
rect 270575 110866 270895 110898
rect 273839 111454 274159 111486
rect 273839 111218 273881 111454
rect 274117 111218 274159 111454
rect 273839 111134 274159 111218
rect 273839 110898 273881 111134
rect 274117 110898 274159 111134
rect 273839 110866 274159 110898
rect 277103 111454 277423 111486
rect 277103 111218 277145 111454
rect 277381 111218 277423 111454
rect 277103 111134 277423 111218
rect 277103 110898 277145 111134
rect 277381 110898 277423 111134
rect 277103 110866 277423 110898
rect 268515 102372 268581 102373
rect 268515 102308 268516 102372
rect 268580 102308 268581 102372
rect 268515 102307 268581 102308
rect 268518 100605 268578 102307
rect 280294 100877 280354 177243
rect 280662 150517 280722 286043
rect 282954 284614 283574 320058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 285627 285972 285693 285973
rect 285627 285908 285628 285972
rect 285692 285908 285693 285972
rect 285627 285907 285693 285908
rect 284339 285700 284405 285701
rect 284339 285636 284340 285700
rect 284404 285636 284405 285700
rect 284339 285635 284405 285636
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 281579 231164 281645 231165
rect 281579 231100 281580 231164
rect 281644 231100 281645 231164
rect 281579 231099 281645 231100
rect 281582 163165 281642 231099
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 281763 186964 281829 186965
rect 281763 186900 281764 186964
rect 281828 186900 281829 186964
rect 281763 186899 281829 186900
rect 281766 166293 281826 186899
rect 282131 182884 282197 182885
rect 282131 182820 282132 182884
rect 282196 182820 282197 182884
rect 282131 182819 282197 182820
rect 281947 181388 282013 181389
rect 281947 181324 281948 181388
rect 282012 181324 282013 181388
rect 281947 181323 282013 181324
rect 281950 174045 282010 181323
rect 281947 174044 282013 174045
rect 281947 173980 281948 174044
rect 282012 173980 282013 174044
rect 281947 173979 282013 173980
rect 281763 166292 281829 166293
rect 281763 166228 281764 166292
rect 281828 166228 281829 166292
rect 281763 166227 281829 166228
rect 282134 163981 282194 182819
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282131 163980 282197 163981
rect 282131 163916 282132 163980
rect 282196 163916 282197 163980
rect 282131 163915 282197 163916
rect 281579 163164 281645 163165
rect 281579 163100 281580 163164
rect 281644 163100 281645 163164
rect 281579 163099 281645 163100
rect 280659 150516 280725 150517
rect 280659 150452 280660 150516
rect 280724 150452 280725 150516
rect 280659 150451 280725 150452
rect 282954 140614 283574 176058
rect 284342 140861 284402 285635
rect 284707 233884 284773 233885
rect 284707 233820 284708 233884
rect 284772 233820 284773 233884
rect 284707 233819 284773 233820
rect 284523 232660 284589 232661
rect 284523 232596 284524 232660
rect 284588 232596 284589 232660
rect 284523 232595 284589 232596
rect 284526 143173 284586 232595
rect 284710 144805 284770 233819
rect 284891 232524 284957 232525
rect 284891 232460 284892 232524
rect 284956 232460 284957 232524
rect 284891 232459 284957 232460
rect 284894 145485 284954 232459
rect 285630 147117 285690 285907
rect 287651 284748 287717 284749
rect 287651 284684 287652 284748
rect 287716 284684 287717 284748
rect 287651 284683 287717 284684
rect 285811 180164 285877 180165
rect 285811 180100 285812 180164
rect 285876 180100 285877 180164
rect 285811 180099 285877 180100
rect 285627 147116 285693 147117
rect 285627 147052 285628 147116
rect 285692 147052 285693 147116
rect 285627 147051 285693 147052
rect 284891 145484 284957 145485
rect 284891 145420 284892 145484
rect 284956 145420 284957 145484
rect 284891 145419 284957 145420
rect 284707 144804 284773 144805
rect 284707 144740 284708 144804
rect 284772 144740 284773 144804
rect 284707 144739 284773 144740
rect 284523 143172 284589 143173
rect 284523 143108 284524 143172
rect 284588 143108 284589 143172
rect 284523 143107 284589 143108
rect 284339 140860 284405 140861
rect 284339 140796 284340 140860
rect 284404 140796 284405 140860
rect 284339 140795 284405 140796
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 285814 115565 285874 180099
rect 285811 115564 285877 115565
rect 285811 115500 285812 115564
rect 285876 115500 285877 115564
rect 285811 115499 285877 115500
rect 287654 111893 287714 284683
rect 288939 277540 289005 277541
rect 288939 277476 288940 277540
rect 289004 277476 289005 277540
rect 288939 277475 289005 277476
rect 288942 151877 289002 277475
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 288939 151876 289005 151877
rect 288939 151812 288940 151876
rect 289004 151812 289005 151876
rect 288939 151811 289005 151812
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 287651 111892 287717 111893
rect 287651 111828 287652 111892
rect 287716 111828 287717 111892
rect 287651 111827 287717 111828
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 280291 100876 280357 100877
rect 280291 100812 280292 100876
rect 280356 100812 280357 100876
rect 280291 100811 280357 100812
rect 268515 100604 268581 100605
rect 268515 100540 268516 100604
rect 268580 100540 268581 100604
rect 268515 100539 268581 100540
rect 268331 97204 268397 97205
rect 268331 97140 268332 97204
rect 268396 97140 268397 97204
rect 268331 97139 268397 97140
rect 267779 96932 267845 96933
rect 267779 96868 267780 96932
rect 267844 96930 267845 96932
rect 268334 96930 268394 97139
rect 267844 96870 268394 96930
rect 267844 96868 267845 96870
rect 267779 96867 267845 96868
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 93454 272414 94000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 94000
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 94000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 219810 273218 220046 273454
rect 219810 272898 220046 273134
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 204450 255218 204686 255454
rect 204450 254898 204686 255134
rect 235170 255218 235406 255454
rect 235170 254898 235406 255134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 221249 165218 221485 165454
rect 221249 164898 221485 165134
rect 224513 165218 224749 165454
rect 224513 164898 224749 165134
rect 219617 147218 219853 147454
rect 219617 146898 219853 147134
rect 222881 147218 223117 147454
rect 222881 146898 223117 147134
rect 226145 147218 226381 147454
rect 226145 146898 226381 147134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 221249 129218 221485 129454
rect 221249 128898 221485 129134
rect 224513 129218 224749 129454
rect 224513 128898 224749 129134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 219617 111218 219853 111454
rect 219617 110898 219853 111134
rect 222881 111218 223117 111454
rect 222881 110898 223117 111134
rect 226145 111218 226381 111454
rect 226145 110898 226381 111134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 272249 165218 272485 165454
rect 272249 164898 272485 165134
rect 275513 165218 275749 165454
rect 275513 164898 275749 165134
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 270617 147218 270853 147454
rect 270617 146898 270853 147134
rect 273881 147218 274117 147454
rect 273881 146898 274117 147134
rect 277145 147218 277381 147454
rect 277145 146898 277381 147134
rect 272249 129218 272485 129454
rect 272249 128898 272485 129134
rect 275513 129218 275749 129454
rect 275513 128898 275749 129134
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 270617 111218 270853 111454
rect 270617 110898 270853 111134
rect 273881 111218 274117 111454
rect 273881 110898 274117 111134
rect 277145 111218 277381 111454
rect 277145 110898 277381 111134
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219810 273454
rect 220046 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219810 273134
rect 220046 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204450 255454
rect 204686 255218 235170 255454
rect 235406 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204450 255134
rect 204686 254898 235170 255134
rect 235406 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 221249 165454
rect 221485 165218 224513 165454
rect 224749 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 272249 165454
rect 272485 165218 275513 165454
rect 275749 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 221249 165134
rect 221485 164898 224513 165134
rect 224749 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 272249 165134
rect 272485 164898 275513 165134
rect 275749 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 219617 147454
rect 219853 147218 222881 147454
rect 223117 147218 226145 147454
rect 226381 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 270617 147454
rect 270853 147218 273881 147454
rect 274117 147218 277145 147454
rect 277381 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 219617 147134
rect 219853 146898 222881 147134
rect 223117 146898 226145 147134
rect 226381 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 270617 147134
rect 270853 146898 273881 147134
rect 274117 146898 277145 147134
rect 277381 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 221249 129454
rect 221485 129218 224513 129454
rect 224749 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 272249 129454
rect 272485 129218 275513 129454
rect 275749 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 221249 129134
rect 221485 128898 224513 129134
rect 224749 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 272249 129134
rect 272485 128898 275513 129134
rect 275749 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 219617 111454
rect 219853 111218 222881 111454
rect 223117 111218 226145 111454
rect 226381 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 270617 111454
rect 270853 111218 273881 111454
rect 274117 111218 277145 111454
rect 277381 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 219617 111134
rect 219853 110898 222881 111134
rect 223117 110898 226145 111134
rect 226381 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 270617 111134
rect 270853 110898 273881 111134
rect 274117 110898 277145 111134
rect 277381 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 268000 0 1 96000
box 0 0 12000 79688
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 12000 79688
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 200200 0 1 240182
box 0 0 44000 44000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 238182 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 286182 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 238182 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 286182 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 238182 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 286182 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 238182 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 286182 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 286182 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 286182 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 178000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 238182 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 286182 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 286182 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 286182 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 178000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 286182 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 286182 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 178000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
