magic
tech sky130A
magscale 1 2
timestamp 1647532009
<< metal1 >>
rect 201494 703264 201500 703316
rect 201552 703304 201558 703316
rect 202782 703304 202788 703316
rect 201552 703276 202788 703304
rect 201552 703264 201558 703276
rect 202782 703264 202788 703276
rect 202840 703264 202846 703316
rect 77938 703196 77944 703248
rect 77996 703236 78002 703248
rect 267642 703236 267648 703248
rect 77996 703208 267648 703236
rect 77996 703196 78002 703208
rect 267642 703196 267648 703208
rect 267700 703196 267706 703248
rect 95142 703128 95148 703180
rect 95200 703168 95206 703180
rect 332502 703168 332508 703180
rect 95200 703140 332508 703168
rect 95200 703128 95206 703140
rect 332502 703128 332508 703140
rect 332560 703128 332566 703180
rect 110322 703060 110328 703112
rect 110380 703100 110386 703112
rect 348786 703100 348792 703112
rect 110380 703072 348792 703100
rect 110380 703060 110386 703072
rect 348786 703060 348792 703072
rect 348844 703060 348850 703112
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 76558 702992 76564 703044
rect 76616 703032 76622 703044
rect 364978 703032 364984 703044
rect 76616 703004 364984 703032
rect 76616 702992 76622 703004
rect 364978 702992 364984 703004
rect 365036 702992 365042 703044
rect 104802 702924 104808 702976
rect 104860 702964 104866 702976
rect 413646 702964 413652 702976
rect 104860 702936 413652 702964
rect 104860 702924 104866 702936
rect 413646 702924 413652 702936
rect 413704 702924 413710 702976
rect 111702 702856 111708 702908
rect 111760 702896 111766 702908
rect 462314 702896 462320 702908
rect 111760 702868 462320 702896
rect 111760 702856 111766 702868
rect 462314 702856 462320 702868
rect 462372 702856 462378 702908
rect 75178 702788 75184 702840
rect 75236 702828 75242 702840
rect 381538 702828 381544 702840
rect 75236 702800 381544 702828
rect 75236 702788 75242 702800
rect 381538 702788 381544 702800
rect 381596 702828 381602 702840
rect 386414 702828 386420 702840
rect 381596 702800 386420 702828
rect 381596 702788 381602 702800
rect 386414 702788 386420 702800
rect 386472 702788 386478 702840
rect 424962 702788 424968 702840
rect 425020 702828 425026 702840
rect 429838 702828 429844 702840
rect 425020 702800 429844 702828
rect 425020 702788 425026 702800
rect 429838 702788 429844 702800
rect 429896 702788 429902 702840
rect 117222 702720 117228 702772
rect 117280 702760 117286 702772
rect 478506 702760 478512 702772
rect 117280 702732 478512 702760
rect 117280 702720 117286 702732
rect 478506 702720 478512 702732
rect 478564 702720 478570 702772
rect 113082 702652 113088 702704
rect 113140 702692 113146 702704
rect 494790 702692 494796 702704
rect 113140 702664 494796 702692
rect 113140 702652 113146 702664
rect 494790 702652 494796 702664
rect 494848 702652 494854 702704
rect 79318 702584 79324 702636
rect 79376 702624 79382 702636
rect 527174 702624 527180 702636
rect 79376 702596 527180 702624
rect 79376 702584 79382 702596
rect 527174 702584 527180 702596
rect 527232 702584 527238 702636
rect 108942 702516 108948 702568
rect 109000 702556 109006 702568
rect 465718 702556 465724 702568
rect 109000 702528 465724 702556
rect 109000 702516 109006 702528
rect 465718 702516 465724 702528
rect 465776 702516 465782 702568
rect 550542 702516 550548 702568
rect 550600 702556 550606 702568
rect 559650 702556 559656 702568
rect 550600 702528 559656 702556
rect 550600 702516 550606 702528
rect 559650 702516 559656 702528
rect 559708 702516 559714 702568
rect 68922 702448 68928 702500
rect 68980 702488 68986 702500
rect 543458 702488 543464 702500
rect 68980 702460 543464 702488
rect 68980 702448 68986 702460
rect 543458 702448 543464 702460
rect 543516 702448 543522 702500
rect 69658 700340 69664 700392
rect 69716 700380 69722 700392
rect 154114 700380 154120 700392
rect 69716 700352 154120 700380
rect 69716 700340 69722 700352
rect 154114 700340 154120 700352
rect 154172 700340 154178 700392
rect 155218 700340 155224 700392
rect 155276 700380 155282 700392
rect 218974 700380 218980 700392
rect 155276 700352 218980 700380
rect 155276 700340 155282 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 62022 700272 62028 700324
rect 62080 700312 62086 700324
rect 235166 700312 235172 700324
rect 62080 700284 235172 700312
rect 62080 700272 62086 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 238018 700272 238024 700324
rect 238076 700312 238082 700324
rect 283834 700312 283840 700324
rect 238076 700284 283840 700312
rect 238076 700272 238082 700284
rect 283834 700272 283840 700284
rect 283892 700272 283898 700324
rect 386414 700272 386420 700324
rect 386472 700312 386478 700324
rect 424962 700312 424968 700324
rect 386472 700284 424968 700312
rect 386472 700272 386478 700284
rect 424962 700272 424968 700284
rect 425020 700272 425026 700324
rect 465718 700272 465724 700324
rect 465776 700312 465782 700324
rect 550542 700312 550548 700324
rect 465776 700284 550548 700312
rect 465776 700272 465782 700284
rect 550542 700272 550548 700284
rect 550600 700272 550606 700324
rect 24302 698912 24308 698964
rect 24360 698952 24366 698964
rect 106274 698952 106280 698964
rect 24360 698924 106280 698952
rect 24360 698912 24366 698924
rect 106274 698912 106280 698924
rect 106332 698912 106338 698964
rect 159358 683136 159364 683188
rect 159416 683176 159422 683188
rect 579614 683176 579620 683188
rect 159416 683148 579620 683176
rect 159416 683136 159422 683148
rect 579614 683136 579620 683148
rect 579672 683136 579678 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 54478 670732 54484 670744
rect 3568 670704 54484 670732
rect 3568 670692 3574 670704
rect 54478 670692 54484 670704
rect 54536 670692 54542 670744
rect 90358 670692 90364 670744
rect 90416 670732 90422 670744
rect 579614 670732 579620 670744
rect 90416 670704 579620 670732
rect 90416 670692 90422 670704
rect 579614 670692 579620 670704
rect 579672 670732 579678 670744
rect 579982 670732 579988 670744
rect 579672 670704 579988 670732
rect 579672 670692 579678 670704
rect 579982 670692 579988 670704
rect 580040 670692 580046 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 11698 656928 11704 656940
rect 3568 656900 11704 656928
rect 3568 656888 3574 656900
rect 11698 656888 11704 656900
rect 11756 656888 11762 656940
rect 457438 643696 457444 643748
rect 457496 643736 457502 643748
rect 579614 643736 579620 643748
rect 457496 643708 579620 643736
rect 457496 643696 457502 643708
rect 579614 643696 579620 643708
rect 579672 643696 579678 643748
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 130378 630640 130384 630692
rect 130436 630680 130442 630692
rect 580166 630680 580172 630692
rect 130436 630652 580172 630680
rect 130436 630640 130442 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 86954 618304 86960 618316
rect 3568 618276 86960 618304
rect 3568 618264 3574 618276
rect 86954 618264 86960 618276
rect 87012 618264 87018 618316
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 35158 605860 35164 605872
rect 3568 605832 35164 605860
rect 3568 605820 3574 605832
rect 35158 605820 35164 605832
rect 35216 605820 35222 605872
rect 6914 598204 6920 598256
rect 6972 598244 6978 598256
rect 52362 598244 52368 598256
rect 6972 598216 52368 598244
rect 6972 598204 6978 598216
rect 52362 598204 52368 598216
rect 52420 598204 52426 598256
rect 52362 597524 52368 597576
rect 52420 597564 52426 597576
rect 85574 597564 85580 597576
rect 52420 597536 85580 597564
rect 52420 597524 52426 597536
rect 85574 597524 85580 597536
rect 85632 597524 85638 597576
rect 68738 596776 68744 596828
rect 68796 596816 68802 596828
rect 136634 596816 136640 596828
rect 68796 596788 136640 596816
rect 68796 596776 68802 596788
rect 136634 596776 136640 596788
rect 136692 596776 136698 596828
rect 3418 595416 3424 595468
rect 3476 595456 3482 595468
rect 42794 595456 42800 595468
rect 3476 595428 42800 595456
rect 3476 595416 3482 595428
rect 42794 595416 42800 595428
rect 42852 595416 42858 595468
rect 42794 594804 42800 594856
rect 42852 594844 42858 594856
rect 44082 594844 44088 594856
rect 42852 594816 44088 594844
rect 42852 594804 42858 594816
rect 44082 594804 44088 594816
rect 44140 594844 44146 594856
rect 71866 594844 71872 594856
rect 44140 594816 71872 594844
rect 44140 594804 44146 594816
rect 71866 594804 71872 594816
rect 71924 594804 71930 594856
rect 69014 594056 69020 594108
rect 69072 594096 69078 594108
rect 580258 594096 580264 594108
rect 69072 594068 580264 594096
rect 69072 594056 69078 594068
rect 580258 594056 580264 594068
rect 580316 594056 580322 594108
rect 81802 591268 81808 591320
rect 81860 591308 81866 591320
rect 90358 591308 90364 591320
rect 81860 591280 90364 591308
rect 81860 591268 81866 591280
rect 90358 591268 90364 591280
rect 90416 591268 90422 591320
rect 40034 590656 40040 590708
rect 40092 590696 40098 590708
rect 48222 590696 48228 590708
rect 40092 590668 48228 590696
rect 40092 590656 40098 590668
rect 48222 590656 48228 590668
rect 48280 590696 48286 590708
rect 74626 590696 74632 590708
rect 48280 590668 74632 590696
rect 48280 590656 48286 590668
rect 74626 590656 74632 590668
rect 74684 590656 74690 590708
rect 556798 590656 556804 590708
rect 556856 590696 556862 590708
rect 580166 590696 580172 590708
rect 556856 590668 580172 590696
rect 556856 590656 556862 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 91462 589296 91468 589348
rect 91520 589336 91526 589348
rect 124214 589336 124220 589348
rect 91520 589308 124220 589336
rect 91520 589296 91526 589308
rect 124214 589296 124220 589308
rect 124272 589296 124278 589348
rect 86954 588956 86960 589008
rect 87012 588996 87018 589008
rect 88242 588996 88248 589008
rect 87012 588968 88248 588996
rect 87012 588956 87018 588968
rect 88242 588956 88248 588968
rect 88300 588956 88306 589008
rect 11698 588548 11704 588600
rect 11756 588588 11762 588600
rect 87690 588588 87696 588600
rect 11756 588560 87696 588588
rect 11756 588548 11762 588560
rect 87690 588548 87696 588560
rect 87748 588548 87754 588600
rect 88334 588548 88340 588600
rect 88392 588588 88398 588600
rect 116118 588588 116124 588600
rect 88392 588560 116124 588588
rect 88392 588548 88398 588560
rect 116118 588548 116124 588560
rect 116176 588548 116182 588600
rect 56410 587868 56416 587920
rect 56468 587908 56474 587920
rect 86954 587908 86960 587920
rect 56468 587880 86960 587908
rect 56468 587868 56474 587880
rect 86954 587868 86960 587880
rect 87012 587868 87018 587920
rect 121454 587120 121460 587172
rect 121512 587160 121518 587172
rect 155218 587160 155224 587172
rect 121512 587132 155224 587160
rect 121512 587120 121518 587132
rect 155218 587120 155224 587132
rect 155276 587120 155282 587172
rect 59170 586644 59176 586696
rect 59228 586684 59234 586696
rect 83182 586684 83188 586696
rect 59228 586656 83188 586684
rect 59228 586644 59234 586656
rect 83182 586644 83188 586656
rect 83240 586644 83246 586696
rect 94866 586644 94872 586696
rect 94924 586684 94930 586696
rect 125594 586684 125600 586696
rect 94924 586656 125600 586684
rect 94924 586644 94930 586656
rect 125594 586644 125600 586656
rect 125652 586644 125658 586696
rect 39758 586576 39764 586628
rect 39816 586616 39822 586628
rect 79318 586616 79324 586628
rect 39816 586588 79324 586616
rect 39816 586576 39822 586588
rect 79318 586576 79324 586588
rect 79376 586576 79382 586628
rect 87690 586576 87696 586628
rect 87748 586616 87754 586628
rect 120166 586616 120172 586628
rect 87748 586588 120172 586616
rect 87748 586576 87754 586588
rect 120166 586576 120172 586588
rect 120224 586576 120230 586628
rect 42610 586508 42616 586560
rect 42668 586548 42674 586560
rect 82998 586548 83004 586560
rect 42668 586520 83004 586548
rect 42668 586508 42674 586520
rect 82998 586508 83004 586520
rect 83056 586508 83062 586560
rect 85298 586508 85304 586560
rect 85356 586548 85362 586560
rect 118694 586548 118700 586560
rect 85356 586520 118700 586548
rect 85356 586508 85362 586520
rect 118694 586508 118700 586520
rect 118752 586508 118758 586560
rect 68830 585760 68836 585812
rect 68888 585800 68894 585812
rect 238018 585800 238024 585812
rect 68888 585772 238024 585800
rect 68888 585760 68894 585772
rect 238018 585760 238024 585772
rect 238076 585760 238082 585812
rect 103514 585420 103520 585472
rect 103572 585460 103578 585472
rect 104802 585460 104808 585472
rect 103572 585432 104808 585460
rect 103572 585420 103578 585432
rect 104802 585420 104808 585432
rect 104860 585460 104866 585472
rect 122834 585460 122840 585472
rect 104860 585432 122840 585460
rect 104860 585420 104866 585432
rect 122834 585420 122840 585432
rect 122892 585420 122898 585472
rect 102410 585352 102416 585404
rect 102468 585392 102474 585404
rect 121454 585392 121460 585404
rect 102468 585364 121460 585392
rect 102468 585352 102474 585364
rect 121454 585352 121460 585364
rect 121512 585352 121518 585404
rect 52270 585284 52276 585336
rect 52328 585324 52334 585336
rect 76558 585324 76564 585336
rect 52328 585296 76564 585324
rect 52328 585284 52334 585296
rect 76558 585284 76564 585296
rect 76616 585284 76622 585336
rect 95142 585284 95148 585336
rect 95200 585324 95206 585336
rect 114554 585324 114560 585336
rect 95200 585296 114560 585324
rect 95200 585284 95206 585296
rect 114554 585284 114560 585296
rect 114612 585284 114618 585336
rect 53466 585216 53472 585268
rect 53524 585256 53530 585268
rect 78030 585256 78036 585268
rect 53524 585228 78036 585256
rect 53524 585216 53530 585228
rect 78030 585216 78036 585228
rect 78088 585216 78094 585268
rect 94130 585216 94136 585268
rect 94188 585256 94194 585268
rect 116210 585256 116216 585268
rect 94188 585228 116216 585256
rect 94188 585216 94194 585228
rect 116210 585216 116216 585228
rect 116268 585216 116274 585268
rect 41138 585148 41144 585200
rect 41196 585188 41202 585200
rect 80606 585188 80612 585200
rect 41196 585160 80612 585188
rect 41196 585148 41202 585160
rect 80606 585148 80612 585160
rect 80664 585148 80670 585200
rect 89622 585148 89628 585200
rect 89680 585188 89686 585200
rect 121546 585188 121552 585200
rect 89680 585160 121552 585188
rect 89680 585148 89686 585160
rect 121546 585148 121552 585160
rect 121604 585148 121610 585200
rect 88242 585080 88248 585132
rect 88300 585120 88306 585132
rect 95418 585120 95424 585132
rect 88300 585092 95424 585120
rect 88300 585080 88306 585092
rect 95418 585080 95424 585092
rect 95476 585080 95482 585132
rect 98730 585012 98736 585064
rect 98788 585052 98794 585064
rect 102410 585052 102416 585064
rect 98788 585024 102416 585052
rect 98788 585012 98794 585024
rect 102410 585012 102416 585024
rect 102468 585012 102474 585064
rect 73338 584100 73344 584112
rect 64846 584072 73344 584100
rect 57790 583992 57796 584044
rect 57848 584032 57854 584044
rect 64846 584032 64874 584072
rect 73338 584060 73344 584072
rect 73396 584060 73402 584112
rect 102594 584060 102600 584112
rect 102652 584100 102658 584112
rect 106642 584100 106648 584112
rect 102652 584072 106648 584100
rect 102652 584060 102658 584072
rect 106642 584060 106648 584072
rect 106700 584060 106706 584112
rect 70394 584032 70400 584044
rect 57848 584004 64874 584032
rect 68388 584004 70400 584032
rect 57848 583992 57854 584004
rect 53742 583924 53748 583976
rect 53800 583964 53806 583976
rect 68388 583964 68416 584004
rect 70394 583992 70400 584004
rect 70452 583992 70458 584044
rect 77846 583992 77852 584044
rect 77904 584032 77910 584044
rect 79226 584032 79232 584044
rect 77904 584004 79232 584032
rect 77904 583992 77910 584004
rect 79226 583992 79232 584004
rect 79284 583992 79290 584044
rect 104618 583992 104624 584044
rect 104676 584032 104682 584044
rect 136634 584032 136640 584044
rect 104676 584004 136640 584032
rect 104676 583992 104682 584004
rect 136634 583992 136640 584004
rect 136692 583992 136698 584044
rect 53800 583936 68416 583964
rect 53800 583924 53806 583936
rect 68462 583924 68468 583976
rect 68520 583964 68526 583976
rect 69658 583964 69664 583976
rect 68520 583936 69664 583964
rect 68520 583924 68526 583936
rect 69658 583924 69664 583936
rect 69716 583924 69722 583976
rect 101306 583924 101312 583976
rect 101364 583964 101370 583976
rect 113358 583964 113364 583976
rect 101364 583936 113364 583964
rect 101364 583924 101370 583936
rect 113358 583924 113364 583936
rect 113416 583924 113422 583976
rect 60642 583856 60648 583908
rect 60700 583896 60706 583908
rect 81894 583896 81900 583908
rect 60700 583868 81900 583896
rect 60700 583856 60706 583868
rect 81894 583856 81900 583868
rect 81952 583856 81958 583908
rect 96522 583856 96528 583908
rect 96580 583896 96586 583908
rect 110506 583896 110512 583908
rect 96580 583868 110512 583896
rect 96580 583856 96586 583868
rect 110506 583856 110512 583868
rect 110564 583856 110570 583908
rect 45370 583788 45376 583840
rect 45428 583828 45434 583840
rect 78674 583828 78680 583840
rect 45428 583800 78680 583828
rect 45428 583788 45434 583800
rect 78674 583788 78680 583800
rect 78732 583788 78738 583840
rect 99282 583788 99288 583840
rect 99340 583828 99346 583840
rect 128354 583828 128360 583840
rect 99340 583800 128360 583828
rect 99340 583788 99346 583800
rect 128354 583788 128360 583800
rect 128412 583788 128418 583840
rect 41322 583720 41328 583772
rect 41380 583760 41386 583772
rect 77846 583760 77852 583772
rect 41380 583732 77852 583760
rect 41380 583720 41386 583732
rect 77846 583720 77852 583732
rect 77904 583720 77910 583772
rect 105538 583720 105544 583772
rect 105596 583760 105602 583772
rect 114646 583760 114652 583772
rect 105596 583732 114652 583760
rect 105596 583720 105602 583732
rect 114646 583720 114652 583732
rect 114704 583720 114710 583772
rect 59078 582972 59084 583024
rect 59136 583012 59142 583024
rect 71774 583012 71780 583024
rect 59136 582984 71780 583012
rect 59136 582972 59142 582984
rect 71774 582972 71780 582984
rect 71832 582972 71838 583024
rect 97442 582700 97448 582752
rect 97500 582740 97506 582752
rect 120258 582740 120264 582752
rect 97500 582712 120264 582740
rect 97500 582700 97506 582712
rect 120258 582700 120264 582712
rect 120316 582700 120322 582752
rect 92842 582632 92848 582684
rect 92900 582672 92906 582684
rect 117406 582672 117412 582684
rect 92900 582644 117412 582672
rect 92900 582632 92906 582644
rect 117406 582632 117412 582644
rect 117464 582632 117470 582684
rect 43990 582564 43996 582616
rect 44048 582604 44054 582616
rect 76742 582604 76748 582616
rect 44048 582576 76748 582604
rect 44048 582564 44054 582576
rect 76742 582564 76748 582576
rect 76800 582564 76806 582616
rect 90266 582564 90272 582616
rect 90324 582604 90330 582616
rect 118786 582604 118792 582616
rect 90324 582576 118792 582604
rect 90324 582564 90330 582576
rect 118786 582564 118792 582576
rect 118844 582564 118850 582616
rect 46658 582496 46664 582548
rect 46716 582536 46722 582548
rect 84470 582536 84476 582548
rect 46716 582508 84476 582536
rect 46716 582496 46722 582508
rect 84470 582496 84476 582508
rect 84528 582496 84534 582548
rect 91002 582496 91008 582548
rect 91060 582536 91066 582548
rect 122926 582536 122932 582548
rect 91060 582508 122932 582536
rect 91060 582496 91066 582508
rect 122926 582496 122932 582508
rect 122984 582496 122990 582548
rect 3418 582428 3424 582480
rect 3476 582468 3482 582480
rect 107654 582468 107660 582480
rect 3476 582440 107660 582468
rect 3476 582428 3482 582440
rect 107654 582428 107660 582440
rect 107712 582428 107718 582480
rect 69198 582360 69204 582412
rect 69256 582400 69262 582412
rect 580166 582400 580172 582412
rect 69256 582372 580172 582400
rect 69256 582360 69262 582372
rect 580166 582360 580172 582372
rect 580224 582360 580230 582412
rect 66162 581816 66168 581868
rect 66220 581856 66226 581868
rect 70946 581856 70952 581868
rect 66220 581828 70952 581856
rect 66220 581816 66226 581828
rect 70946 581816 70952 581828
rect 71004 581816 71010 581868
rect 75454 581788 75460 581800
rect 64846 581760 75460 581788
rect 37090 581272 37096 581324
rect 37148 581312 37154 581324
rect 64846 581312 64874 581760
rect 75454 581748 75460 581760
rect 75512 581748 75518 581800
rect 104434 581748 104440 581800
rect 104492 581788 104498 581800
rect 108666 581788 108672 581800
rect 104492 581760 108672 581788
rect 104492 581748 104498 581760
rect 108666 581748 108672 581760
rect 108724 581748 108730 581800
rect 68738 581680 68744 581732
rect 68796 581720 68802 581732
rect 72234 581720 72240 581732
rect 68796 581692 72240 581720
rect 68796 581680 68802 581692
rect 72234 581680 72240 581692
rect 72292 581680 72298 581732
rect 84010 581720 84016 581732
rect 74506 581692 84016 581720
rect 37148 581284 64874 581312
rect 37148 581272 37154 581284
rect 50338 581204 50344 581256
rect 50396 581244 50402 581256
rect 67634 581244 67640 581256
rect 50396 581216 67640 581244
rect 50396 581204 50402 581216
rect 67634 581204 67640 581216
rect 67692 581204 67698 581256
rect 57882 581136 57888 581188
rect 57940 581176 57946 581188
rect 74506 581176 74534 581692
rect 84010 581680 84016 581692
rect 84068 581680 84074 581732
rect 97902 581680 97908 581732
rect 97960 581720 97966 581732
rect 97960 581692 103514 581720
rect 97960 581680 97966 581692
rect 57940 581148 74534 581176
rect 57940 581136 57946 581148
rect 35802 581068 35808 581120
rect 35860 581108 35866 581120
rect 68738 581108 68744 581120
rect 35860 581080 68744 581108
rect 35860 581068 35866 581080
rect 68738 581068 68744 581080
rect 68796 581068 68802 581120
rect 103486 581040 103514 581692
rect 103882 581680 103888 581732
rect 103940 581720 103946 581732
rect 103940 581692 113174 581720
rect 103940 581680 103946 581692
rect 113146 581176 113174 581692
rect 113266 581176 113272 581188
rect 113146 581148 113272 581176
rect 113266 581136 113272 581148
rect 113324 581136 113330 581188
rect 108666 581068 108672 581120
rect 108724 581108 108730 581120
rect 128446 581108 128452 581120
rect 108724 581080 128452 581108
rect 108724 581068 108730 581080
rect 128446 581068 128452 581080
rect 128504 581068 128510 581120
rect 128630 581040 128636 581052
rect 103486 581012 128636 581040
rect 128630 581000 128636 581012
rect 128688 581000 128694 581052
rect 106642 580932 106648 580984
rect 106700 580972 106706 580984
rect 114830 580972 114836 580984
rect 106700 580944 114836 580972
rect 106700 580932 106706 580944
rect 114830 580932 114836 580944
rect 114888 580932 114894 580984
rect 39942 580252 39948 580304
rect 40000 580292 40006 580304
rect 67818 580292 67824 580304
rect 40000 580264 67824 580292
rect 40000 580252 40006 580264
rect 67818 580252 67824 580264
rect 67876 580252 67882 580304
rect 108942 579708 108948 579760
rect 109000 579748 109006 579760
rect 126974 579748 126980 579760
rect 109000 579720 126980 579748
rect 109000 579708 109006 579720
rect 126974 579708 126980 579720
rect 127032 579708 127038 579760
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 53098 579680 53104 579692
rect 3384 579652 53104 579680
rect 3384 579640 3390 579652
rect 53098 579640 53104 579652
rect 53156 579640 53162 579692
rect 69106 579028 69112 579080
rect 69164 579068 69170 579080
rect 69750 579068 69756 579080
rect 69164 579040 69756 579068
rect 69164 579028 69170 579040
rect 69750 579028 69756 579040
rect 69808 579028 69814 579080
rect 59262 578280 59268 578332
rect 59320 578320 59326 578332
rect 67634 578320 67640 578332
rect 59320 578292 67640 578320
rect 59320 578280 59326 578292
rect 67634 578280 67640 578292
rect 67692 578280 67698 578332
rect 108390 578280 108396 578332
rect 108448 578320 108454 578332
rect 111886 578320 111892 578332
rect 108448 578292 111892 578320
rect 108448 578280 108454 578292
rect 111886 578280 111892 578292
rect 111944 578280 111950 578332
rect 108942 578212 108948 578264
rect 109000 578252 109006 578264
rect 131114 578252 131120 578264
rect 109000 578224 131120 578252
rect 109000 578212 109006 578224
rect 131114 578212 131120 578224
rect 131172 578212 131178 578264
rect 108850 577464 108856 577516
rect 108908 577504 108914 577516
rect 115934 577504 115940 577516
rect 108908 577476 115940 577504
rect 108908 577464 108914 577476
rect 115934 577464 115940 577476
rect 115992 577464 115998 577516
rect 66070 577396 66076 577448
rect 66128 577436 66134 577448
rect 68186 577436 68192 577448
rect 66128 577408 68192 577436
rect 66128 577396 66134 577408
rect 68186 577396 68192 577408
rect 68244 577396 68250 577448
rect 108942 576852 108948 576904
rect 109000 576892 109006 576904
rect 138014 576892 138020 576904
rect 109000 576864 138020 576892
rect 109000 576852 109006 576864
rect 138014 576852 138020 576864
rect 138072 576852 138078 576904
rect 108942 576104 108948 576156
rect 109000 576144 109006 576156
rect 123110 576144 123116 576156
rect 109000 576116 123116 576144
rect 109000 576104 109006 576116
rect 123110 576104 123116 576116
rect 123168 576104 123174 576156
rect 38562 575492 38568 575544
rect 38620 575532 38626 575544
rect 67634 575532 67640 575544
rect 38620 575504 67640 575532
rect 38620 575492 38626 575504
rect 67634 575492 67640 575504
rect 67692 575492 67698 575544
rect 108482 575492 108488 575544
rect 108540 575532 108546 575544
rect 117314 575532 117320 575544
rect 108540 575504 117320 575532
rect 108540 575492 108546 575504
rect 117314 575492 117320 575504
rect 117372 575492 117378 575544
rect 123110 575492 123116 575544
rect 123168 575532 123174 575544
rect 429838 575532 429844 575544
rect 123168 575504 429844 575532
rect 123168 575492 123174 575504
rect 429838 575492 429844 575504
rect 429896 575492 429902 575544
rect 52178 574064 52184 574116
rect 52236 574104 52242 574116
rect 67634 574104 67640 574116
rect 52236 574076 67640 574104
rect 52236 574064 52242 574076
rect 67634 574064 67640 574076
rect 67692 574064 67698 574116
rect 126882 573996 126888 574048
rect 126940 574036 126946 574048
rect 159358 574036 159364 574048
rect 126940 574008 159364 574036
rect 126940 573996 126946 574008
rect 159358 573996 159364 574008
rect 159416 573996 159422 574048
rect 108942 573316 108948 573368
rect 109000 573356 109006 573368
rect 126146 573356 126152 573368
rect 109000 573328 126152 573356
rect 109000 573316 109006 573328
rect 126146 573316 126152 573328
rect 126204 573356 126210 573368
rect 126882 573356 126888 573368
rect 126204 573328 126888 573356
rect 126204 573316 126210 573328
rect 126882 573316 126888 573328
rect 126940 573316 126946 573368
rect 105630 572840 105636 572892
rect 105688 572880 105694 572892
rect 110598 572880 110604 572892
rect 105688 572852 110604 572880
rect 105688 572840 105694 572852
rect 110598 572840 110604 572852
rect 110656 572840 110662 572892
rect 65978 572772 65984 572824
rect 66036 572812 66042 572824
rect 67726 572812 67732 572824
rect 66036 572784 67732 572812
rect 66036 572772 66042 572784
rect 67726 572772 67732 572784
rect 67784 572772 67790 572824
rect 61930 572704 61936 572756
rect 61988 572744 61994 572756
rect 67634 572744 67640 572756
rect 61988 572716 67640 572744
rect 61988 572704 61994 572716
rect 67634 572704 67640 572716
rect 67692 572704 67698 572756
rect 107654 572704 107660 572756
rect 107712 572744 107718 572756
rect 110414 572744 110420 572756
rect 107712 572716 110420 572744
rect 107712 572704 107718 572716
rect 110414 572704 110420 572716
rect 110472 572704 110478 572756
rect 55030 572024 55036 572076
rect 55088 572064 55094 572076
rect 67818 572064 67824 572076
rect 55088 572036 67824 572064
rect 55088 572024 55094 572036
rect 67818 572024 67824 572036
rect 67876 572024 67882 572076
rect 49510 571956 49516 572008
rect 49568 571996 49574 572008
rect 67910 571996 67916 572008
rect 49568 571968 67916 571996
rect 49568 571956 49574 571968
rect 67910 571956 67916 571968
rect 67968 571956 67974 572008
rect 108942 571344 108948 571396
rect 109000 571384 109006 571396
rect 130010 571384 130016 571396
rect 109000 571356 130016 571384
rect 109000 571344 109006 571356
rect 130010 571344 130016 571356
rect 130068 571344 130074 571396
rect 66162 571276 66168 571328
rect 66220 571316 66226 571328
rect 68278 571316 68284 571328
rect 66220 571288 68284 571316
rect 66220 571276 66226 571288
rect 68278 571276 68284 571288
rect 68336 571276 68342 571328
rect 108850 569984 108856 570036
rect 108908 570024 108914 570036
rect 136726 570024 136732 570036
rect 108908 569996 136732 570024
rect 108908 569984 108914 569996
rect 136726 569984 136732 569996
rect 136784 569984 136790 570036
rect 63218 569916 63224 569968
rect 63276 569956 63282 569968
rect 67634 569956 67640 569968
rect 63276 569928 67640 569956
rect 63276 569916 63282 569928
rect 67634 569916 67640 569928
rect 67692 569916 67698 569968
rect 108942 569916 108948 569968
rect 109000 569956 109006 569968
rect 139394 569956 139400 569968
rect 109000 569928 139400 569956
rect 109000 569916 109006 569928
rect 139394 569916 139400 569928
rect 139452 569916 139458 569968
rect 66162 568624 66168 568676
rect 66220 568664 66226 568676
rect 67726 568664 67732 568676
rect 66220 568636 67732 568664
rect 66220 568624 66226 568636
rect 67726 568624 67732 568636
rect 67784 568624 67790 568676
rect 34238 568556 34244 568608
rect 34296 568596 34302 568608
rect 67634 568596 67640 568608
rect 34296 568568 67640 568596
rect 34296 568556 34302 568568
rect 67634 568556 67640 568568
rect 67692 568556 67698 568608
rect 108942 568556 108948 568608
rect 109000 568596 109006 568608
rect 124858 568596 124864 568608
rect 109000 568568 124864 568596
rect 109000 568556 109006 568568
rect 124858 568556 124864 568568
rect 124916 568556 124922 568608
rect 108942 567536 108948 567588
rect 109000 567576 109006 567588
rect 113818 567576 113824 567588
rect 109000 567548 113824 567576
rect 109000 567536 109006 567548
rect 113818 567536 113824 567548
rect 113876 567536 113882 567588
rect 64598 567264 64604 567316
rect 64656 567304 64662 567316
rect 67634 567304 67640 567316
rect 64656 567276 67640 567304
rect 64656 567264 64662 567276
rect 67634 567264 67640 567276
rect 67692 567264 67698 567316
rect 60458 567196 60464 567248
rect 60516 567236 60522 567248
rect 67726 567236 67732 567248
rect 60516 567208 67732 567236
rect 60516 567196 60522 567208
rect 67726 567196 67732 567208
rect 67784 567196 67790 567248
rect 108942 567196 108948 567248
rect 109000 567236 109006 567248
rect 117958 567236 117964 567248
rect 109000 567208 117964 567236
rect 109000 567196 109006 567208
rect 117958 567196 117964 567208
rect 118016 567196 118022 567248
rect 106918 566448 106924 566500
rect 106976 566488 106982 566500
rect 121638 566488 121644 566500
rect 106976 566460 121644 566488
rect 106976 566448 106982 566460
rect 121638 566448 121644 566460
rect 121696 566448 121702 566500
rect 108390 565904 108396 565956
rect 108448 565944 108454 565956
rect 111978 565944 111984 565956
rect 108448 565916 111984 565944
rect 108448 565904 108454 565916
rect 111978 565904 111984 565916
rect 112036 565904 112042 565956
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 25498 565876 25504 565888
rect 3292 565848 25504 565876
rect 3292 565836 3298 565848
rect 25498 565836 25504 565848
rect 25556 565836 25562 565888
rect 64690 565836 64696 565888
rect 64748 565876 64754 565888
rect 67634 565876 67640 565888
rect 64748 565848 67640 565876
rect 64748 565836 64754 565848
rect 67634 565836 67640 565848
rect 67692 565836 67698 565888
rect 108942 565836 108948 565888
rect 109000 565876 109006 565888
rect 140866 565876 140872 565888
rect 109000 565848 140872 565876
rect 109000 565836 109006 565848
rect 140866 565836 140872 565848
rect 140924 565836 140930 565888
rect 48038 564476 48044 564528
rect 48096 564516 48102 564528
rect 67634 564516 67640 564528
rect 48096 564488 67640 564516
rect 48096 564476 48102 564488
rect 67634 564476 67640 564488
rect 67692 564476 67698 564528
rect 117222 564476 117228 564528
rect 117280 564516 117286 564528
rect 132586 564516 132592 564528
rect 117280 564488 132592 564516
rect 117280 564476 117286 564488
rect 132586 564476 132592 564488
rect 132644 564476 132650 564528
rect 108942 564408 108948 564460
rect 109000 564448 109006 564460
rect 143442 564448 143448 564460
rect 109000 564420 143448 564448
rect 109000 564408 109006 564420
rect 143442 564408 143448 564420
rect 143500 564448 143506 564460
rect 204898 564448 204904 564460
rect 143500 564420 204904 564448
rect 143500 564408 143506 564420
rect 204898 564408 204904 564420
rect 204956 564408 204962 564460
rect 108390 564340 108396 564392
rect 108448 564380 108454 564392
rect 117222 564380 117228 564392
rect 108448 564352 117228 564380
rect 108448 564340 108454 564352
rect 117222 564340 117228 564352
rect 117280 564340 117286 564392
rect 374638 563660 374644 563712
rect 374696 563700 374702 563712
rect 429838 563700 429844 563712
rect 374696 563672 429844 563700
rect 374696 563660 374702 563672
rect 429838 563660 429844 563672
rect 429896 563700 429902 563712
rect 580166 563700 580172 563712
rect 429896 563672 580172 563700
rect 429896 563660 429902 563672
rect 580166 563660 580172 563672
rect 580224 563660 580230 563712
rect 63126 563116 63132 563168
rect 63184 563156 63190 563168
rect 67634 563156 67640 563168
rect 63184 563128 67640 563156
rect 63184 563116 63190 563128
rect 67634 563116 67640 563128
rect 67692 563116 67698 563168
rect 56502 563048 56508 563100
rect 56560 563088 56566 563100
rect 67726 563088 67732 563100
rect 56560 563060 67732 563088
rect 56560 563048 56566 563060
rect 67726 563048 67732 563060
rect 67784 563048 67790 563100
rect 60734 562300 60740 562352
rect 60792 562340 60798 562352
rect 62022 562340 62028 562352
rect 60792 562312 62028 562340
rect 60792 562300 60798 562312
rect 62022 562300 62028 562312
rect 62080 562340 62086 562352
rect 67634 562340 67640 562352
rect 62080 562312 67640 562340
rect 62080 562300 62086 562312
rect 67634 562300 67640 562312
rect 67692 562300 67698 562352
rect 61746 561688 61752 561740
rect 61804 561728 61810 561740
rect 67634 561728 67640 561740
rect 61804 561700 67640 561728
rect 61804 561688 61810 561700
rect 67634 561688 67640 561700
rect 67692 561688 67698 561740
rect 108942 561688 108948 561740
rect 109000 561728 109006 561740
rect 135438 561728 135444 561740
rect 109000 561700 135444 561728
rect 109000 561688 109006 561700
rect 135438 561688 135444 561700
rect 135496 561688 135502 561740
rect 53558 560940 53564 560992
rect 53616 560980 53622 560992
rect 60734 560980 60740 560992
rect 53616 560952 60740 560980
rect 53616 560940 53622 560952
rect 60734 560940 60740 560952
rect 60792 560940 60798 560992
rect 58986 560328 58992 560380
rect 59044 560368 59050 560380
rect 67726 560368 67732 560380
rect 59044 560340 67732 560368
rect 59044 560328 59050 560340
rect 67726 560328 67732 560340
rect 67784 560328 67790 560380
rect 108206 560328 108212 560380
rect 108264 560368 108270 560380
rect 131390 560368 131396 560380
rect 108264 560340 131396 560368
rect 108264 560328 108270 560340
rect 131390 560328 131396 560340
rect 131448 560328 131454 560380
rect 55122 560260 55128 560312
rect 55180 560300 55186 560312
rect 67634 560300 67640 560312
rect 55180 560272 67640 560300
rect 55180 560260 55186 560272
rect 67634 560260 67640 560272
rect 67692 560260 67698 560312
rect 108942 560260 108948 560312
rect 109000 560300 109006 560312
rect 133966 560300 133972 560312
rect 109000 560272 133972 560300
rect 109000 560260 109006 560272
rect 133966 560260 133972 560272
rect 134024 560260 134030 560312
rect 135162 559512 135168 559564
rect 135220 559552 135226 559564
rect 201494 559552 201500 559564
rect 135220 559524 201500 559552
rect 135220 559512 135226 559524
rect 201494 559512 201500 559524
rect 201552 559512 201558 559564
rect 108942 558968 108948 559020
rect 109000 559008 109006 559020
rect 132770 559008 132776 559020
rect 109000 558980 132776 559008
rect 109000 558968 109006 558980
rect 132770 558968 132776 558980
rect 132828 558968 132834 559020
rect 41230 558900 41236 558952
rect 41288 558940 41294 558952
rect 67634 558940 67640 558952
rect 41288 558912 67640 558940
rect 41288 558900 41294 558912
rect 67634 558900 67640 558912
rect 67692 558900 67698 558952
rect 108850 558900 108856 558952
rect 108908 558940 108914 558952
rect 133874 558940 133880 558952
rect 108908 558912 133880 558940
rect 108908 558900 108914 558912
rect 133874 558900 133880 558912
rect 133932 558940 133938 558952
rect 135162 558940 135168 558952
rect 133932 558912 135168 558940
rect 133932 558900 133938 558912
rect 135162 558900 135168 558912
rect 135220 558900 135226 558952
rect 64782 558220 64788 558272
rect 64840 558260 64846 558272
rect 68830 558260 68836 558272
rect 64840 558232 68836 558260
rect 64840 558220 64846 558232
rect 68830 558220 68836 558232
rect 68888 558220 68894 558272
rect 59170 558152 59176 558204
rect 59228 558192 59234 558204
rect 69750 558192 69756 558204
rect 59228 558164 69756 558192
rect 59228 558152 59234 558164
rect 69750 558152 69756 558164
rect 69808 558152 69814 558204
rect 108942 557540 108948 557592
rect 109000 557580 109006 557592
rect 116026 557580 116032 557592
rect 109000 557552 116032 557580
rect 109000 557540 109006 557552
rect 116026 557540 116032 557552
rect 116084 557540 116090 557592
rect 48130 556248 48136 556300
rect 48188 556288 48194 556300
rect 67634 556288 67640 556300
rect 48188 556260 67640 556288
rect 48188 556248 48194 556260
rect 67634 556248 67640 556260
rect 67692 556248 67698 556300
rect 42702 556180 42708 556232
rect 42760 556220 42766 556232
rect 67726 556220 67732 556232
rect 42760 556192 67732 556220
rect 42760 556180 42766 556192
rect 67726 556180 67732 556192
rect 67784 556180 67790 556232
rect 108942 556180 108948 556232
rect 109000 556220 109006 556232
rect 136818 556220 136824 556232
rect 109000 556192 136824 556220
rect 109000 556180 109006 556192
rect 136818 556180 136824 556192
rect 136876 556180 136882 556232
rect 108850 556112 108856 556164
rect 108908 556152 108914 556164
rect 110598 556152 110604 556164
rect 108908 556124 110604 556152
rect 108908 556112 108914 556124
rect 110598 556112 110604 556124
rect 110656 556112 110662 556164
rect 110598 555432 110604 555484
rect 110656 555472 110662 555484
rect 125962 555472 125968 555484
rect 110656 555444 125968 555472
rect 110656 555432 110662 555444
rect 125962 555432 125968 555444
rect 126020 555432 126026 555484
rect 57606 554820 57612 554872
rect 57664 554860 57670 554872
rect 67634 554860 67640 554872
rect 57664 554832 67640 554860
rect 57664 554820 57670 554832
rect 67634 554820 67640 554832
rect 67692 554820 67698 554872
rect 36538 554752 36544 554804
rect 36596 554792 36602 554804
rect 67726 554792 67732 554804
rect 36596 554764 67732 554792
rect 36596 554752 36602 554764
rect 67726 554752 67732 554764
rect 67784 554752 67790 554804
rect 140958 554004 140964 554056
rect 141016 554044 141022 554056
rect 556798 554044 556804 554056
rect 141016 554016 556804 554044
rect 141016 554004 141022 554016
rect 556798 554004 556804 554016
rect 556856 554004 556862 554056
rect 58618 553392 58624 553444
rect 58676 553432 58682 553444
rect 67634 553432 67640 553444
rect 58676 553404 67640 553432
rect 58676 553392 58682 553404
rect 67634 553392 67640 553404
rect 67692 553392 67698 553444
rect 108942 553392 108948 553444
rect 109000 553432 109006 553444
rect 140958 553432 140964 553444
rect 109000 553404 140964 553432
rect 109000 553392 109006 553404
rect 140958 553392 140964 553404
rect 141016 553392 141022 553444
rect 54938 552032 54944 552084
rect 54996 552072 55002 552084
rect 67634 552072 67640 552084
rect 54996 552044 67640 552072
rect 54996 552032 55002 552044
rect 67634 552032 67640 552044
rect 67692 552032 67698 552084
rect 35710 550604 35716 550656
rect 35768 550644 35774 550656
rect 67634 550644 67640 550656
rect 35768 550616 67640 550644
rect 35768 550604 35774 550616
rect 67634 550604 67640 550616
rect 67692 550604 67698 550656
rect 108942 550604 108948 550656
rect 109000 550644 109006 550656
rect 120074 550644 120080 550656
rect 109000 550616 120080 550644
rect 109000 550604 109006 550616
rect 120074 550604 120080 550616
rect 120132 550604 120138 550656
rect 63310 549312 63316 549364
rect 63368 549352 63374 549364
rect 67634 549352 67640 549364
rect 63368 549324 67640 549352
rect 63368 549312 63374 549324
rect 67634 549312 67640 549324
rect 67692 549312 67698 549364
rect 108850 549312 108856 549364
rect 108908 549352 108914 549364
rect 134242 549352 134248 549364
rect 108908 549324 134248 549352
rect 108908 549312 108914 549324
rect 134242 549312 134248 549324
rect 134300 549312 134306 549364
rect 61838 549244 61844 549296
rect 61896 549284 61902 549296
rect 67726 549284 67732 549296
rect 61896 549256 67732 549284
rect 61896 549244 61902 549256
rect 67726 549244 67732 549256
rect 67784 549244 67790 549296
rect 108942 549244 108948 549296
rect 109000 549284 109006 549296
rect 142154 549284 142160 549296
rect 109000 549256 142160 549284
rect 109000 549244 109006 549256
rect 142154 549244 142160 549256
rect 142212 549244 142218 549296
rect 34330 547884 34336 547936
rect 34388 547924 34394 547936
rect 67634 547924 67640 547936
rect 34388 547896 67640 547924
rect 34388 547884 34394 547896
rect 67634 547884 67640 547896
rect 67692 547884 67698 547936
rect 108942 547884 108948 547936
rect 109000 547924 109006 547936
rect 139578 547924 139584 547936
rect 109000 547896 139584 547924
rect 109000 547884 109006 547896
rect 139578 547884 139584 547896
rect 139636 547884 139642 547936
rect 60550 546456 60556 546508
rect 60608 546496 60614 546508
rect 67634 546496 67640 546508
rect 60608 546468 67640 546496
rect 60608 546456 60614 546468
rect 67634 546456 67640 546468
rect 67692 546456 67698 546508
rect 108942 546456 108948 546508
rect 109000 546496 109006 546508
rect 135346 546496 135352 546508
rect 109000 546468 135352 546496
rect 109000 546456 109006 546468
rect 135346 546456 135352 546468
rect 135404 546456 135410 546508
rect 108942 545708 108948 545760
rect 109000 545748 109006 545760
rect 113082 545748 113088 545760
rect 109000 545720 113088 545748
rect 109000 545708 109006 545720
rect 113082 545708 113088 545720
rect 113140 545748 113146 545760
rect 119338 545748 119344 545760
rect 113140 545720 119344 545748
rect 113140 545708 113146 545720
rect 119338 545708 119344 545720
rect 119396 545708 119402 545760
rect 108942 545096 108948 545148
rect 109000 545136 109006 545148
rect 138198 545136 138204 545148
rect 109000 545108 138204 545136
rect 109000 545096 109006 545108
rect 138198 545096 138204 545108
rect 138256 545096 138262 545148
rect 25498 544348 25504 544400
rect 25556 544388 25562 544400
rect 67726 544388 67732 544400
rect 25556 544360 67732 544388
rect 25556 544348 25562 544360
rect 67726 544348 67732 544360
rect 67784 544348 67790 544400
rect 60274 542444 60280 542496
rect 60332 542484 60338 542496
rect 67634 542484 67640 542496
rect 60332 542456 67640 542484
rect 60332 542444 60338 542456
rect 67634 542444 67640 542456
rect 67692 542444 67698 542496
rect 49602 542376 49608 542428
rect 49660 542416 49666 542428
rect 68002 542416 68008 542428
rect 49660 542388 68008 542416
rect 49660 542376 49666 542388
rect 68002 542376 68008 542388
rect 68060 542376 68066 542428
rect 108942 542376 108948 542428
rect 109000 542416 109006 542428
rect 134150 542416 134156 542428
rect 109000 542388 134156 542416
rect 109000 542376 109006 542388
rect 134150 542376 134156 542388
rect 134208 542376 134214 542428
rect 60642 541628 60648 541680
rect 60700 541668 60706 541680
rect 69658 541668 69664 541680
rect 60700 541640 69664 541668
rect 60700 541628 60706 541640
rect 69658 541628 69664 541640
rect 69716 541628 69722 541680
rect 128538 541628 128544 541680
rect 128596 541668 128602 541680
rect 299474 541668 299480 541680
rect 128596 541640 299480 541668
rect 128596 541628 128602 541640
rect 299474 541628 299480 541640
rect 299532 541628 299538 541680
rect 64138 541016 64144 541068
rect 64196 541056 64202 541068
rect 67726 541056 67732 541068
rect 64196 541028 67732 541056
rect 64196 541016 64202 541028
rect 67726 541016 67732 541028
rect 67784 541016 67790 541068
rect 63402 540948 63408 541000
rect 63460 540988 63466 541000
rect 67634 540988 67640 541000
rect 63460 540960 67640 540988
rect 63460 540948 63466 540960
rect 67634 540948 67640 540960
rect 67692 540948 67698 541000
rect 109678 540948 109684 541000
rect 109736 540988 109742 541000
rect 128538 540988 128544 541000
rect 109736 540960 128544 540988
rect 109736 540948 109742 540960
rect 128538 540948 128544 540960
rect 128596 540948 128602 541000
rect 108942 539656 108948 539708
rect 109000 539696 109006 539708
rect 110322 539696 110328 539708
rect 109000 539668 110328 539696
rect 109000 539656 109006 539668
rect 110322 539656 110328 539668
rect 110380 539696 110386 539708
rect 114738 539696 114744 539708
rect 110380 539668 114744 539696
rect 110380 539656 110386 539668
rect 114738 539656 114744 539668
rect 114796 539656 114802 539708
rect 62022 539588 62028 539640
rect 62080 539628 62086 539640
rect 67634 539628 67640 539640
rect 62080 539600 67640 539628
rect 62080 539588 62086 539600
rect 67634 539588 67640 539600
rect 67692 539588 67698 539640
rect 107838 539588 107844 539640
rect 107896 539628 107902 539640
rect 127066 539628 127072 539640
rect 107896 539600 127072 539628
rect 107896 539588 107902 539600
rect 127066 539588 127072 539600
rect 127124 539588 127130 539640
rect 35158 539520 35164 539572
rect 35216 539560 35222 539572
rect 105814 539560 105820 539572
rect 35216 539532 105820 539560
rect 35216 539520 35222 539532
rect 105814 539520 105820 539532
rect 105872 539520 105878 539572
rect 54478 538908 54484 538960
rect 54536 538948 54542 538960
rect 73154 538948 73160 538960
rect 54536 538920 73160 538948
rect 54536 538908 54542 538920
rect 73154 538908 73160 538920
rect 73212 538908 73218 538960
rect 95050 538908 95056 538960
rect 95108 538948 95114 538960
rect 109126 538948 109132 538960
rect 95108 538920 109132 538948
rect 95108 538908 95114 538920
rect 109126 538908 109132 538920
rect 109184 538908 109190 538960
rect 4798 538840 4804 538892
rect 4856 538880 4862 538892
rect 82262 538880 82268 538892
rect 4856 538852 82268 538880
rect 4856 538840 4862 538852
rect 82262 538840 82268 538852
rect 82320 538840 82326 538892
rect 95142 538840 95148 538892
rect 95200 538880 95206 538892
rect 116210 538880 116216 538892
rect 95200 538852 116216 538880
rect 95200 538840 95206 538852
rect 116210 538840 116216 538852
rect 116268 538840 116274 538892
rect 122098 538840 122104 538892
rect 122156 538880 122162 538892
rect 580350 538880 580356 538892
rect 122156 538852 580356 538880
rect 122156 538840 122162 538852
rect 580350 538840 580356 538852
rect 580408 538840 580414 538892
rect 122098 538268 122104 538280
rect 110340 538240 122104 538268
rect 53098 538160 53104 538212
rect 53156 538200 53162 538212
rect 98362 538200 98368 538212
rect 53156 538172 98368 538200
rect 53156 538160 53162 538172
rect 98362 538160 98368 538172
rect 98420 538160 98426 538212
rect 103514 538160 103520 538212
rect 103572 538200 103578 538212
rect 109678 538200 109684 538212
rect 103572 538172 109684 538200
rect 103572 538160 103578 538172
rect 109678 538160 109684 538172
rect 109736 538160 109742 538212
rect 88058 538092 88064 538144
rect 88116 538132 88122 538144
rect 110340 538132 110368 538240
rect 122098 538228 122104 538240
rect 122156 538228 122162 538280
rect 204898 538160 204904 538212
rect 204956 538200 204962 538212
rect 580166 538200 580172 538212
rect 204956 538172 580172 538200
rect 204956 538160 204962 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 88116 538104 110368 538132
rect 88116 538092 88122 538104
rect 73154 538024 73160 538076
rect 73212 538064 73218 538076
rect 91278 538064 91284 538076
rect 73212 538036 91284 538064
rect 73212 538024 73218 538036
rect 91278 538024 91284 538036
rect 91336 538024 91342 538076
rect 82262 537956 82268 538008
rect 82320 537996 82326 538008
rect 99006 537996 99012 538008
rect 82320 537968 99012 537996
rect 82320 537956 82326 537968
rect 99006 537956 99012 537968
rect 99064 537956 99070 538008
rect 57882 537752 57888 537804
rect 57940 537792 57946 537804
rect 79318 537792 79324 537804
rect 57940 537764 79324 537792
rect 57940 537752 57946 537764
rect 79318 537752 79324 537764
rect 79376 537752 79382 537804
rect 94498 537684 94504 537736
rect 94556 537724 94562 537736
rect 104710 537724 104716 537736
rect 94556 537696 104716 537724
rect 94556 537684 94562 537696
rect 104710 537684 104716 537696
rect 104768 537684 104774 537736
rect 57882 537616 57888 537668
rect 57940 537656 57946 537668
rect 81618 537656 81624 537668
rect 57940 537628 81624 537656
rect 57940 537616 57946 537628
rect 81618 537616 81624 537628
rect 81676 537616 81682 537668
rect 95786 537616 95792 537668
rect 95844 537656 95850 537668
rect 123018 537656 123024 537668
rect 95844 537628 123024 537656
rect 95844 537616 95850 537628
rect 123018 537616 123024 537628
rect 123076 537616 123082 537668
rect 43806 537548 43812 537600
rect 43864 537588 43870 537600
rect 72602 537588 72608 537600
rect 43864 537560 72608 537588
rect 43864 537548 43870 537560
rect 72602 537548 72608 537560
rect 72660 537548 72666 537600
rect 102226 537548 102232 537600
rect 102284 537588 102290 537600
rect 129826 537588 129832 537600
rect 102284 537560 129832 537588
rect 102284 537548 102290 537560
rect 129826 537548 129832 537560
rect 129884 537548 129890 537600
rect 50982 537480 50988 537532
rect 51040 537520 51046 537532
rect 82906 537520 82912 537532
rect 51040 537492 82912 537520
rect 51040 537480 51046 537492
rect 82906 537480 82912 537492
rect 82964 537480 82970 537532
rect 102870 537480 102876 537532
rect 102928 537520 102934 537532
rect 132678 537520 132684 537532
rect 102928 537492 132684 537520
rect 102928 537480 102934 537492
rect 132678 537480 132684 537492
rect 132736 537480 132742 537532
rect 73154 536868 73160 536920
rect 73212 536908 73218 536920
rect 73798 536908 73804 536920
rect 73212 536880 73804 536908
rect 73212 536868 73218 536880
rect 73798 536868 73804 536880
rect 73856 536868 73862 536920
rect 84838 536868 84844 536920
rect 84896 536908 84902 536920
rect 90358 536908 90364 536920
rect 84896 536880 90364 536908
rect 84896 536868 84902 536880
rect 90358 536868 90364 536880
rect 90416 536868 90422 536920
rect 70118 536800 70124 536852
rect 70176 536840 70182 536852
rect 75914 536840 75920 536852
rect 70176 536812 75920 536840
rect 70176 536800 70182 536812
rect 75914 536800 75920 536812
rect 75972 536800 75978 536852
rect 82262 536800 82268 536852
rect 82320 536840 82326 536852
rect 82722 536840 82728 536852
rect 82320 536812 82728 536840
rect 82320 536800 82326 536812
rect 82722 536800 82728 536812
rect 82780 536800 82786 536852
rect 84102 536800 84108 536852
rect 84160 536840 84166 536852
rect 85482 536840 85488 536852
rect 84160 536812 85488 536840
rect 84160 536800 84166 536812
rect 85482 536800 85488 536812
rect 85540 536800 85546 536852
rect 102042 536800 102048 536852
rect 102100 536840 102106 536852
rect 105538 536840 105544 536852
rect 102100 536812 105544 536840
rect 102100 536800 102106 536812
rect 105538 536800 105544 536812
rect 105596 536800 105602 536852
rect 59078 536732 59084 536784
rect 59136 536772 59142 536784
rect 73890 536772 73896 536784
rect 59136 536744 73896 536772
rect 59136 536732 59142 536744
rect 73890 536732 73896 536744
rect 73948 536732 73954 536784
rect 57606 536188 57612 536240
rect 57664 536228 57670 536240
rect 65886 536228 65892 536240
rect 57664 536200 65892 536228
rect 57664 536188 57670 536200
rect 65886 536188 65892 536200
rect 65944 536188 65950 536240
rect 45462 536120 45468 536172
rect 45520 536160 45526 536172
rect 59078 536160 59084 536172
rect 45520 536132 59084 536160
rect 45520 536120 45526 536132
rect 59078 536120 59084 536132
rect 59136 536120 59142 536172
rect 104710 536120 104716 536172
rect 104768 536160 104774 536172
rect 109126 536160 109132 536172
rect 104768 536132 109132 536160
rect 104768 536120 104774 536132
rect 109126 536120 109132 536132
rect 109184 536160 109190 536172
rect 116118 536160 116124 536172
rect 109184 536132 116124 536160
rect 109184 536120 109190 536132
rect 116118 536120 116124 536132
rect 116176 536120 116182 536172
rect 37182 536052 37188 536104
rect 37240 536092 37246 536104
rect 71314 536092 71320 536104
rect 37240 536064 71320 536092
rect 37240 536052 37246 536064
rect 71314 536052 71320 536064
rect 71372 536052 71378 536104
rect 97902 536052 97908 536104
rect 97960 536092 97966 536104
rect 114830 536092 114836 536104
rect 97960 536064 114836 536092
rect 97960 536052 97966 536064
rect 114830 536052 114836 536064
rect 114888 536052 114894 536104
rect 56318 535440 56324 535492
rect 56376 535480 56382 535492
rect 57606 535480 57612 535492
rect 56376 535452 57612 535480
rect 56376 535440 56382 535452
rect 57606 535440 57612 535452
rect 57664 535440 57670 535492
rect 65886 535372 65892 535424
rect 65944 535412 65950 535424
rect 169754 535412 169760 535424
rect 65944 535384 169760 535412
rect 65944 535372 65950 535384
rect 169754 535372 169760 535384
rect 169812 535372 169818 535424
rect 72418 534896 72424 534948
rect 72476 534936 72482 534948
rect 77754 534936 77760 534948
rect 72476 534908 77760 534936
rect 72476 534896 72482 534908
rect 77754 534896 77760 534908
rect 77812 534896 77818 534948
rect 99282 534896 99288 534948
rect 99340 534936 99346 534948
rect 113266 534936 113272 534948
rect 99340 534908 113272 534936
rect 99340 534896 99346 534908
rect 113266 534896 113272 534908
rect 113324 534896 113330 534948
rect 53650 534828 53656 534880
rect 53708 534868 53714 534880
rect 75178 534868 75184 534880
rect 53708 534840 75184 534868
rect 53708 534828 53714 534840
rect 75178 534828 75184 534840
rect 75236 534828 75242 534880
rect 98638 534828 98644 534880
rect 98696 534868 98702 534880
rect 117406 534868 117412 534880
rect 98696 534840 117412 534868
rect 98696 534828 98702 534840
rect 117406 534828 117412 534840
rect 117464 534828 117470 534880
rect 46842 534760 46848 534812
rect 46900 534800 46906 534812
rect 78398 534800 78404 534812
rect 46900 534772 78404 534800
rect 46900 534760 46906 534772
rect 78398 534760 78404 534772
rect 78456 534760 78462 534812
rect 93854 534760 93860 534812
rect 93912 534800 93918 534812
rect 125778 534800 125784 534812
rect 93912 534772 125784 534800
rect 93912 534760 93918 534772
rect 125778 534760 125784 534772
rect 125836 534760 125842 534812
rect 39850 534692 39856 534744
rect 39908 534732 39914 534744
rect 73246 534732 73252 534744
rect 39908 534704 73252 534732
rect 39908 534692 39914 534704
rect 73246 534692 73252 534704
rect 73304 534692 73310 534744
rect 89990 534692 89996 534744
rect 90048 534732 90054 534744
rect 124398 534732 124404 534744
rect 90048 534704 124404 534732
rect 90048 534692 90054 534704
rect 124398 534692 124404 534704
rect 124456 534692 124462 534744
rect 69290 533332 69296 533384
rect 69348 533372 69354 533384
rect 69750 533372 69756 533384
rect 69348 533344 69756 533372
rect 69348 533332 69354 533344
rect 69750 533332 69756 533344
rect 69808 533332 69814 533384
rect 49326 532108 49332 532160
rect 49384 532148 49390 532160
rect 76466 532148 76472 532160
rect 49384 532120 76472 532148
rect 49384 532108 49390 532120
rect 76466 532108 76472 532120
rect 76524 532108 76530 532160
rect 51994 532040 52000 532092
rect 52052 532080 52058 532092
rect 83550 532080 83556 532092
rect 52052 532052 83556 532080
rect 52052 532040 52058 532052
rect 83550 532040 83556 532052
rect 83608 532040 83614 532092
rect 89346 532040 89352 532092
rect 89404 532080 89410 532092
rect 113266 532080 113272 532092
rect 89404 532052 113272 532080
rect 89404 532040 89410 532052
rect 113266 532040 113272 532052
rect 113324 532040 113330 532092
rect 47946 531972 47952 532024
rect 48004 532012 48010 532024
rect 79042 532012 79048 532024
rect 48004 531984 79048 532012
rect 48004 531972 48010 531984
rect 79042 531972 79048 531984
rect 79100 531972 79106 532024
rect 93762 531972 93768 532024
rect 93820 532012 93826 532024
rect 124214 532012 124220 532024
rect 93820 531984 124220 532012
rect 93820 531972 93826 531984
rect 124214 531972 124220 531984
rect 124272 531972 124278 532024
rect 54846 529320 54852 529372
rect 54904 529360 54910 529372
rect 77110 529360 77116 529372
rect 54904 529332 77116 529360
rect 54904 529320 54910 529332
rect 77110 529320 77116 529332
rect 77168 529320 77174 529372
rect 41046 529252 41052 529304
rect 41104 529292 41110 529304
rect 70394 529292 70400 529304
rect 41104 529264 70400 529292
rect 41104 529252 41110 529264
rect 70394 529252 70400 529264
rect 70452 529252 70458 529304
rect 42518 529184 42524 529236
rect 42576 529224 42582 529236
rect 74534 529224 74540 529236
rect 42576 529196 74540 529224
rect 42576 529184 42582 529196
rect 74534 529184 74540 529196
rect 74592 529184 74598 529236
rect 107010 528612 107016 528624
rect 106246 528584 107016 528612
rect 3142 528504 3148 528556
rect 3200 528544 3206 528556
rect 106246 528544 106274 528584
rect 107010 528572 107016 528584
rect 107068 528612 107074 528624
rect 124950 528612 124956 528624
rect 107068 528584 124956 528612
rect 107068 528572 107074 528584
rect 124950 528572 124956 528584
rect 125008 528572 125014 528624
rect 3200 528516 106274 528544
rect 3200 528504 3206 528516
rect 39666 526396 39672 526448
rect 39724 526436 39730 526448
rect 71958 526436 71964 526448
rect 39724 526408 71964 526436
rect 39724 526396 39730 526408
rect 71958 526396 71964 526408
rect 72016 526396 72022 526448
rect 34146 525784 34152 525836
rect 34204 525824 34210 525836
rect 64138 525824 64144 525836
rect 34204 525796 64144 525824
rect 34204 525784 34210 525796
rect 64138 525784 64144 525796
rect 64196 525824 64202 525836
rect 64196 525796 64874 525824
rect 64196 525784 64202 525796
rect 64846 525756 64874 525796
rect 579798 525756 579804 525768
rect 64846 525728 579804 525756
rect 579798 525716 579804 525728
rect 579856 525716 579862 525768
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 7558 514808 7564 514820
rect 3476 514780 7564 514808
rect 3476 514768 3482 514780
rect 7558 514768 7564 514780
rect 7616 514768 7622 514820
rect 59262 511980 59268 512032
rect 59320 512020 59326 512032
rect 67450 512020 67456 512032
rect 59320 511992 67456 512020
rect 59320 511980 59326 511992
rect 67450 511980 67456 511992
rect 67508 511980 67514 512032
rect 67450 511232 67456 511284
rect 67508 511272 67514 511284
rect 405734 511272 405740 511284
rect 67508 511244 405740 511272
rect 67508 511232 67514 511244
rect 405734 511232 405740 511244
rect 405792 511232 405798 511284
rect 405734 510620 405740 510672
rect 405792 510660 405798 510672
rect 580166 510660 580172 510672
rect 405792 510632 580172 510660
rect 405792 510620 405798 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 93210 500420 93216 500472
rect 93268 500460 93274 500472
rect 116118 500460 116124 500472
rect 93268 500432 116124 500460
rect 93268 500420 93274 500432
rect 116118 500420 116124 500432
rect 116176 500420 116182 500472
rect 84102 500352 84108 500404
rect 84160 500392 84166 500404
rect 110598 500392 110604 500404
rect 84160 500364 110604 500392
rect 84160 500352 84166 500364
rect 110598 500352 110604 500364
rect 110656 500352 110662 500404
rect 91094 500284 91100 500336
rect 91152 500324 91158 500336
rect 128630 500324 128636 500336
rect 91152 500296 128636 500324
rect 91152 500284 91158 500296
rect 128630 500284 128636 500296
rect 128688 500324 128694 500336
rect 128688 500296 132494 500324
rect 128688 500284 128694 500296
rect 7558 500216 7564 500268
rect 7616 500256 7622 500268
rect 91738 500256 91744 500268
rect 7616 500228 91744 500256
rect 7616 500216 7622 500228
rect 91738 500216 91744 500228
rect 91796 500216 91802 500268
rect 91922 500216 91928 500268
rect 91980 500256 91986 500268
rect 124306 500256 124312 500268
rect 91980 500228 124312 500256
rect 91980 500216 91986 500228
rect 124306 500216 124312 500228
rect 124364 500216 124370 500268
rect 132466 500256 132494 500296
rect 135254 500256 135260 500268
rect 132466 500228 135260 500256
rect 135254 500216 135260 500228
rect 135312 500216 135318 500268
rect 84194 498788 84200 498840
rect 84252 498828 84258 498840
rect 118878 498828 118884 498840
rect 84252 498800 118884 498828
rect 84252 498788 84258 498800
rect 118878 498788 118884 498800
rect 118936 498788 118942 498840
rect 81434 498176 81440 498228
rect 81492 498216 81498 498228
rect 114922 498216 114928 498228
rect 81492 498188 114928 498216
rect 81492 498176 81498 498188
rect 114922 498176 114928 498188
rect 114980 498176 114986 498228
rect 87414 497564 87420 497616
rect 87472 497604 87478 497616
rect 112070 497604 112076 497616
rect 87472 497576 112076 497604
rect 87472 497564 87478 497576
rect 112070 497564 112076 497576
rect 112128 497564 112134 497616
rect 90634 497496 90640 497548
rect 90692 497536 90698 497548
rect 120442 497536 120448 497548
rect 90692 497508 120448 497536
rect 90692 497496 90698 497508
rect 120442 497496 120448 497508
rect 120500 497496 120506 497548
rect 69658 497428 69664 497480
rect 69716 497468 69722 497480
rect 75822 497468 75828 497480
rect 69716 497440 75828 497468
rect 69716 497428 69722 497440
rect 75822 497428 75828 497440
rect 75880 497468 75886 497480
rect 81434 497468 81440 497480
rect 75880 497440 81440 497468
rect 75880 497428 75886 497440
rect 81434 497428 81440 497440
rect 81492 497428 81498 497480
rect 83826 497428 83832 497480
rect 83884 497468 83890 497480
rect 118786 497468 118792 497480
rect 83884 497440 118792 497468
rect 83884 497428 83890 497440
rect 118786 497428 118792 497440
rect 118844 497468 118850 497480
rect 131206 497468 131212 497480
rect 118844 497440 131212 497468
rect 118844 497428 118850 497440
rect 131206 497428 131212 497440
rect 131264 497428 131270 497480
rect 88242 496136 88248 496188
rect 88300 496176 88306 496188
rect 121638 496176 121644 496188
rect 88300 496148 121644 496176
rect 88300 496136 88306 496148
rect 121638 496136 121644 496148
rect 121696 496176 121702 496188
rect 128998 496176 129004 496188
rect 121696 496148 129004 496176
rect 121696 496136 121702 496148
rect 128998 496136 129004 496148
rect 129056 496136 129062 496188
rect 50706 496068 50712 496120
rect 50764 496108 50770 496120
rect 80974 496108 80980 496120
rect 50764 496080 80980 496108
rect 50764 496068 50770 496080
rect 80974 496068 80980 496080
rect 81032 496068 81038 496120
rect 93210 496068 93216 496120
rect 93268 496108 93274 496120
rect 128354 496108 128360 496120
rect 93268 496080 128360 496108
rect 93268 496068 93274 496080
rect 128354 496068 128360 496080
rect 128412 496108 128418 496120
rect 136910 496108 136916 496120
rect 128412 496080 136916 496108
rect 128412 496068 128418 496080
rect 136910 496068 136916 496080
rect 136968 496068 136974 496120
rect 42610 495592 42616 495644
rect 42668 495632 42674 495644
rect 76098 495632 76104 495644
rect 42668 495604 76104 495632
rect 42668 495592 42674 495604
rect 76098 495592 76104 495604
rect 76156 495592 76162 495644
rect 39758 495524 39764 495576
rect 39816 495564 39822 495576
rect 73246 495564 73252 495576
rect 39816 495536 73252 495564
rect 39816 495524 39822 495536
rect 73246 495524 73252 495536
rect 73304 495524 73310 495576
rect 41138 495456 41144 495508
rect 41196 495496 41202 495508
rect 74534 495496 74540 495508
rect 41196 495468 74540 495496
rect 41196 495456 41202 495468
rect 74534 495456 74540 495468
rect 74592 495456 74598 495508
rect 3418 495388 3424 495440
rect 3476 495428 3482 495440
rect 83826 495428 83832 495440
rect 3476 495400 83832 495428
rect 3476 495388 3482 495400
rect 83826 495388 83832 495400
rect 83884 495388 83890 495440
rect 96430 494980 96436 495032
rect 96488 495020 96494 495032
rect 113174 495020 113180 495032
rect 96488 494992 113180 495020
rect 96488 494980 96494 494992
rect 113174 494980 113180 494992
rect 113232 494980 113238 495032
rect 98730 494912 98736 494964
rect 98788 494952 98794 494964
rect 121638 494952 121644 494964
rect 98788 494924 121644 494952
rect 98788 494912 98794 494924
rect 121638 494912 121644 494924
rect 121696 494912 121702 494964
rect 82262 494844 82268 494896
rect 82320 494884 82326 494896
rect 111794 494884 111800 494896
rect 82320 494856 111800 494884
rect 82320 494844 82326 494856
rect 111794 494844 111800 494856
rect 111852 494844 111858 494896
rect 82722 494776 82728 494828
rect 82780 494816 82786 494828
rect 120350 494816 120356 494828
rect 82780 494788 120356 494816
rect 82780 494776 82786 494788
rect 120350 494776 120356 494788
rect 120408 494776 120414 494828
rect 80974 494708 80980 494760
rect 81032 494748 81038 494760
rect 120166 494748 120172 494760
rect 81032 494720 120172 494748
rect 81032 494708 81038 494720
rect 120166 494708 120172 494720
rect 120224 494748 120230 494760
rect 128354 494748 128360 494760
rect 120224 494720 128360 494748
rect 120224 494708 120230 494720
rect 128354 494708 128360 494720
rect 128412 494708 128418 494760
rect 85482 494164 85488 494216
rect 85540 494204 85546 494216
rect 89622 494204 89628 494216
rect 85540 494176 89628 494204
rect 85540 494164 85546 494176
rect 89622 494164 89628 494176
rect 89680 494164 89686 494216
rect 79318 494028 79324 494080
rect 79376 494068 79382 494080
rect 79962 494068 79968 494080
rect 79376 494040 79968 494068
rect 79376 494028 79382 494040
rect 79962 494028 79968 494040
rect 80020 494068 80026 494080
rect 123110 494068 123116 494080
rect 80020 494040 123116 494068
rect 80020 494028 80026 494040
rect 123110 494028 123116 494040
rect 123168 494028 123174 494080
rect 97718 493960 97724 494012
rect 97776 494000 97782 494012
rect 102134 494000 102140 494012
rect 97776 493972 102140 494000
rect 97776 493960 97782 493972
rect 102134 493960 102140 493972
rect 102192 493960 102198 494012
rect 70854 493688 70860 493740
rect 70912 493728 70918 493740
rect 72418 493728 72424 493740
rect 70912 493700 72424 493728
rect 70912 493688 70918 493700
rect 72418 493688 72424 493700
rect 72476 493688 72482 493740
rect 95234 493484 95240 493536
rect 95292 493524 95298 493536
rect 95292 493496 113174 493524
rect 95292 493484 95298 493496
rect 81618 493416 81624 493468
rect 81676 493456 81682 493468
rect 88242 493456 88248 493468
rect 81676 493428 88248 493456
rect 81676 493416 81682 493428
rect 88242 493416 88248 493428
rect 88300 493416 88306 493468
rect 90266 493416 90272 493468
rect 90324 493456 90330 493468
rect 110506 493456 110512 493468
rect 90324 493428 110512 493456
rect 90324 493416 90330 493428
rect 110506 493416 110512 493428
rect 110564 493416 110570 493468
rect 113146 493456 113174 493496
rect 113358 493456 113364 493468
rect 113146 493428 113364 493456
rect 113358 493416 113364 493428
rect 113416 493456 113422 493468
rect 132494 493456 132500 493468
rect 113416 493428 132500 493456
rect 113416 493416 113422 493428
rect 132494 493416 132500 493428
rect 132552 493416 132558 493468
rect 57698 493348 57704 493400
rect 57756 493388 57762 493400
rect 74810 493388 74816 493400
rect 57756 493360 74816 493388
rect 57756 493348 57762 493360
rect 74810 493348 74816 493360
rect 74868 493348 74874 493400
rect 82906 493348 82912 493400
rect 82964 493388 82970 493400
rect 121546 493388 121552 493400
rect 82964 493360 121552 493388
rect 82964 493348 82970 493360
rect 121546 493348 121552 493360
rect 121604 493388 121610 493400
rect 127158 493388 127164 493400
rect 121604 493360 127164 493388
rect 121604 493348 121610 493360
rect 127158 493348 127164 493360
rect 127216 493348 127222 493400
rect 43714 493280 43720 493332
rect 43772 493320 43778 493332
rect 53466 493320 53472 493332
rect 43772 493292 53472 493320
rect 43772 493280 43778 493292
rect 53466 493280 53472 493292
rect 53524 493320 53530 493332
rect 71774 493320 71780 493332
rect 53524 493292 71780 493320
rect 53524 493280 53530 493292
rect 71774 493280 71780 493292
rect 71832 493280 71838 493332
rect 79686 493280 79692 493332
rect 79744 493320 79750 493332
rect 118694 493320 118700 493332
rect 79744 493292 118700 493320
rect 79744 493280 79750 493292
rect 118694 493280 118700 493292
rect 118752 493320 118758 493332
rect 125870 493320 125876 493332
rect 118752 493292 125876 493320
rect 118752 493280 118758 493292
rect 125870 493280 125876 493292
rect 125928 493280 125934 493332
rect 51902 492804 51908 492856
rect 51960 492844 51966 492856
rect 52270 492844 52276 492856
rect 51960 492816 52276 492844
rect 51960 492804 51966 492816
rect 52270 492804 52276 492816
rect 52328 492844 52334 492856
rect 70026 492844 70032 492856
rect 52328 492816 70032 492844
rect 52328 492804 52334 492816
rect 70026 492804 70032 492816
rect 70084 492804 70090 492856
rect 58894 492736 58900 492788
rect 58952 492776 58958 492788
rect 90266 492776 90272 492788
rect 58952 492748 90272 492776
rect 58952 492736 58958 492748
rect 90266 492736 90272 492748
rect 90324 492736 90330 492788
rect 56410 492668 56416 492720
rect 56468 492708 56474 492720
rect 89714 492708 89720 492720
rect 56468 492680 89720 492708
rect 56468 492668 56474 492680
rect 89714 492668 89720 492680
rect 89772 492668 89778 492720
rect 77754 492600 77760 492652
rect 77812 492640 77818 492652
rect 79962 492640 79968 492652
rect 77812 492612 79968 492640
rect 77812 492600 77818 492612
rect 79962 492600 79968 492612
rect 80020 492600 80026 492652
rect 91278 492600 91284 492652
rect 91336 492640 91342 492652
rect 91738 492640 91744 492652
rect 91336 492612 91744 492640
rect 91336 492600 91342 492612
rect 91738 492600 91744 492612
rect 91796 492640 91802 492652
rect 120258 492640 120264 492652
rect 91796 492612 120264 492640
rect 91796 492600 91802 492612
rect 120258 492600 120264 492612
rect 120316 492600 120322 492652
rect 120258 492328 120264 492380
rect 120316 492368 120322 492380
rect 121546 492368 121552 492380
rect 120316 492340 121552 492368
rect 120316 492328 120322 492340
rect 121546 492328 121552 492340
rect 121604 492328 121610 492380
rect 97718 492260 97724 492312
rect 97776 492300 97782 492312
rect 99282 492300 99288 492312
rect 97776 492272 99288 492300
rect 97776 492260 97782 492272
rect 99282 492260 99288 492272
rect 99340 492260 99346 492312
rect 96430 492056 96436 492108
rect 96488 492096 96494 492108
rect 97902 492096 97908 492108
rect 96488 492068 97908 492096
rect 96488 492056 96494 492068
rect 97902 492056 97908 492068
rect 97960 492056 97966 492108
rect 38470 491988 38476 492040
rect 38528 492028 38534 492040
rect 43990 492028 43996 492040
rect 38528 492000 43996 492028
rect 38528 491988 38534 492000
rect 43990 491988 43996 492000
rect 44048 492028 44054 492040
rect 70394 492028 70400 492040
rect 44048 492000 70400 492028
rect 44048 491988 44054 492000
rect 70394 491988 70400 492000
rect 70452 491988 70458 492040
rect 43898 491920 43904 491972
rect 43956 491960 43962 491972
rect 45370 491960 45376 491972
rect 43956 491932 45376 491960
rect 43956 491920 43962 491932
rect 45370 491920 45376 491932
rect 45428 491960 45434 491972
rect 72234 491960 72240 491972
rect 45428 491932 72240 491960
rect 45428 491920 45434 491932
rect 72234 491920 72240 491932
rect 72292 491920 72298 491972
rect 97920 491960 97948 492056
rect 99282 491988 99288 492040
rect 99340 492028 99346 492040
rect 111058 492028 111064 492040
rect 99340 492000 111064 492028
rect 99340 491988 99346 492000
rect 111058 491988 111064 492000
rect 111116 491988 111122 492040
rect 109770 491960 109776 491972
rect 97920 491932 109776 491960
rect 109770 491920 109776 491932
rect 109828 491920 109834 491972
rect 88702 491580 88708 491632
rect 88760 491620 88766 491632
rect 100662 491620 100668 491632
rect 88760 491592 100668 491620
rect 88760 491580 88766 491592
rect 100662 491580 100668 491592
rect 100720 491580 100726 491632
rect 84838 491512 84844 491564
rect 84896 491552 84902 491564
rect 122926 491552 122932 491564
rect 84896 491524 122932 491552
rect 84896 491512 84902 491524
rect 122926 491512 122932 491524
rect 122984 491512 122990 491564
rect 99006 491444 99012 491496
rect 99064 491484 99070 491496
rect 110506 491484 110512 491496
rect 99064 491456 110512 491484
rect 99064 491444 99070 491456
rect 110506 491444 110512 491456
rect 110564 491444 110570 491496
rect 41322 491376 41328 491428
rect 41380 491416 41386 491428
rect 41380 491388 45554 491416
rect 41380 491376 41386 491388
rect 45526 491348 45554 491388
rect 52362 491376 52368 491428
rect 52420 491416 52426 491428
rect 80054 491416 80060 491428
rect 52420 491388 80060 491416
rect 52420 491376 52426 491388
rect 80054 491376 80060 491388
rect 80112 491376 80118 491428
rect 86770 491376 86776 491428
rect 86828 491416 86834 491428
rect 86828 491388 98040 491416
rect 86828 491376 86834 491388
rect 70946 491348 70952 491360
rect 45526 491320 70952 491348
rect 70946 491308 70952 491320
rect 71004 491308 71010 491360
rect 86126 491308 86132 491360
rect 86184 491348 86190 491360
rect 93762 491348 93768 491360
rect 86184 491320 93768 491348
rect 86184 491308 86190 491320
rect 93762 491308 93768 491320
rect 93820 491308 93826 491360
rect 58618 491240 58624 491292
rect 58676 491280 58682 491292
rect 63494 491280 63500 491292
rect 58676 491252 63500 491280
rect 58676 491240 58682 491252
rect 63494 491240 63500 491252
rect 63552 491240 63558 491292
rect 98012 491280 98040 491388
rect 99650 491376 99656 491428
rect 99708 491416 99714 491428
rect 114646 491416 114652 491428
rect 99708 491388 114652 491416
rect 99708 491376 99714 491388
rect 114646 491376 114652 491388
rect 114704 491416 114710 491428
rect 115474 491416 115480 491428
rect 114704 491388 115480 491416
rect 114704 491376 114710 491388
rect 115474 491376 115480 491388
rect 115532 491376 115538 491428
rect 98638 491280 98644 491292
rect 98012 491252 98644 491280
rect 98638 491240 98644 491252
rect 98696 491280 98702 491292
rect 101398 491280 101404 491292
rect 98696 491252 101404 491280
rect 98696 491240 98702 491252
rect 101398 491240 101404 491252
rect 101456 491240 101462 491292
rect 110506 491240 110512 491292
rect 110564 491280 110570 491292
rect 111702 491280 111708 491292
rect 110564 491252 111708 491280
rect 110564 491240 110570 491252
rect 111702 491240 111708 491252
rect 111760 491280 111766 491292
rect 136634 491280 136640 491292
rect 111760 491252 136640 491280
rect 111760 491240 111766 491252
rect 136634 491240 136640 491252
rect 136692 491240 136698 491292
rect 100662 491172 100668 491224
rect 100720 491212 100726 491224
rect 114554 491212 114560 491224
rect 100720 491184 114560 491212
rect 100720 491172 100726 491184
rect 114554 491172 114560 491184
rect 114612 491172 114618 491224
rect 115474 491172 115480 491224
rect 115532 491212 115538 491224
rect 118786 491212 118792 491224
rect 115532 491184 118792 491212
rect 115532 491172 115538 491184
rect 118786 491172 118792 491184
rect 118844 491172 118850 491224
rect 59078 490764 59084 490816
rect 59136 490804 59142 490816
rect 73798 490804 73804 490816
rect 59136 490776 73804 490804
rect 59136 490764 59142 490776
rect 73798 490764 73804 490776
rect 73856 490764 73862 490816
rect 93854 490764 93860 490816
rect 93912 490804 93918 490816
rect 100018 490804 100024 490816
rect 93912 490776 100024 490804
rect 93912 490764 93918 490776
rect 100018 490764 100024 490776
rect 100076 490764 100082 490816
rect 56226 490696 56232 490748
rect 56284 490736 56290 490748
rect 79594 490736 79600 490748
rect 56284 490708 79600 490736
rect 56284 490696 56290 490708
rect 79594 490696 79600 490708
rect 79652 490696 79658 490748
rect 45370 490628 45376 490680
rect 45428 490668 45434 490680
rect 46658 490668 46664 490680
rect 45428 490640 46664 490668
rect 45428 490628 45434 490640
rect 46658 490628 46664 490640
rect 46716 490668 46722 490680
rect 78030 490668 78036 490680
rect 46716 490640 78036 490668
rect 46716 490628 46722 490640
rect 78030 490628 78036 490640
rect 78088 490628 78094 490680
rect 92842 490628 92848 490680
rect 92900 490668 92906 490680
rect 106274 490668 106280 490680
rect 92900 490640 106280 490668
rect 92900 490628 92906 490640
rect 106274 490628 106280 490640
rect 106332 490628 106338 490680
rect 35526 490560 35532 490612
rect 35584 490600 35590 490612
rect 37090 490600 37096 490612
rect 35584 490572 37096 490600
rect 35584 490560 35590 490572
rect 37090 490560 37096 490572
rect 37148 490600 37154 490612
rect 69750 490600 69756 490612
rect 37148 490572 69756 490600
rect 37148 490560 37154 490572
rect 69750 490560 69756 490572
rect 69808 490560 69814 490612
rect 94130 490560 94136 490612
rect 94188 490600 94194 490612
rect 94958 490600 94964 490612
rect 94188 490572 94964 490600
rect 94188 490560 94194 490572
rect 94958 490560 94964 490572
rect 95016 490600 95022 490612
rect 109678 490600 109684 490612
rect 95016 490572 109684 490600
rect 95016 490560 95022 490572
rect 109678 490560 109684 490572
rect 109736 490560 109742 490612
rect 114830 490560 114836 490612
rect 114888 490600 114894 490612
rect 125594 490600 125600 490612
rect 114888 490572 125600 490600
rect 114888 490560 114894 490572
rect 125594 490560 125600 490572
rect 125652 490560 125658 490612
rect 75914 490152 75920 490204
rect 75972 490192 75978 490204
rect 77064 490192 77070 490204
rect 75972 490164 77070 490192
rect 75972 490152 75978 490164
rect 77064 490152 77070 490164
rect 77122 490152 77128 490204
rect 88242 489948 88248 490000
rect 88300 489988 88306 490000
rect 114830 489988 114836 490000
rect 88300 489960 114836 489988
rect 88300 489948 88306 489960
rect 114830 489948 114836 489960
rect 114888 489948 114894 490000
rect 77294 489880 77300 489932
rect 77352 489920 77358 489932
rect 111794 489920 111800 489932
rect 77352 489892 111800 489920
rect 77352 489880 77358 489892
rect 111794 489880 111800 489892
rect 111852 489880 111858 489932
rect 69842 489812 69848 489864
rect 69900 489852 69906 489864
rect 70854 489852 70860 489864
rect 69900 489824 70860 489852
rect 69900 489812 69906 489824
rect 70854 489812 70860 489824
rect 70912 489812 70918 489864
rect 98730 489812 98736 489864
rect 98788 489852 98794 489864
rect 99282 489852 99288 489864
rect 98788 489824 99288 489852
rect 98788 489812 98794 489824
rect 99282 489812 99288 489824
rect 99340 489812 99346 489864
rect 106274 489812 106280 489864
rect 106332 489852 106338 489864
rect 107378 489852 107384 489864
rect 106332 489824 107384 489852
rect 106332 489812 106338 489824
rect 107378 489812 107384 489824
rect 107436 489852 107442 489864
rect 121454 489852 121460 489864
rect 107436 489824 121460 489852
rect 107436 489812 107442 489824
rect 121454 489812 121460 489824
rect 121512 489812 121518 489864
rect 115842 489132 115848 489184
rect 115900 489172 115906 489184
rect 126974 489172 126980 489184
rect 115900 489144 126980 489172
rect 115900 489132 115906 489144
rect 126974 489132 126980 489144
rect 127032 489132 127038 489184
rect 103422 488588 103428 488640
rect 103480 488628 103486 488640
rect 115842 488628 115848 488640
rect 103480 488600 115848 488628
rect 103480 488588 103486 488600
rect 115842 488588 115848 488600
rect 115900 488588 115906 488640
rect 99282 488520 99288 488572
rect 99340 488560 99346 488572
rect 99340 488532 113174 488560
rect 99340 488520 99346 488532
rect 103330 488452 103336 488504
rect 103388 488492 103394 488504
rect 111886 488492 111892 488504
rect 103388 488464 111892 488492
rect 103388 488452 103394 488464
rect 111886 488452 111892 488464
rect 111944 488452 111950 488504
rect 113146 488492 113174 488532
rect 122926 488520 122932 488572
rect 122984 488560 122990 488572
rect 131482 488560 131488 488572
rect 122984 488532 131488 488560
rect 122984 488520 122990 488532
rect 131482 488520 131488 488532
rect 131540 488520 131546 488572
rect 114370 488492 114376 488504
rect 113146 488464 114376 488492
rect 114370 488452 114376 488464
rect 114428 488492 114434 488504
rect 128446 488492 128452 488504
rect 114428 488464 128452 488492
rect 114428 488452 114434 488464
rect 128446 488452 128452 488464
rect 128504 488452 128510 488504
rect 102870 488384 102876 488436
rect 102928 488424 102934 488436
rect 109034 488424 109040 488436
rect 102928 488396 109040 488424
rect 102928 488384 102934 488396
rect 109034 488384 109040 488396
rect 109092 488384 109098 488436
rect 111886 487908 111892 487960
rect 111944 487948 111950 487960
rect 116210 487948 116216 487960
rect 111944 487920 116216 487948
rect 111944 487908 111950 487920
rect 116210 487908 116216 487920
rect 116268 487908 116274 487960
rect 48222 487840 48228 487892
rect 48280 487880 48286 487892
rect 57238 487880 57244 487892
rect 48280 487852 57244 487880
rect 48280 487840 48286 487852
rect 57238 487840 57244 487852
rect 57296 487840 57302 487892
rect 109034 487840 109040 487892
rect 109092 487880 109098 487892
rect 122926 487880 122932 487892
rect 109092 487852 122932 487880
rect 109092 487840 109098 487852
rect 122926 487840 122932 487852
rect 122984 487840 122990 487892
rect 50798 487772 50804 487824
rect 50856 487812 50862 487824
rect 67634 487812 67640 487824
rect 50856 487784 67640 487812
rect 50856 487772 50862 487784
rect 67634 487772 67640 487784
rect 67692 487772 67698 487824
rect 106274 487772 106280 487824
rect 106332 487812 106338 487824
rect 138014 487812 138020 487824
rect 106332 487784 138020 487812
rect 106332 487772 106338 487784
rect 138014 487772 138020 487784
rect 138072 487812 138078 487824
rect 147674 487812 147680 487824
rect 138072 487784 147680 487812
rect 138072 487772 138078 487784
rect 147674 487772 147680 487784
rect 147732 487772 147738 487824
rect 56594 487160 56600 487212
rect 56652 487200 56658 487212
rect 57238 487200 57244 487212
rect 56652 487172 57244 487200
rect 56652 487160 56658 487172
rect 57238 487160 57244 487172
rect 57296 487200 57302 487212
rect 67634 487200 67640 487212
rect 57296 487172 67640 487200
rect 57296 487160 57302 487172
rect 67634 487160 67640 487172
rect 67692 487160 67698 487212
rect 35802 487092 35808 487144
rect 35860 487132 35866 487144
rect 68094 487132 68100 487144
rect 35860 487104 68100 487132
rect 35860 487092 35866 487104
rect 68094 487092 68100 487104
rect 68152 487092 68158 487144
rect 103330 487092 103336 487144
rect 103388 487132 103394 487144
rect 131114 487132 131120 487144
rect 103388 487104 131120 487132
rect 103388 487092 103394 487104
rect 131114 487092 131120 487104
rect 131172 487132 131178 487144
rect 131298 487132 131304 487144
rect 131172 487104 131304 487132
rect 131172 487092 131178 487104
rect 131298 487092 131304 487104
rect 131356 487092 131362 487144
rect 131298 486412 131304 486464
rect 131356 486452 131362 486464
rect 142338 486452 142344 486464
rect 131356 486424 142344 486452
rect 131356 486412 131362 486424
rect 142338 486412 142344 486424
rect 142396 486412 142402 486464
rect 103422 486004 103428 486056
rect 103480 486044 103486 486056
rect 106274 486044 106280 486056
rect 103480 486016 106280 486044
rect 103480 486004 103486 486016
rect 106274 486004 106280 486016
rect 106332 486004 106338 486056
rect 65518 485840 65524 485852
rect 64846 485812 65524 485840
rect 57790 485732 57796 485784
rect 57848 485772 57854 485784
rect 64846 485772 64874 485812
rect 65518 485800 65524 485812
rect 65576 485840 65582 485852
rect 67634 485840 67640 485852
rect 65576 485812 67640 485840
rect 65576 485800 65582 485812
rect 67634 485800 67640 485812
rect 67692 485800 67698 485852
rect 57848 485744 64874 485772
rect 57848 485732 57854 485744
rect 102226 485732 102232 485784
rect 102284 485772 102290 485784
rect 115934 485772 115940 485784
rect 102284 485744 115940 485772
rect 102284 485732 102290 485744
rect 115934 485732 115940 485744
rect 115992 485772 115998 485784
rect 117222 485772 117228 485784
rect 115992 485744 117228 485772
rect 115992 485732 115998 485744
rect 117222 485732 117228 485744
rect 117280 485732 117286 485784
rect 131298 485052 131304 485104
rect 131356 485092 131362 485104
rect 131482 485092 131488 485104
rect 131356 485064 131488 485092
rect 131356 485052 131362 485064
rect 131482 485052 131488 485064
rect 131540 485052 131546 485104
rect 64506 484508 64512 484560
rect 64564 484548 64570 484560
rect 68370 484548 68376 484560
rect 64564 484520 68376 484548
rect 64564 484508 64570 484520
rect 68370 484508 68376 484520
rect 68428 484508 68434 484560
rect 53282 484412 53288 484424
rect 52472 484384 53288 484412
rect 44082 484304 44088 484356
rect 44140 484344 44146 484356
rect 52472 484344 52500 484384
rect 53282 484372 53288 484384
rect 53340 484412 53346 484424
rect 67634 484412 67640 484424
rect 53340 484384 67640 484412
rect 53340 484372 53346 484384
rect 67634 484372 67640 484384
rect 67692 484372 67698 484424
rect 102226 484372 102232 484424
rect 102284 484412 102290 484424
rect 102284 484384 113174 484412
rect 102284 484372 102290 484384
rect 113146 484356 113174 484384
rect 44140 484316 52500 484344
rect 44140 484304 44146 484316
rect 113082 484304 113088 484356
rect 113140 484344 113174 484356
rect 117314 484344 117320 484356
rect 113140 484316 117320 484344
rect 113140 484304 113146 484316
rect 117314 484304 117320 484316
rect 117372 484304 117378 484356
rect 102226 483624 102232 483676
rect 102284 483664 102290 483676
rect 123202 483664 123208 483676
rect 102284 483636 123208 483664
rect 102284 483624 102290 483636
rect 123202 483624 123208 483636
rect 123260 483624 123266 483676
rect 37090 483012 37096 483064
rect 37148 483052 37154 483064
rect 50338 483052 50344 483064
rect 37148 483024 50344 483052
rect 37148 483012 37154 483024
rect 50338 483012 50344 483024
rect 50396 483012 50402 483064
rect 104710 483012 104716 483064
rect 104768 483052 104774 483064
rect 125686 483052 125692 483064
rect 104768 483024 125692 483052
rect 104768 483012 104774 483024
rect 125686 483012 125692 483024
rect 125744 483012 125750 483064
rect 50356 482984 50384 483012
rect 67634 482984 67640 482996
rect 50356 482956 67640 482984
rect 67634 482944 67640 482956
rect 67692 482944 67698 482996
rect 102318 482944 102324 482996
rect 102376 482984 102382 482996
rect 106366 482984 106372 482996
rect 102376 482956 106372 482984
rect 102376 482944 102382 482956
rect 106366 482944 106372 482956
rect 106424 482984 106430 482996
rect 107562 482984 107568 482996
rect 106424 482956 107568 482984
rect 106424 482944 106430 482956
rect 107562 482944 107568 482956
rect 107620 482944 107626 482996
rect 115842 482944 115848 482996
rect 115900 482984 115906 482996
rect 117682 482984 117688 482996
rect 115900 482956 117688 482984
rect 115900 482944 115906 482956
rect 117682 482944 117688 482956
rect 117740 482944 117746 482996
rect 102226 482604 102232 482656
rect 102284 482644 102290 482656
rect 104710 482644 104716 482656
rect 102284 482616 104716 482644
rect 102284 482604 102290 482616
rect 104710 482604 104716 482616
rect 104768 482604 104774 482656
rect 107562 481720 107568 481772
rect 107620 481760 107626 481772
rect 115290 481760 115296 481772
rect 107620 481732 115296 481760
rect 107620 481720 107626 481732
rect 115290 481720 115296 481732
rect 115348 481720 115354 481772
rect 103486 481664 103744 481692
rect 102226 481584 102232 481636
rect 102284 481624 102290 481636
rect 103486 481624 103514 481664
rect 102284 481596 103514 481624
rect 103716 481624 103744 481664
rect 106182 481652 106188 481704
rect 106240 481692 106246 481704
rect 150618 481692 150624 481704
rect 106240 481664 150624 481692
rect 106240 481652 106246 481664
rect 150618 481652 150624 481664
rect 150676 481652 150682 481704
rect 110414 481624 110420 481636
rect 103716 481596 110420 481624
rect 102284 481584 102290 481596
rect 110414 481584 110420 481596
rect 110472 481624 110478 481636
rect 111150 481624 111156 481636
rect 110472 481596 111156 481624
rect 110472 481584 110478 481596
rect 111150 481584 111156 481596
rect 111208 481584 111214 481636
rect 102318 481516 102324 481568
rect 102376 481556 102382 481568
rect 102376 481528 103514 481556
rect 102376 481516 102382 481528
rect 103486 481488 103514 481528
rect 106182 481488 106188 481500
rect 103486 481460 106188 481488
rect 106182 481448 106188 481460
rect 106240 481448 106246 481500
rect 39942 480904 39948 480956
rect 40000 480944 40006 480956
rect 67634 480944 67640 480956
rect 40000 480916 67640 480944
rect 40000 480904 40006 480916
rect 67634 480904 67640 480916
rect 67692 480904 67698 480956
rect 101950 480904 101956 480956
rect 102008 480944 102014 480956
rect 130010 480944 130016 480956
rect 102008 480916 130016 480944
rect 102008 480904 102014 480916
rect 130010 480904 130016 480916
rect 130068 480944 130074 480956
rect 147858 480944 147864 480956
rect 130068 480916 147864 480944
rect 130068 480904 130074 480916
rect 147858 480904 147864 480916
rect 147916 480904 147922 480956
rect 59262 480224 59268 480276
rect 59320 480264 59326 480276
rect 67542 480264 67548 480276
rect 59320 480236 67548 480264
rect 59320 480224 59326 480236
rect 67542 480224 67548 480236
rect 67600 480224 67606 480276
rect 111150 480224 111156 480276
rect 111208 480264 111214 480276
rect 113358 480264 113364 480276
rect 111208 480236 113364 480264
rect 111208 480224 111214 480236
rect 113358 480224 113364 480236
rect 113416 480224 113422 480276
rect 102226 480156 102232 480208
rect 102284 480196 102290 480208
rect 104894 480196 104900 480208
rect 102284 480168 104900 480196
rect 102284 480156 102290 480168
rect 104894 480156 104900 480168
rect 104952 480156 104958 480208
rect 66070 479680 66076 479732
rect 66128 479720 66134 479732
rect 68370 479720 68376 479732
rect 66128 479692 68376 479720
rect 66128 479680 66134 479692
rect 68370 479680 68376 479692
rect 68428 479680 68434 479732
rect 124858 478864 124864 478916
rect 124916 478904 124922 478916
rect 137002 478904 137008 478916
rect 124916 478876 137008 478904
rect 124916 478864 124922 478876
rect 137002 478864 137008 478876
rect 137060 478864 137066 478916
rect 105538 477572 105544 477624
rect 105596 477612 105602 477624
rect 107930 477612 107936 477624
rect 105596 477584 107936 477612
rect 105596 477572 105602 477584
rect 107930 477572 107936 477584
rect 107988 477572 107994 477624
rect 102870 477504 102876 477556
rect 102928 477544 102934 477556
rect 111886 477544 111892 477556
rect 102928 477516 111892 477544
rect 102928 477504 102934 477516
rect 111886 477504 111892 477516
rect 111944 477504 111950 477556
rect 113818 477544 113824 477556
rect 113146 477516 113824 477544
rect 102318 477436 102324 477488
rect 102376 477476 102382 477488
rect 113146 477476 113174 477516
rect 113818 477504 113824 477516
rect 113876 477544 113882 477556
rect 118694 477544 118700 477556
rect 113876 477516 118700 477544
rect 113876 477504 113882 477516
rect 118694 477504 118700 477516
rect 118752 477504 118758 477556
rect 102376 477448 113174 477476
rect 102376 477436 102382 477448
rect 102226 477368 102232 477420
rect 102284 477408 102290 477420
rect 124858 477408 124864 477420
rect 102284 477380 124864 477408
rect 102284 477368 102290 477380
rect 124858 477368 124864 477380
rect 124916 477368 124922 477420
rect 111886 477300 111892 477352
rect 111944 477340 111950 477352
rect 113082 477340 113088 477352
rect 111944 477312 113088 477340
rect 111944 477300 111950 477312
rect 113082 477300 113088 477312
rect 113140 477340 113146 477352
rect 136726 477340 136732 477352
rect 113140 477312 136732 477340
rect 113140 477300 113146 477312
rect 136726 477300 136732 477312
rect 136784 477300 136790 477352
rect 34422 476076 34428 476128
rect 34480 476116 34486 476128
rect 67634 476116 67640 476128
rect 34480 476088 67640 476116
rect 34480 476076 34486 476088
rect 67634 476076 67640 476088
rect 67692 476076 67698 476128
rect 117958 476076 117964 476128
rect 118016 476116 118022 476128
rect 128446 476116 128452 476128
rect 118016 476088 128452 476116
rect 118016 476076 118022 476088
rect 128446 476076 128452 476088
rect 128504 476076 128510 476128
rect 102410 476008 102416 476060
rect 102468 476048 102474 476060
rect 103330 476048 103336 476060
rect 102468 476020 103336 476048
rect 102468 476008 102474 476020
rect 103330 476008 103336 476020
rect 103388 476048 103394 476060
rect 139394 476048 139400 476060
rect 103388 476020 139400 476048
rect 103388 476008 103394 476020
rect 139394 476008 139400 476020
rect 139452 476008 139458 476060
rect 102226 475940 102232 475992
rect 102284 475980 102290 475992
rect 117958 475980 117964 475992
rect 102284 475952 117964 475980
rect 102284 475940 102290 475952
rect 117958 475940 117964 475952
rect 118016 475940 118022 475992
rect 102318 475872 102324 475924
rect 102376 475912 102382 475924
rect 111886 475912 111892 475924
rect 102376 475884 111892 475912
rect 102376 475872 102382 475884
rect 111886 475872 111892 475884
rect 111944 475872 111950 475924
rect 51074 475396 51080 475448
rect 51132 475436 51138 475448
rect 52178 475436 52184 475448
rect 51132 475408 52184 475436
rect 51132 475396 51138 475408
rect 52178 475396 52184 475408
rect 52236 475436 52242 475448
rect 67634 475436 67640 475448
rect 52236 475408 67640 475436
rect 52236 475396 52242 475408
rect 67634 475396 67640 475408
rect 67692 475396 67698 475448
rect 35618 475328 35624 475380
rect 35676 475368 35682 475380
rect 65978 475368 65984 475380
rect 35676 475340 65984 475368
rect 35676 475328 35682 475340
rect 65978 475328 65984 475340
rect 66036 475368 66042 475380
rect 67726 475368 67732 475380
rect 66036 475340 67732 475368
rect 66036 475328 66042 475340
rect 67726 475328 67732 475340
rect 67784 475328 67790 475380
rect 111886 475328 111892 475380
rect 111944 475368 111950 475380
rect 121454 475368 121460 475380
rect 111944 475340 121460 475368
rect 111944 475328 111950 475340
rect 121454 475328 121460 475340
rect 121512 475328 121518 475380
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 25498 474756 25504 474768
rect 3476 474728 25504 474756
rect 3476 474716 3482 474728
rect 25498 474716 25504 474728
rect 25556 474716 25562 474768
rect 60366 474648 60372 474700
rect 60424 474688 60430 474700
rect 61930 474688 61936 474700
rect 60424 474660 61936 474688
rect 60424 474648 60430 474660
rect 61930 474648 61936 474660
rect 61988 474688 61994 474700
rect 67634 474688 67640 474700
rect 61988 474660 67640 474688
rect 61988 474648 61994 474660
rect 67634 474648 67640 474660
rect 67692 474648 67698 474700
rect 102226 474648 102232 474700
rect 102284 474688 102290 474700
rect 140866 474688 140872 474700
rect 102284 474660 140872 474688
rect 102284 474648 102290 474660
rect 140866 474648 140872 474660
rect 140924 474688 140930 474700
rect 141234 474688 141240 474700
rect 140924 474660 141240 474688
rect 140924 474648 140930 474660
rect 141234 474648 141240 474660
rect 141292 474648 141298 474700
rect 44082 473968 44088 474020
rect 44140 474008 44146 474020
rect 51074 474008 51080 474020
rect 44140 473980 51080 474008
rect 44140 473968 44146 473980
rect 51074 473968 51080 473980
rect 51132 473968 51138 474020
rect 113082 473968 113088 474020
rect 113140 474008 113146 474020
rect 117314 474008 117320 474020
rect 113140 473980 117320 474008
rect 113140 473968 113146 473980
rect 117314 473968 117320 473980
rect 117372 473968 117378 474020
rect 141234 473968 141240 474020
rect 141292 474008 141298 474020
rect 144914 474008 144920 474020
rect 141292 473980 144920 474008
rect 141292 473968 141298 473980
rect 144914 473968 144920 473980
rect 144972 473968 144978 474020
rect 65610 473396 65616 473408
rect 64846 473368 65616 473396
rect 49510 473288 49516 473340
rect 49568 473328 49574 473340
rect 64846 473328 64874 473368
rect 65610 473356 65616 473368
rect 65668 473396 65674 473408
rect 67634 473396 67640 473408
rect 65668 473368 67640 473396
rect 65668 473356 65674 473368
rect 67634 473356 67640 473368
rect 67692 473356 67698 473408
rect 49568 473300 64874 473328
rect 49568 473288 49574 473300
rect 100294 473288 100300 473340
rect 100352 473328 100358 473340
rect 100754 473328 100760 473340
rect 100352 473300 100760 473328
rect 100352 473288 100358 473300
rect 100754 473288 100760 473300
rect 100812 473288 100818 473340
rect 102318 472676 102324 472728
rect 102376 472716 102382 472728
rect 103422 472716 103428 472728
rect 102376 472688 103428 472716
rect 102376 472676 102382 472688
rect 103422 472676 103428 472688
rect 103480 472716 103486 472728
rect 109034 472716 109040 472728
rect 103480 472688 109040 472716
rect 103480 472676 103486 472688
rect 109034 472676 109040 472688
rect 109092 472676 109098 472728
rect 55030 472608 55036 472660
rect 55088 472648 55094 472660
rect 67634 472648 67640 472660
rect 55088 472620 67640 472648
rect 55088 472608 55094 472620
rect 67634 472608 67640 472620
rect 67692 472608 67698 472660
rect 102226 472608 102232 472660
rect 102284 472648 102290 472660
rect 143534 472648 143540 472660
rect 102284 472620 143540 472648
rect 102284 472608 102290 472620
rect 143534 472608 143540 472620
rect 143592 472608 143598 472660
rect 132586 472036 132592 472048
rect 106200 472008 132592 472036
rect 61930 471928 61936 471980
rect 61988 471968 61994 471980
rect 63218 471968 63224 471980
rect 61988 471940 63224 471968
rect 61988 471928 61994 471940
rect 63218 471928 63224 471940
rect 63276 471968 63282 471980
rect 67634 471968 67640 471980
rect 63276 471940 67640 471968
rect 63276 471928 63282 471940
rect 67634 471928 67640 471940
rect 67692 471928 67698 471980
rect 102226 471928 102232 471980
rect 102284 471968 102290 471980
rect 106200 471968 106228 472008
rect 132586 471996 132592 472008
rect 132644 471996 132650 472048
rect 102284 471940 106228 471968
rect 102284 471928 102290 471940
rect 102778 471316 102784 471368
rect 102836 471356 102842 471368
rect 135438 471356 135444 471368
rect 102836 471328 135444 471356
rect 102836 471316 102842 471328
rect 135438 471316 135444 471328
rect 135496 471356 135502 471368
rect 143626 471356 143632 471368
rect 135496 471328 143632 471356
rect 135496 471316 135502 471328
rect 143626 471316 143632 471328
rect 143684 471316 143690 471368
rect 109034 471248 109040 471300
rect 109092 471288 109098 471300
rect 146294 471288 146300 471300
rect 109092 471260 146300 471288
rect 109092 471248 109098 471260
rect 146294 471248 146300 471260
rect 146352 471248 146358 471300
rect 146294 470568 146300 470620
rect 146352 470608 146358 470620
rect 579982 470608 579988 470620
rect 146352 470580 579988 470608
rect 146352 470568 146358 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 66162 469888 66168 469940
rect 66220 469928 66226 469940
rect 67634 469928 67640 469940
rect 66220 469900 67640 469928
rect 66220 469888 66226 469900
rect 67634 469888 67640 469900
rect 67692 469888 67698 469940
rect 103514 469888 103520 469940
rect 103572 469928 103578 469940
rect 131390 469928 131396 469940
rect 103572 469900 131396 469928
rect 103572 469888 103578 469900
rect 131390 469888 131396 469900
rect 131448 469928 131454 469940
rect 139486 469928 139492 469940
rect 131448 469900 139492 469928
rect 131448 469888 131454 469900
rect 139486 469888 139492 469900
rect 139544 469888 139550 469940
rect 46658 469820 46664 469872
rect 46716 469860 46722 469872
rect 66180 469860 66208 469888
rect 46716 469832 66208 469860
rect 46716 469820 46722 469832
rect 102226 469820 102232 469872
rect 102284 469860 102290 469872
rect 134058 469860 134064 469872
rect 102284 469832 134064 469860
rect 102284 469820 102290 469832
rect 134058 469820 134064 469832
rect 134116 469820 134122 469872
rect 34238 469140 34244 469192
rect 34296 469180 34302 469192
rect 66990 469180 66996 469192
rect 34296 469152 66996 469180
rect 34296 469140 34302 469152
rect 66990 469140 66996 469152
rect 67048 469180 67054 469192
rect 67542 469180 67548 469192
rect 67048 469152 67548 469180
rect 67048 469140 67054 469152
rect 67542 469140 67548 469152
rect 67600 469140 67606 469192
rect 64598 467848 64604 467900
rect 64656 467888 64662 467900
rect 65978 467888 65984 467900
rect 64656 467860 65984 467888
rect 64656 467848 64662 467860
rect 65978 467848 65984 467860
rect 66036 467888 66042 467900
rect 67634 467888 67640 467900
rect 66036 467860 67640 467888
rect 66036 467848 66042 467860
rect 67634 467848 67640 467860
rect 67692 467848 67698 467900
rect 125502 467100 125508 467152
rect 125560 467140 125566 467152
rect 133874 467140 133880 467152
rect 125560 467112 133880 467140
rect 125560 467100 125566 467112
rect 133874 467100 133880 467112
rect 133932 467100 133938 467152
rect 108390 466556 108396 466608
rect 108448 466596 108454 466608
rect 113266 466596 113272 466608
rect 108448 466568 113272 466596
rect 108448 466556 108454 466568
rect 113266 466556 113272 466568
rect 113324 466556 113330 466608
rect 105630 466488 105636 466540
rect 105688 466528 105694 466540
rect 107838 466528 107844 466540
rect 105688 466500 107844 466528
rect 105688 466488 105694 466500
rect 107838 466488 107844 466500
rect 107896 466488 107902 466540
rect 64690 466420 64696 466472
rect 64748 466460 64754 466472
rect 67634 466460 67640 466472
rect 64748 466432 67640 466460
rect 64748 466420 64754 466432
rect 67634 466420 67640 466432
rect 67692 466420 67698 466472
rect 102226 466420 102232 466472
rect 102284 466460 102290 466472
rect 125502 466460 125508 466472
rect 102284 466432 125508 466460
rect 102284 466420 102290 466432
rect 125502 466420 125508 466432
rect 125560 466420 125566 466472
rect 102318 465808 102324 465860
rect 102376 465848 102382 465860
rect 107746 465848 107752 465860
rect 102376 465820 107752 465848
rect 102376 465808 102382 465820
rect 107746 465808 107752 465820
rect 107804 465848 107810 465860
rect 116578 465848 116584 465860
rect 107804 465820 116584 465848
rect 107804 465808 107810 465820
rect 116578 465808 116584 465820
rect 116636 465808 116642 465860
rect 102226 465740 102232 465792
rect 102284 465780 102290 465792
rect 116026 465780 116032 465792
rect 102284 465752 116032 465780
rect 102284 465740 102290 465752
rect 116026 465740 116032 465752
rect 116084 465780 116090 465792
rect 116670 465780 116676 465792
rect 116084 465752 116676 465780
rect 116084 465740 116090 465752
rect 116670 465740 116676 465752
rect 116728 465740 116734 465792
rect 103514 465672 103520 465724
rect 103572 465712 103578 465724
rect 136818 465712 136824 465724
rect 103572 465684 136824 465712
rect 103572 465672 103578 465684
rect 136818 465672 136824 465684
rect 136876 465712 136882 465724
rect 138106 465712 138112 465724
rect 136876 465684 138112 465712
rect 136876 465672 136882 465684
rect 138106 465672 138112 465684
rect 138164 465672 138170 465724
rect 67634 465100 67640 465112
rect 50356 465072 67640 465100
rect 50356 465044 50384 465072
rect 67634 465060 67640 465072
rect 67692 465060 67698 465112
rect 48038 464992 48044 465044
rect 48096 465032 48102 465044
rect 50338 465032 50344 465044
rect 48096 465004 50344 465032
rect 48096 464992 48102 465004
rect 50338 464992 50344 465004
rect 50396 464992 50402 465044
rect 59170 464992 59176 465044
rect 59228 465032 59234 465044
rect 63126 465032 63132 465044
rect 59228 465004 63132 465032
rect 59228 464992 59234 465004
rect 63126 464992 63132 465004
rect 63184 465032 63190 465044
rect 67726 465032 67732 465044
rect 63184 465004 67732 465032
rect 63184 464992 63190 465004
rect 67726 464992 67732 465004
rect 67784 464992 67790 465044
rect 104710 464108 104716 464160
rect 104768 464148 104774 464160
rect 107654 464148 107660 464160
rect 104768 464120 107660 464148
rect 104768 464108 104774 464120
rect 107654 464108 107660 464120
rect 107712 464108 107718 464160
rect 67634 463740 67640 463752
rect 57256 463712 67640 463740
rect 57256 463684 57284 463712
rect 67634 463700 67640 463712
rect 67692 463700 67698 463752
rect 56502 463632 56508 463684
rect 56560 463672 56566 463684
rect 57238 463672 57244 463684
rect 56560 463644 57244 463672
rect 56560 463632 56566 463644
rect 57238 463632 57244 463644
rect 57296 463632 57302 463684
rect 125594 463632 125600 463684
rect 125652 463672 125658 463684
rect 125962 463672 125968 463684
rect 125652 463644 125968 463672
rect 125652 463632 125658 463644
rect 125962 463632 125968 463644
rect 126020 463632 126026 463684
rect 52454 462952 52460 463004
rect 52512 462992 52518 463004
rect 53558 462992 53564 463004
rect 52512 462964 53564 462992
rect 52512 462952 52518 462964
rect 53558 462952 53564 462964
rect 53616 462992 53622 463004
rect 67634 462992 67640 463004
rect 53616 462964 67640 462992
rect 53616 462952 53622 462964
rect 67634 462952 67640 462964
rect 67692 462952 67698 463004
rect 102226 462952 102232 463004
rect 102284 462992 102290 463004
rect 125594 462992 125600 463004
rect 102284 462964 125600 462992
rect 102284 462952 102290 462964
rect 125594 462952 125600 462964
rect 125652 462952 125658 463004
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4798 462584 4804 462596
rect 2832 462556 4804 462584
rect 2832 462544 2838 462556
rect 4798 462544 4804 462556
rect 4856 462544 4862 462596
rect 61746 462340 61752 462392
rect 61804 462380 61810 462392
rect 64598 462380 64604 462392
rect 61804 462352 64604 462380
rect 61804 462340 61810 462352
rect 64598 462340 64604 462352
rect 64656 462380 64662 462392
rect 67634 462380 67640 462392
rect 64656 462352 67640 462380
rect 64656 462340 64662 462352
rect 67634 462340 67640 462352
rect 67692 462340 67698 462392
rect 107562 462340 107568 462392
rect 107620 462380 107626 462392
rect 140958 462380 140964 462392
rect 107620 462352 140964 462380
rect 107620 462340 107626 462352
rect 140958 462340 140964 462352
rect 141016 462340 141022 462392
rect 48222 462272 48228 462324
rect 48280 462312 48286 462324
rect 52454 462312 52460 462324
rect 48280 462284 52460 462312
rect 48280 462272 48286 462284
rect 52454 462272 52460 462284
rect 52512 462272 52518 462324
rect 58986 462272 58992 462324
rect 59044 462312 59050 462324
rect 63126 462312 63132 462324
rect 59044 462284 63132 462312
rect 59044 462272 59050 462284
rect 63126 462272 63132 462284
rect 63184 462272 63190 462324
rect 102318 462272 102324 462324
rect 102376 462312 102382 462324
rect 129918 462312 129924 462324
rect 102376 462284 129924 462312
rect 102376 462272 102382 462284
rect 129918 462272 129924 462284
rect 129976 462312 129982 462324
rect 130378 462312 130384 462324
rect 129976 462284 130384 462312
rect 129976 462272 129982 462284
rect 130378 462272 130384 462284
rect 130436 462272 130442 462324
rect 102226 462204 102232 462256
rect 102284 462244 102290 462256
rect 107562 462244 107568 462256
rect 102284 462216 107568 462244
rect 102284 462204 102290 462216
rect 107562 462204 107568 462216
rect 107620 462204 107626 462256
rect 116670 462204 116676 462256
rect 116728 462244 116734 462256
rect 120718 462244 120724 462256
rect 116728 462216 120724 462244
rect 116728 462204 116734 462216
rect 120718 462204 120724 462216
rect 120776 462204 120782 462256
rect 63126 460912 63132 460964
rect 63184 460952 63190 460964
rect 67634 460952 67640 460964
rect 63184 460924 67640 460952
rect 63184 460912 63190 460924
rect 67634 460912 67640 460924
rect 67692 460912 67698 460964
rect 102318 460844 102324 460896
rect 102376 460884 102382 460896
rect 106642 460884 106648 460896
rect 102376 460856 106648 460884
rect 102376 460844 102382 460856
rect 106642 460844 106648 460856
rect 106700 460844 106706 460896
rect 102134 460300 102140 460352
rect 102192 460340 102198 460352
rect 105538 460340 105544 460352
rect 102192 460312 105544 460340
rect 102192 460300 102198 460312
rect 105538 460300 105544 460312
rect 105596 460300 105602 460352
rect 54202 460232 54208 460284
rect 54260 460272 54266 460284
rect 55122 460272 55128 460284
rect 54260 460244 55128 460272
rect 54260 460232 54266 460244
rect 55122 460232 55128 460244
rect 55180 460272 55186 460284
rect 67634 460272 67640 460284
rect 55180 460244 67640 460272
rect 55180 460232 55186 460244
rect 67634 460232 67640 460244
rect 67692 460232 67698 460284
rect 41230 460164 41236 460216
rect 41288 460204 41294 460216
rect 67726 460204 67732 460216
rect 41288 460176 67732 460204
rect 41288 460164 41294 460176
rect 67726 460164 67732 460176
rect 67784 460164 67790 460216
rect 40954 459552 40960 459604
rect 41012 459592 41018 459604
rect 41230 459592 41236 459604
rect 41012 459564 41236 459592
rect 41012 459552 41018 459564
rect 41230 459552 41236 459564
rect 41288 459552 41294 459604
rect 107010 459552 107016 459604
rect 107068 459592 107074 459604
rect 114738 459592 114744 459604
rect 107068 459564 114744 459592
rect 107068 459552 107074 459564
rect 114738 459552 114744 459564
rect 114796 459552 114802 459604
rect 124950 459552 124956 459604
rect 125008 459592 125014 459604
rect 133966 459592 133972 459604
rect 125008 459564 133972 459592
rect 125008 459552 125014 459564
rect 133966 459552 133972 459564
rect 134024 459552 134030 459604
rect 102134 459484 102140 459536
rect 102192 459524 102198 459536
rect 124968 459524 124996 459552
rect 102192 459496 124996 459524
rect 102192 459484 102198 459496
rect 108206 458804 108212 458856
rect 108264 458844 108270 458856
rect 134242 458844 134248 458856
rect 108264 458816 134248 458844
rect 108264 458804 108270 458816
rect 134242 458804 134248 458816
rect 134300 458844 134306 458856
rect 149238 458844 149244 458856
rect 134300 458816 149244 458844
rect 134300 458804 134306 458816
rect 149238 458804 149244 458816
rect 149296 458804 149302 458856
rect 48038 458192 48044 458244
rect 48096 458232 48102 458244
rect 54202 458232 54208 458244
rect 48096 458204 54208 458232
rect 48096 458192 48102 458204
rect 54202 458192 54208 458204
rect 54260 458192 54266 458244
rect 64782 458192 64788 458244
rect 64840 458232 64846 458244
rect 67634 458232 67640 458244
rect 64840 458204 67640 458232
rect 64840 458192 64846 458204
rect 67634 458192 67640 458204
rect 67692 458192 67698 458244
rect 102134 458192 102140 458244
rect 102192 458232 102198 458244
rect 102192 458204 115888 458232
rect 102192 458192 102198 458204
rect 115860 458176 115888 458204
rect 102318 458124 102324 458176
rect 102376 458164 102382 458176
rect 108206 458164 108212 458176
rect 102376 458136 108212 458164
rect 102376 458124 102382 458136
rect 108206 458124 108212 458136
rect 108264 458124 108270 458176
rect 115842 458164 115848 458176
rect 115755 458136 115848 458164
rect 115842 458124 115848 458136
rect 115900 458164 115906 458176
rect 120074 458164 120080 458176
rect 115900 458136 120080 458164
rect 115900 458124 115906 458136
rect 120074 458124 120080 458136
rect 120132 458124 120138 458176
rect 103514 457444 103520 457496
rect 103572 457484 103578 457496
rect 139578 457484 139584 457496
rect 103572 457456 139584 457484
rect 103572 457444 103578 457456
rect 139578 457444 139584 457456
rect 139636 457484 139642 457496
rect 142246 457484 142252 457496
rect 139636 457456 142252 457484
rect 139636 457444 139642 457456
rect 142246 457444 142252 457456
rect 142304 457444 142310 457496
rect 52454 456832 52460 456884
rect 52512 456872 52518 456884
rect 53190 456872 53196 456884
rect 52512 456844 53196 456872
rect 52512 456832 52518 456844
rect 53190 456832 53196 456844
rect 53248 456872 53254 456884
rect 67634 456872 67640 456884
rect 53248 456844 67640 456872
rect 53248 456832 53254 456844
rect 67634 456832 67640 456844
rect 67692 456832 67698 456884
rect 67726 456804 67732 456816
rect 45526 456776 67732 456804
rect 42702 456696 42708 456748
rect 42760 456736 42766 456748
rect 44818 456736 44824 456748
rect 42760 456708 44824 456736
rect 42760 456696 42766 456708
rect 44818 456696 44824 456708
rect 44876 456736 44882 456748
rect 45526 456736 45554 456776
rect 67726 456764 67732 456776
rect 67784 456764 67790 456816
rect 377398 456764 377404 456816
rect 377456 456804 377462 456816
rect 580166 456804 580172 456816
rect 377456 456776 580172 456804
rect 377456 456764 377462 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 44876 456708 45554 456736
rect 44876 456696 44882 456708
rect 48130 456696 48136 456748
rect 48188 456736 48194 456748
rect 52454 456736 52460 456748
rect 48188 456708 52460 456736
rect 48188 456696 48194 456708
rect 52454 456696 52460 456708
rect 52512 456696 52518 456748
rect 102134 456696 102140 456748
rect 102192 456736 102198 456748
rect 142154 456736 142160 456748
rect 102192 456708 142160 456736
rect 102192 456696 102198 456708
rect 142154 456696 142160 456708
rect 142212 456736 142218 456748
rect 143442 456736 143448 456748
rect 142212 456708 143448 456736
rect 142212 456696 142218 456708
rect 143442 456696 143448 456708
rect 143500 456696 143506 456748
rect 143442 456016 143448 456068
rect 143500 456056 143506 456068
rect 151906 456056 151912 456068
rect 143500 456028 151912 456056
rect 143500 456016 143506 456028
rect 151906 456016 151912 456028
rect 151964 456016 151970 456068
rect 30282 455404 30288 455456
rect 30340 455444 30346 455456
rect 67634 455444 67640 455456
rect 30340 455416 35894 455444
rect 30340 455404 30346 455416
rect 35866 455376 35894 455416
rect 64846 455416 67640 455444
rect 36538 455376 36544 455388
rect 35866 455348 36544 455376
rect 36538 455336 36544 455348
rect 36596 455376 36602 455388
rect 64846 455376 64874 455416
rect 67634 455404 67640 455416
rect 67692 455404 67698 455456
rect 36596 455348 64874 455376
rect 36596 455336 36602 455348
rect 102870 455336 102876 455388
rect 102928 455376 102934 455388
rect 105630 455376 105636 455388
rect 102928 455348 105636 455376
rect 102928 455336 102934 455348
rect 105630 455336 105636 455348
rect 105688 455336 105694 455388
rect 56318 455268 56324 455320
rect 56376 455308 56382 455320
rect 56502 455308 56508 455320
rect 56376 455280 56508 455308
rect 56376 455268 56382 455280
rect 56502 455268 56508 455280
rect 56560 455268 56566 455320
rect 106182 454792 106188 454844
rect 106240 454832 106246 454844
rect 114830 454832 114836 454844
rect 106240 454804 114836 454832
rect 106240 454792 106246 454804
rect 114830 454792 114836 454804
rect 114888 454792 114894 454844
rect 108206 454724 108212 454776
rect 108264 454764 108270 454776
rect 138198 454764 138204 454776
rect 108264 454736 138204 454764
rect 108264 454724 108270 454736
rect 138198 454724 138204 454736
rect 138256 454764 138262 454776
rect 150526 454764 150532 454776
rect 138256 454736 150532 454764
rect 138256 454724 138262 454736
rect 150526 454724 150532 454736
rect 150584 454724 150590 454776
rect 56502 454656 56508 454708
rect 56560 454696 56566 454708
rect 67634 454696 67640 454708
rect 56560 454668 67640 454696
rect 56560 454656 56566 454668
rect 67634 454656 67640 454668
rect 67692 454656 67698 454708
rect 102134 454656 102140 454708
rect 102192 454696 102198 454708
rect 135346 454696 135352 454708
rect 102192 454668 135352 454696
rect 102192 454656 102198 454668
rect 135346 454656 135352 454668
rect 135404 454656 135410 454708
rect 102134 453976 102140 454028
rect 102192 454016 102198 454028
rect 118970 454016 118976 454028
rect 102192 453988 118976 454016
rect 102192 453976 102198 453988
rect 118970 453976 118976 453988
rect 119028 453976 119034 454028
rect 102318 453908 102324 453960
rect 102376 453948 102382 453960
rect 108206 453948 108212 453960
rect 102376 453920 108212 453948
rect 102376 453908 102382 453920
rect 108206 453908 108212 453920
rect 108264 453908 108270 453960
rect 55122 453364 55128 453416
rect 55180 453404 55186 453416
rect 57698 453404 57704 453416
rect 55180 453376 57704 453404
rect 55180 453364 55186 453376
rect 57698 453364 57704 453376
rect 57756 453404 57762 453416
rect 67634 453404 67640 453416
rect 57756 453376 67640 453404
rect 57756 453364 57762 453376
rect 67634 453364 67640 453376
rect 67692 453364 67698 453416
rect 54938 453296 54944 453348
rect 54996 453336 55002 453348
rect 67726 453336 67732 453348
rect 54996 453308 67732 453336
rect 54996 453296 55002 453308
rect 67726 453296 67732 453308
rect 67784 453296 67790 453348
rect 52086 451936 52092 451988
rect 52144 451976 52150 451988
rect 54938 451976 54944 451988
rect 52144 451948 54944 451976
rect 52144 451936 52150 451948
rect 54938 451936 54944 451948
rect 54996 451936 55002 451988
rect 102134 451936 102140 451988
rect 102192 451976 102198 451988
rect 115934 451976 115940 451988
rect 102192 451948 115940 451976
rect 102192 451936 102198 451948
rect 115934 451936 115940 451948
rect 115992 451936 115998 451988
rect 102502 451868 102508 451920
rect 102560 451908 102566 451920
rect 134150 451908 134156 451920
rect 102560 451880 134156 451908
rect 102560 451868 102566 451880
rect 134150 451868 134156 451880
rect 134208 451908 134214 451920
rect 147766 451908 147772 451920
rect 134208 451880 147772 451908
rect 134208 451868 134214 451880
rect 147766 451868 147772 451880
rect 147824 451868 147830 451920
rect 101950 451188 101956 451240
rect 102008 451228 102014 451240
rect 105722 451228 105728 451240
rect 102008 451200 105728 451228
rect 102008 451188 102014 451200
rect 105722 451188 105728 451200
rect 105780 451188 105786 451240
rect 100110 450508 100116 450560
rect 100168 450548 100174 450560
rect 109126 450548 109132 450560
rect 100168 450520 109132 450548
rect 100168 450508 100174 450520
rect 109126 450508 109132 450520
rect 109184 450508 109190 450560
rect 61838 449896 61844 449948
rect 61896 449936 61902 449948
rect 64414 449936 64420 449948
rect 61896 449908 64420 449936
rect 61896 449896 61902 449908
rect 64414 449896 64420 449908
rect 64472 449936 64478 449948
rect 67634 449936 67640 449948
rect 64472 449908 67640 449936
rect 64472 449896 64478 449908
rect 67634 449896 67640 449908
rect 67692 449896 67698 449948
rect 106918 449896 106924 449948
rect 106976 449936 106982 449948
rect 122834 449936 122840 449948
rect 106976 449908 122840 449936
rect 106976 449896 106982 449908
rect 122834 449896 122840 449908
rect 122892 449896 122898 449948
rect 102318 449828 102324 449880
rect 102376 449868 102382 449880
rect 106936 449868 106964 449896
rect 102376 449840 106964 449868
rect 102376 449828 102382 449840
rect 102134 449760 102140 449812
rect 102192 449800 102198 449812
rect 105354 449800 105360 449812
rect 102192 449772 105360 449800
rect 102192 449760 102198 449772
rect 105354 449760 105360 449772
rect 105412 449760 105418 449812
rect 63310 448536 63316 448588
rect 63368 448576 63374 448588
rect 64690 448576 64696 448588
rect 63368 448548 64696 448576
rect 63368 448536 63374 448548
rect 64690 448536 64696 448548
rect 64748 448576 64754 448588
rect 67634 448576 67640 448588
rect 64748 448548 67640 448576
rect 64748 448536 64754 448548
rect 67634 448536 67640 448548
rect 67692 448536 67698 448588
rect 102134 447924 102140 447976
rect 102192 447964 102198 447976
rect 107010 447964 107016 447976
rect 102192 447936 107016 447964
rect 102192 447924 102198 447936
rect 107010 447924 107016 447936
rect 107068 447924 107074 447976
rect 104710 447856 104716 447908
rect 104768 447896 104774 447908
rect 114922 447896 114928 447908
rect 104768 447868 114928 447896
rect 104768 447856 104774 447868
rect 114922 447856 114928 447868
rect 114980 447856 114986 447908
rect 102318 447788 102324 447840
rect 102376 447828 102382 447840
rect 127066 447828 127072 447840
rect 102376 447800 127072 447828
rect 102376 447788 102382 447800
rect 127066 447788 127072 447800
rect 127124 447788 127130 447840
rect 61378 447148 61384 447160
rect 60752 447120 61384 447148
rect 60752 447080 60780 447120
rect 61378 447108 61384 447120
rect 61436 447148 61442 447160
rect 67634 447148 67640 447160
rect 61436 447120 67640 447148
rect 61436 447108 61442 447120
rect 67634 447108 67640 447120
rect 67692 447108 67698 447160
rect 45526 447052 60780 447080
rect 34330 446972 34336 447024
rect 34388 447012 34394 447024
rect 45526 447012 45554 447052
rect 34388 446984 45554 447012
rect 34388 446972 34394 446984
rect 60734 445748 60740 445800
rect 60792 445788 60798 445800
rect 61746 445788 61752 445800
rect 60792 445760 61752 445788
rect 60792 445748 60798 445760
rect 61746 445748 61752 445760
rect 61804 445788 61810 445800
rect 67634 445788 67640 445800
rect 61804 445760 67640 445788
rect 61804 445748 61810 445760
rect 67634 445748 67640 445760
rect 67692 445748 67698 445800
rect 101030 445748 101036 445800
rect 101088 445788 101094 445800
rect 102042 445788 102048 445800
rect 101088 445760 102048 445788
rect 101088 445748 101094 445760
rect 102042 445748 102048 445760
rect 102100 445788 102106 445800
rect 146386 445788 146392 445800
rect 102100 445760 146392 445788
rect 102100 445748 102106 445760
rect 146386 445748 146392 445760
rect 146444 445748 146450 445800
rect 102134 445680 102140 445732
rect 102192 445720 102198 445732
rect 103698 445720 103704 445732
rect 102192 445692 103704 445720
rect 102192 445680 102198 445692
rect 103698 445680 103704 445692
rect 103756 445720 103762 445732
rect 104158 445720 104164 445732
rect 103756 445692 104164 445720
rect 103756 445680 103762 445692
rect 104158 445680 104164 445692
rect 104216 445680 104222 445732
rect 102318 445272 102324 445324
rect 102376 445312 102382 445324
rect 104894 445312 104900 445324
rect 102376 445284 104900 445312
rect 102376 445272 102382 445284
rect 104894 445272 104900 445284
rect 104952 445312 104958 445324
rect 105630 445312 105636 445324
rect 104952 445284 105636 445312
rect 104952 445272 104958 445284
rect 105630 445272 105636 445284
rect 105688 445272 105694 445324
rect 104802 445068 104808 445120
rect 104860 445108 104866 445120
rect 128538 445108 128544 445120
rect 104860 445080 128544 445108
rect 104860 445068 104866 445080
rect 128538 445068 128544 445080
rect 128596 445068 128602 445120
rect 36998 445000 37004 445052
rect 37056 445040 37062 445052
rect 67634 445040 67640 445052
rect 37056 445012 67640 445040
rect 37056 445000 37062 445012
rect 67634 445000 67640 445012
rect 67692 445000 67698 445052
rect 102134 445000 102140 445052
rect 102192 445040 102198 445052
rect 132678 445040 132684 445052
rect 102192 445012 132684 445040
rect 102192 445000 102198 445012
rect 132678 445000 132684 445012
rect 132736 445040 132742 445052
rect 142154 445040 142160 445052
rect 132736 445012 142160 445040
rect 132736 445000 132742 445012
rect 142154 445000 142160 445012
rect 142212 445000 142218 445052
rect 102318 443980 102324 444032
rect 102376 444020 102382 444032
rect 104802 444020 104808 444032
rect 102376 443992 104808 444020
rect 102376 443980 102382 443992
rect 104802 443980 104808 443992
rect 104860 443980 104866 444032
rect 34330 443640 34336 443692
rect 34388 443680 34394 443692
rect 67634 443680 67640 443692
rect 34388 443652 67640 443680
rect 34388 443640 34394 443652
rect 67634 443640 67640 443652
rect 67692 443640 67698 443692
rect 113082 443640 113088 443692
rect 113140 443680 113146 443692
rect 123110 443680 123116 443692
rect 113140 443652 123116 443680
rect 113140 443640 113146 443652
rect 123110 443640 123116 443652
rect 123168 443640 123174 443692
rect 33042 442892 33048 442944
rect 33100 442932 33106 442944
rect 34146 442932 34152 442944
rect 33100 442904 34152 442932
rect 33100 442892 33106 442904
rect 34146 442892 34152 442904
rect 34204 442932 34210 442944
rect 67634 442932 67640 442944
rect 34204 442904 67640 442932
rect 34204 442892 34210 442904
rect 67634 442892 67640 442904
rect 67692 442892 67698 442944
rect 49602 442824 49608 442876
rect 49660 442864 49666 442876
rect 66254 442864 66260 442876
rect 49660 442836 66260 442864
rect 49660 442824 49666 442836
rect 66254 442824 66260 442836
rect 66312 442824 66318 442876
rect 60274 442756 60280 442808
rect 60332 442796 60338 442808
rect 61838 442796 61844 442808
rect 60332 442768 61844 442796
rect 60332 442756 60338 442768
rect 61838 442756 61844 442768
rect 61896 442796 61902 442808
rect 67726 442796 67732 442808
rect 61896 442768 67732 442796
rect 61896 442756 61902 442768
rect 67726 442756 67732 442768
rect 67784 442756 67790 442808
rect 64414 442280 64420 442332
rect 64472 442320 64478 442332
rect 64782 442320 64788 442332
rect 64472 442292 64788 442320
rect 64472 442280 64478 442292
rect 64782 442280 64788 442292
rect 64840 442280 64846 442332
rect 102134 441600 102140 441652
rect 102192 441640 102198 441652
rect 102192 441612 108988 441640
rect 102192 441600 102198 441612
rect 62022 441532 62028 441584
rect 62080 441572 62086 441584
rect 63310 441572 63316 441584
rect 62080 441544 63316 441572
rect 62080 441532 62086 441544
rect 63310 441532 63316 441544
rect 63368 441532 63374 441584
rect 63402 441532 63408 441584
rect 63460 441572 63466 441584
rect 66162 441572 66168 441584
rect 63460 441544 66168 441572
rect 63460 441532 63466 441544
rect 66162 441532 66168 441544
rect 66220 441532 66226 441584
rect 108960 441572 108988 441612
rect 129826 441572 129832 441584
rect 108960 441544 129832 441572
rect 129826 441532 129832 441544
rect 129884 441532 129890 441584
rect 66162 441124 66168 441176
rect 66220 441164 66226 441176
rect 67634 441164 67640 441176
rect 66220 441136 67640 441164
rect 66220 441124 66226 441136
rect 67634 441124 67640 441136
rect 67692 441124 67698 441176
rect 63310 440988 63316 441040
rect 63368 441028 63374 441040
rect 67634 441028 67640 441040
rect 63368 441000 67640 441028
rect 63368 440988 63374 441000
rect 67634 440988 67640 441000
rect 67692 440988 67698 441040
rect 56226 440920 56232 440972
rect 56284 440960 56290 440972
rect 56284 440932 70394 440960
rect 56284 440920 56290 440932
rect 43806 440852 43812 440904
rect 43864 440892 43870 440904
rect 43864 440864 60734 440892
rect 43864 440852 43870 440864
rect 60706 440688 60734 440864
rect 70366 440756 70394 440932
rect 116118 440892 116124 440904
rect 103486 440864 116124 440892
rect 103486 440756 103514 440864
rect 116118 440852 116124 440864
rect 116176 440852 116182 440904
rect 129826 440852 129832 440904
rect 129884 440892 129890 440904
rect 139578 440892 139584 440904
rect 129884 440864 139584 440892
rect 129884 440852 129890 440864
rect 139578 440852 139584 440864
rect 139636 440852 139642 440904
rect 70366 440728 79364 440756
rect 79336 440700 79364 440728
rect 94148 440728 103514 440756
rect 94148 440700 94176 440728
rect 71774 440688 71780 440700
rect 60706 440660 71780 440688
rect 71774 440648 71780 440660
rect 71832 440688 71838 440700
rect 72326 440688 72332 440700
rect 71832 440660 72332 440688
rect 71832 440648 71838 440660
rect 72326 440648 72332 440660
rect 72384 440648 72390 440700
rect 79318 440648 79324 440700
rect 79376 440648 79382 440700
rect 94130 440648 94136 440700
rect 94188 440648 94194 440700
rect 97442 440648 97448 440700
rect 97500 440688 97506 440700
rect 99926 440688 99932 440700
rect 97500 440660 99932 440688
rect 97500 440648 97506 440660
rect 99926 440648 99932 440660
rect 99984 440648 99990 440700
rect 100754 440308 100760 440360
rect 100812 440348 100818 440360
rect 131114 440348 131120 440360
rect 100812 440320 131120 440348
rect 100812 440308 100818 440320
rect 131114 440308 131120 440320
rect 131172 440308 131178 440360
rect 99466 440240 99472 440292
rect 99524 440280 99530 440292
rect 100846 440280 100852 440292
rect 99524 440252 100852 440280
rect 99524 440240 99530 440252
rect 100846 440240 100852 440252
rect 100904 440280 100910 440292
rect 136818 440280 136824 440292
rect 100904 440252 136824 440280
rect 100904 440240 100910 440252
rect 136818 440240 136824 440252
rect 136876 440240 136882 440292
rect 95326 440172 95332 440224
rect 95384 440212 95390 440224
rect 100110 440212 100116 440224
rect 95384 440184 100116 440212
rect 95384 440172 95390 440184
rect 97276 439952 97304 440184
rect 100110 440172 100116 440184
rect 100168 440172 100174 440224
rect 97902 440104 97908 440156
rect 97960 440144 97966 440156
rect 103606 440144 103612 440156
rect 97960 440116 103612 440144
rect 97960 440104 97966 440116
rect 103606 440104 103612 440116
rect 103664 440104 103670 440156
rect 97258 439900 97264 439952
rect 97316 439900 97322 439952
rect 69198 439560 69204 439612
rect 69256 439600 69262 439612
rect 76558 439600 76564 439612
rect 69256 439572 76564 439600
rect 69256 439560 69262 439572
rect 76558 439560 76564 439572
rect 76616 439560 76622 439612
rect 95142 439560 95148 439612
rect 95200 439600 95206 439612
rect 110598 439600 110604 439612
rect 95200 439572 110604 439600
rect 95200 439560 95206 439572
rect 110598 439560 110604 439572
rect 110656 439560 110662 439612
rect 50706 439492 50712 439544
rect 50764 439532 50770 439544
rect 79318 439532 79324 439544
rect 50764 439504 79324 439532
rect 50764 439492 50770 439504
rect 79318 439492 79324 439504
rect 79376 439532 79382 439544
rect 81434 439532 81440 439544
rect 79376 439504 81440 439532
rect 79376 439492 79382 439504
rect 81434 439492 81440 439504
rect 81492 439492 81498 439544
rect 96522 439492 96528 439544
rect 96580 439532 96586 439544
rect 120442 439532 120448 439544
rect 96580 439504 120448 439532
rect 96580 439492 96586 439504
rect 120442 439492 120448 439504
rect 120500 439492 120506 439544
rect 69106 439016 69112 439068
rect 69164 439056 69170 439068
rect 73798 439056 73804 439068
rect 69164 439028 73804 439056
rect 69164 439016 69170 439028
rect 73798 439016 73804 439028
rect 73856 439016 73862 439068
rect 79778 439016 79784 439068
rect 79836 439056 79842 439068
rect 82814 439056 82820 439068
rect 79836 439028 82820 439056
rect 79836 439016 79842 439028
rect 82814 439016 82820 439028
rect 82872 439016 82878 439068
rect 46750 438948 46756 439000
rect 46808 438988 46814 439000
rect 80974 438988 80980 439000
rect 46808 438960 80980 438988
rect 46808 438948 46814 438960
rect 80974 438948 80980 438960
rect 81032 438948 81038 439000
rect 88702 438948 88708 439000
rect 88760 438988 88766 439000
rect 121638 438988 121644 439000
rect 88760 438960 121644 438988
rect 88760 438948 88766 438960
rect 121638 438948 121644 438960
rect 121696 438948 121702 439000
rect 25498 438880 25504 438932
rect 25556 438920 25562 438932
rect 25556 438892 96476 438920
rect 25556 438880 25562 438892
rect 96448 438864 96476 438892
rect 96614 438880 96620 438932
rect 96672 438920 96678 438932
rect 97718 438920 97724 438932
rect 96672 438892 97724 438920
rect 96672 438880 96678 438892
rect 97718 438880 97724 438892
rect 97776 438880 97782 438932
rect 75178 438812 75184 438864
rect 75236 438852 75242 438864
rect 82262 438852 82268 438864
rect 75236 438824 82268 438852
rect 75236 438812 75242 438824
rect 82262 438812 82268 438824
rect 82320 438812 82326 438864
rect 86126 438812 86132 438864
rect 86184 438852 86190 438864
rect 94498 438852 94504 438864
rect 86184 438824 94504 438852
rect 86184 438812 86190 438824
rect 94498 438812 94504 438824
rect 94556 438852 94562 438864
rect 95142 438852 95148 438864
rect 94556 438824 95148 438852
rect 94556 438812 94562 438824
rect 95142 438812 95148 438824
rect 95200 438812 95206 438864
rect 96430 438812 96436 438864
rect 96488 438852 96494 438864
rect 96488 438824 96660 438852
rect 96488 438812 96494 438824
rect 50890 438744 50896 438796
rect 50948 438784 50954 438796
rect 82906 438784 82912 438796
rect 50948 438756 82912 438784
rect 50948 438744 50954 438756
rect 82906 438744 82912 438756
rect 82964 438744 82970 438796
rect 84194 438744 84200 438796
rect 84252 438784 84258 438796
rect 85574 438784 85580 438796
rect 84252 438756 85580 438784
rect 84252 438744 84258 438756
rect 85574 438744 85580 438756
rect 85632 438744 85638 438796
rect 91278 438744 91284 438796
rect 91336 438784 91342 438796
rect 95234 438784 95240 438796
rect 91336 438756 95240 438784
rect 91336 438744 91342 438756
rect 95234 438744 95240 438756
rect 95292 438784 95298 438796
rect 96522 438784 96528 438796
rect 95292 438756 96528 438784
rect 95292 438744 95298 438756
rect 96522 438744 96528 438756
rect 96580 438744 96586 438796
rect 96632 438784 96660 438824
rect 99006 438812 99012 438864
rect 99064 438852 99070 438864
rect 121730 438852 121736 438864
rect 99064 438824 121736 438852
rect 99064 438812 99070 438824
rect 121730 438812 121736 438824
rect 121788 438852 121794 438864
rect 124214 438852 124220 438864
rect 121788 438824 124220 438852
rect 121788 438812 121794 438824
rect 124214 438812 124220 438824
rect 124272 438812 124278 438864
rect 123018 438784 123024 438796
rect 96632 438756 123024 438784
rect 123018 438744 123024 438756
rect 123076 438744 123082 438796
rect 51994 438676 52000 438728
rect 52052 438716 52058 438728
rect 83550 438716 83556 438728
rect 52052 438688 83556 438716
rect 52052 438676 52058 438688
rect 83550 438676 83556 438688
rect 83608 438676 83614 438728
rect 70394 438608 70400 438660
rect 70452 438648 70458 438660
rect 77110 438648 77116 438660
rect 70452 438620 77116 438648
rect 70452 438608 70458 438620
rect 77110 438608 77116 438620
rect 77168 438608 77174 438660
rect 88242 438608 88248 438660
rect 88300 438648 88306 438660
rect 105722 438648 105728 438660
rect 88300 438620 105728 438648
rect 88300 438608 88306 438620
rect 105722 438608 105728 438620
rect 105780 438608 105786 438660
rect 3418 438540 3424 438592
rect 3476 438580 3482 438592
rect 99374 438580 99380 438592
rect 3476 438552 99380 438580
rect 3476 438540 3482 438552
rect 99374 438540 99380 438552
rect 99432 438540 99438 438592
rect 93578 438472 93584 438524
rect 93636 438512 93642 438524
rect 93946 438512 93952 438524
rect 93636 438484 93952 438512
rect 93636 438472 93642 438484
rect 93946 438472 93952 438484
rect 94004 438472 94010 438524
rect 87414 438268 87420 438320
rect 87472 438308 87478 438320
rect 88242 438308 88248 438320
rect 87472 438280 88248 438308
rect 87472 438268 87478 438280
rect 88242 438268 88248 438280
rect 88300 438268 88306 438320
rect 56318 438200 56324 438252
rect 56376 438240 56382 438252
rect 73890 438240 73896 438252
rect 56376 438212 73896 438240
rect 56376 438200 56382 438212
rect 73890 438200 73896 438212
rect 73948 438200 73954 438252
rect 4798 438132 4804 438184
rect 4856 438172 4862 438184
rect 49510 438172 49516 438184
rect 4856 438144 49516 438172
rect 4856 438132 4862 438144
rect 49510 438132 49516 438144
rect 49568 438172 49574 438184
rect 51994 438172 52000 438184
rect 49568 438144 52000 438172
rect 49568 438132 49574 438144
rect 51994 438132 52000 438144
rect 52052 438132 52058 438184
rect 52454 438132 52460 438184
rect 52512 438172 52518 438184
rect 71314 438172 71320 438184
rect 52512 438144 71320 438172
rect 52512 438132 52518 438144
rect 71314 438132 71320 438144
rect 71372 438132 71378 438184
rect 85574 438132 85580 438184
rect 85632 438172 85638 438184
rect 118878 438172 118884 438184
rect 85632 438144 118884 438172
rect 85632 438132 85638 438144
rect 118878 438132 118884 438144
rect 118936 438132 118942 438184
rect 98362 437996 98368 438048
rect 98420 438036 98426 438048
rect 99282 438036 99288 438048
rect 98420 438008 99288 438036
rect 98420 437996 98426 438008
rect 99282 437996 99288 438008
rect 99340 438036 99346 438048
rect 102226 438036 102232 438048
rect 99340 438008 102232 438036
rect 99340 437996 99346 438008
rect 102226 437996 102232 438008
rect 102284 437996 102290 438048
rect 69106 437452 69112 437504
rect 69164 437492 69170 437504
rect 73246 437492 73252 437504
rect 69164 437464 73252 437492
rect 69164 437452 69170 437464
rect 73246 437452 73252 437464
rect 73304 437452 73310 437504
rect 85022 437452 85028 437504
rect 85080 437492 85086 437504
rect 86770 437492 86776 437504
rect 85080 437464 86776 437492
rect 85080 437452 85086 437464
rect 86770 437452 86776 437464
rect 86828 437452 86834 437504
rect 88058 437452 88064 437504
rect 88116 437492 88122 437504
rect 89622 437492 89628 437504
rect 88116 437464 89628 437492
rect 88116 437452 88122 437464
rect 89622 437452 89628 437464
rect 89680 437452 89686 437504
rect 47946 437384 47952 437436
rect 48004 437424 48010 437436
rect 78674 437424 78680 437436
rect 48004 437396 78680 437424
rect 48004 437384 48010 437396
rect 78674 437384 78680 437396
rect 78732 437424 78738 437436
rect 79042 437424 79048 437436
rect 78732 437396 79048 437424
rect 78732 437384 78738 437396
rect 79042 437384 79048 437396
rect 79100 437384 79106 437436
rect 89990 437384 89996 437436
rect 90048 437424 90054 437436
rect 90358 437424 90364 437436
rect 90048 437396 90364 437424
rect 90048 437384 90054 437396
rect 90358 437384 90364 437396
rect 90416 437424 90422 437436
rect 124398 437424 124404 437436
rect 90416 437396 124404 437424
rect 90416 437384 90422 437396
rect 124398 437384 124404 437396
rect 124456 437384 124462 437436
rect 39850 437316 39856 437368
rect 39908 437356 39914 437368
rect 69106 437356 69112 437368
rect 39908 437328 69112 437356
rect 39908 437316 39914 437328
rect 69106 437316 69112 437328
rect 69164 437316 69170 437368
rect 94958 437316 94964 437368
rect 95016 437356 95022 437368
rect 125778 437356 125784 437368
rect 95016 437328 125784 437356
rect 95016 437316 95022 437328
rect 125778 437316 125784 437328
rect 125836 437316 125842 437368
rect 37182 437248 37188 437300
rect 37240 437288 37246 437300
rect 52454 437288 52460 437300
rect 37240 437260 52460 437288
rect 37240 437248 37246 437260
rect 52454 437248 52460 437260
rect 52512 437288 52518 437300
rect 53098 437288 53104 437300
rect 52512 437260 53104 437288
rect 52512 437248 52518 437260
rect 53098 437248 53104 437260
rect 53156 437248 53162 437300
rect 53650 437248 53656 437300
rect 53708 437288 53714 437300
rect 74626 437288 74632 437300
rect 53708 437260 74632 437288
rect 53708 437248 53714 437260
rect 74626 437248 74632 437260
rect 74684 437288 74690 437300
rect 75822 437288 75828 437300
rect 74684 437260 75828 437288
rect 74684 437248 74690 437260
rect 75822 437248 75828 437260
rect 75880 437248 75886 437300
rect 89346 437248 89352 437300
rect 89404 437288 89410 437300
rect 89530 437288 89536 437300
rect 89404 437260 89536 437288
rect 89404 437248 89410 437260
rect 89530 437248 89536 437260
rect 89588 437288 89594 437300
rect 108390 437288 108396 437300
rect 89588 437260 108396 437288
rect 89588 437248 89594 437260
rect 108390 437248 108396 437260
rect 108448 437248 108454 437300
rect 54846 437180 54852 437232
rect 54904 437220 54910 437232
rect 70394 437220 70400 437232
rect 54904 437192 70400 437220
rect 54904 437180 54910 437192
rect 70394 437180 70400 437192
rect 70452 437180 70458 437232
rect 93210 437180 93216 437232
rect 93268 437220 93274 437232
rect 93670 437220 93676 437232
rect 93268 437192 93676 437220
rect 93268 437180 93274 437192
rect 93670 437180 93676 437192
rect 93728 437220 93734 437232
rect 108482 437220 108488 437232
rect 93728 437192 108488 437220
rect 93728 437180 93734 437192
rect 108482 437180 108488 437192
rect 108540 437180 108546 437232
rect 45462 437112 45468 437164
rect 45520 437152 45526 437164
rect 55858 437152 55864 437164
rect 45520 437124 55864 437152
rect 45520 437112 45526 437124
rect 55858 437112 55864 437124
rect 55916 437152 55922 437164
rect 56318 437152 56324 437164
rect 55916 437124 56324 437152
rect 55916 437112 55922 437124
rect 56318 437112 56324 437124
rect 56376 437112 56382 437164
rect 64506 436704 64512 436756
rect 64564 436744 64570 436756
rect 75178 436744 75184 436756
rect 64564 436716 75184 436744
rect 64564 436704 64570 436716
rect 75178 436704 75184 436716
rect 75236 436704 75242 436756
rect 59078 436024 59084 436076
rect 59136 436064 59142 436076
rect 91738 436064 91744 436076
rect 59136 436036 91744 436064
rect 59136 436024 59142 436036
rect 91738 436024 91744 436036
rect 91796 436024 91802 436076
rect 92566 436024 92572 436076
rect 92624 436064 92630 436076
rect 93762 436064 93768 436076
rect 92624 436036 93768 436064
rect 92624 436024 92630 436036
rect 93762 436024 93768 436036
rect 93820 436064 93826 436076
rect 124306 436064 124312 436076
rect 93820 436036 124312 436064
rect 93820 436024 93826 436036
rect 124306 436024 124312 436036
rect 124364 436024 124370 436076
rect 46842 435956 46848 436008
rect 46900 435996 46906 436008
rect 78582 435996 78588 436008
rect 46900 435968 78588 435996
rect 46900 435956 46906 435968
rect 78582 435956 78588 435968
rect 78640 435956 78646 436008
rect 89622 435956 89628 436008
rect 89680 435996 89686 436008
rect 112070 435996 112076 436008
rect 89680 435968 112076 435996
rect 89680 435956 89686 435968
rect 112070 435956 112076 435968
rect 112128 435956 112134 436008
rect 65518 435344 65524 435396
rect 65576 435384 65582 435396
rect 77938 435384 77944 435396
rect 65576 435356 77944 435384
rect 65576 435344 65582 435356
rect 77938 435344 77944 435356
rect 77996 435344 78002 435396
rect 41046 434664 41052 434716
rect 41104 434704 41110 434716
rect 41230 434704 41236 434716
rect 41104 434676 41236 434704
rect 41104 434664 41110 434676
rect 41230 434664 41236 434676
rect 41288 434664 41294 434716
rect 42518 434664 42524 434716
rect 42576 434704 42582 434716
rect 74534 434704 74540 434716
rect 42576 434676 74540 434704
rect 42576 434664 42582 434676
rect 74534 434664 74540 434676
rect 74592 434664 74598 434716
rect 41248 434636 41276 434664
rect 70670 434636 70676 434648
rect 41248 434608 70676 434636
rect 70670 434596 70676 434608
rect 70728 434596 70734 434648
rect 49326 434528 49332 434580
rect 49384 434568 49390 434580
rect 49602 434568 49608 434580
rect 49384 434540 49608 434568
rect 49384 434528 49390 434540
rect 49602 434528 49608 434540
rect 49660 434568 49666 434580
rect 76466 434568 76472 434580
rect 49660 434540 76472 434568
rect 49660 434528 49666 434540
rect 76466 434528 76472 434540
rect 76524 434528 76530 434580
rect 45278 433984 45284 434036
rect 45336 434024 45342 434036
rect 49602 434024 49608 434036
rect 45336 433996 49608 434024
rect 45336 433984 45342 433996
rect 49602 433984 49608 433996
rect 49660 433984 49666 434036
rect 78582 431944 78588 431996
rect 78640 431984 78646 431996
rect 80146 431984 80152 431996
rect 78640 431956 80152 431984
rect 78640 431944 78646 431956
rect 80146 431944 80152 431956
rect 80204 431984 80210 431996
rect 580902 431984 580908 431996
rect 80204 431956 580908 431984
rect 80204 431944 80210 431956
rect 580902 431944 580908 431956
rect 580960 431944 580966 431996
rect 39666 431876 39672 431928
rect 39724 431916 39730 431928
rect 71866 431916 71872 431928
rect 39724 431888 71872 431916
rect 39724 431876 39730 431888
rect 71866 431876 71872 431888
rect 71924 431876 71930 431928
rect 100754 430584 100760 430636
rect 100812 430624 100818 430636
rect 101950 430624 101956 430636
rect 100812 430596 101956 430624
rect 100812 430584 100818 430596
rect 101950 430584 101956 430596
rect 102008 430624 102014 430636
rect 104250 430624 104256 430636
rect 102008 430596 104256 430624
rect 102008 430584 102014 430596
rect 104250 430584 104256 430596
rect 104308 430584 104314 430636
rect 3418 429836 3424 429888
rect 3476 429876 3482 429888
rect 100754 429876 100760 429888
rect 3476 429848 100760 429876
rect 3476 429836 3482 429848
rect 100754 429836 100760 429848
rect 100812 429836 100818 429888
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 3568 422300 110184 422328
rect 3568 422288 3574 422300
rect 110156 422260 110184 422300
rect 118786 422260 118792 422272
rect 110156 422232 118792 422260
rect 118786 422220 118792 422232
rect 118844 422220 118850 422272
rect 121638 404336 121644 404388
rect 121696 404376 121702 404388
rect 579614 404376 579620 404388
rect 121696 404348 579620 404376
rect 121696 404336 121702 404348
rect 579614 404336 579620 404348
rect 579672 404336 579678 404388
rect 70394 404268 70400 404320
rect 70452 404308 70458 404320
rect 71038 404308 71044 404320
rect 70452 404280 71044 404308
rect 70452 404268 70458 404280
rect 71038 404268 71044 404280
rect 71096 404268 71102 404320
rect 93578 403656 93584 403708
rect 93636 403696 93642 403708
rect 129918 403696 129924 403708
rect 93636 403668 129924 403696
rect 93636 403656 93642 403668
rect 129918 403656 129924 403668
rect 129976 403656 129982 403708
rect 104158 403588 104164 403640
rect 104216 403628 104222 403640
rect 141050 403628 141056 403640
rect 104216 403600 141056 403628
rect 104216 403588 104222 403600
rect 141050 403588 141056 403600
rect 141108 403588 141114 403640
rect 70394 402976 70400 403028
rect 70452 403016 70458 403028
rect 341518 403016 341524 403028
rect 70452 402988 341524 403016
rect 70452 402976 70458 402988
rect 341518 402976 341524 402988
rect 341576 402976 341582 403028
rect 74810 401616 74816 401668
rect 74868 401656 74874 401668
rect 304258 401656 304264 401668
rect 74868 401628 304264 401656
rect 74868 401616 74874 401628
rect 304258 401616 304264 401628
rect 304316 401616 304322 401668
rect 96614 400868 96620 400920
rect 96672 400908 96678 400920
rect 132678 400908 132684 400920
rect 96672 400880 132684 400908
rect 96672 400868 96678 400880
rect 132678 400868 132684 400880
rect 132736 400868 132742 400920
rect 89530 399576 89536 399628
rect 89588 399616 89594 399628
rect 125962 399616 125968 399628
rect 89588 399588 125968 399616
rect 89588 399576 89594 399588
rect 125962 399576 125968 399588
rect 126020 399576 126026 399628
rect 41138 399508 41144 399560
rect 41196 399548 41202 399560
rect 86218 399548 86224 399560
rect 41196 399520 86224 399548
rect 41196 399508 41202 399520
rect 86218 399508 86224 399520
rect 86276 399508 86282 399560
rect 93670 399508 93676 399560
rect 93728 399548 93734 399560
rect 127250 399548 127256 399560
rect 93728 399520 127256 399548
rect 93728 399508 93734 399520
rect 127250 399508 127256 399520
rect 127308 399508 127314 399560
rect 39758 399440 39764 399492
rect 39816 399480 39822 399492
rect 85114 399480 85120 399492
rect 39816 399452 85120 399480
rect 39816 399440 39822 399452
rect 85114 399440 85120 399452
rect 85172 399440 85178 399492
rect 92658 399440 92664 399492
rect 92716 399480 92722 399492
rect 125870 399480 125876 399492
rect 92716 399452 125876 399480
rect 92716 399440 92722 399452
rect 125870 399440 125876 399452
rect 125928 399480 125934 399492
rect 197998 399480 198004 399492
rect 125928 399452 198004 399480
rect 125928 399440 125934 399452
rect 197998 399440 198004 399452
rect 198056 399440 198062 399492
rect 65978 398828 65984 398880
rect 66036 398868 66042 398880
rect 170398 398868 170404 398880
rect 66036 398840 170404 398868
rect 66036 398828 66042 398840
rect 170398 398828 170404 398840
rect 170456 398828 170462 398880
rect 100662 398760 100668 398812
rect 100720 398800 100726 398812
rect 104158 398800 104164 398812
rect 100720 398772 104164 398800
rect 100720 398760 100726 398772
rect 104158 398760 104164 398772
rect 104216 398760 104222 398812
rect 104250 398216 104256 398268
rect 104308 398256 104314 398268
rect 135438 398256 135444 398268
rect 104308 398228 135444 398256
rect 104308 398216 104314 398228
rect 135438 398216 135444 398228
rect 135496 398216 135502 398268
rect 97258 398148 97264 398200
rect 97316 398188 97322 398200
rect 130010 398188 130016 398200
rect 97316 398160 130016 398188
rect 97316 398148 97322 398160
rect 130010 398148 130016 398160
rect 130068 398148 130074 398200
rect 43990 398080 43996 398132
rect 44048 398120 44054 398132
rect 77294 398120 77300 398132
rect 44048 398092 77300 398120
rect 44048 398080 44054 398092
rect 77294 398080 77300 398092
rect 77352 398080 77358 398132
rect 91738 398080 91744 398132
rect 91796 398120 91802 398132
rect 128538 398120 128544 398132
rect 91796 398092 128544 398120
rect 91796 398080 91802 398092
rect 128538 398080 128544 398092
rect 128596 398080 128602 398132
rect 128354 397672 128360 397724
rect 128412 397712 128418 397724
rect 128722 397712 128728 397724
rect 128412 397684 128728 397712
rect 128412 397672 128418 397684
rect 128722 397672 128728 397684
rect 128780 397672 128786 397724
rect 128354 397536 128360 397588
rect 128412 397576 128418 397588
rect 128998 397576 129004 397588
rect 128412 397548 129004 397576
rect 128412 397536 128418 397548
rect 128998 397536 129004 397548
rect 129056 397576 129062 397588
rect 215938 397576 215944 397588
rect 129056 397548 215944 397576
rect 129056 397536 129062 397548
rect 215938 397536 215944 397548
rect 215996 397536 216002 397588
rect 61930 397468 61936 397520
rect 61988 397508 61994 397520
rect 291838 397508 291844 397520
rect 61988 397480 291844 397508
rect 61988 397468 61994 397480
rect 291838 397468 291844 397480
rect 291896 397468 291902 397520
rect 77938 397400 77944 397452
rect 77996 397440 78002 397452
rect 121638 397440 121644 397452
rect 77996 397412 121644 397440
rect 77996 397400 78002 397412
rect 121638 397400 121644 397412
rect 121696 397400 121702 397452
rect 56410 396896 56416 396908
rect 45526 396868 56416 396896
rect 39850 396788 39856 396840
rect 39908 396828 39914 396840
rect 45526 396828 45554 396868
rect 56410 396856 56416 396868
rect 56468 396896 56474 396908
rect 89714 396896 89720 396908
rect 56468 396868 89720 396896
rect 56468 396856 56474 396868
rect 89714 396856 89720 396868
rect 89772 396856 89778 396908
rect 93762 396856 93768 396908
rect 93820 396896 93826 396908
rect 128630 396896 128636 396908
rect 93820 396868 128636 396896
rect 93820 396856 93826 396868
rect 128630 396856 128636 396868
rect 128688 396856 128694 396908
rect 39908 396800 45554 396828
rect 39908 396788 39914 396800
rect 84102 396788 84108 396840
rect 84160 396828 84166 396840
rect 120810 396828 120816 396840
rect 84160 396800 120816 396828
rect 84160 396788 84166 396800
rect 120810 396788 120816 396800
rect 120868 396788 120874 396840
rect 42610 396720 42616 396772
rect 42668 396760 42674 396772
rect 88334 396760 88340 396772
rect 42668 396732 88340 396760
rect 42668 396720 42674 396732
rect 88334 396720 88340 396732
rect 88392 396720 88398 396772
rect 94130 396720 94136 396772
rect 94188 396760 94194 396772
rect 128354 396760 128360 396772
rect 94188 396732 128360 396760
rect 94188 396720 94194 396732
rect 128354 396720 128360 396732
rect 128412 396720 128418 396772
rect 88334 396040 88340 396092
rect 88392 396080 88398 396092
rect 195238 396080 195244 396092
rect 88392 396052 195244 396080
rect 88392 396040 88398 396052
rect 195238 396040 195244 396052
rect 195296 396040 195302 396092
rect 43898 395428 43904 395480
rect 43956 395468 43962 395480
rect 50982 395468 50988 395480
rect 43956 395440 50988 395468
rect 43956 395428 43962 395440
rect 50982 395428 50988 395440
rect 51040 395428 51046 395480
rect 59262 395428 59268 395480
rect 59320 395468 59326 395480
rect 84194 395468 84200 395480
rect 59320 395440 84200 395468
rect 59320 395428 59326 395440
rect 84194 395428 84200 395440
rect 84252 395428 84258 395480
rect 89714 395428 89720 395480
rect 89772 395468 89778 395480
rect 103790 395468 103796 395480
rect 89772 395440 103796 395468
rect 89772 395428 89778 395440
rect 103790 395428 103796 395440
rect 103848 395428 103854 395480
rect 43714 395360 43720 395412
rect 43772 395400 43778 395412
rect 82814 395400 82820 395412
rect 43772 395372 82820 395400
rect 43772 395360 43778 395372
rect 82814 395360 82820 395372
rect 82872 395360 82878 395412
rect 95142 395360 95148 395412
rect 95200 395400 95206 395412
rect 125778 395400 125784 395412
rect 95200 395372 125784 395400
rect 95200 395360 95206 395372
rect 125778 395360 125784 395372
rect 125836 395360 125842 395412
rect 38470 395292 38476 395344
rect 38528 395332 38534 395344
rect 81434 395332 81440 395344
rect 38528 395304 81440 395332
rect 38528 395292 38534 395304
rect 81434 395292 81440 395304
rect 81492 395292 81498 395344
rect 97994 395292 98000 395344
rect 98052 395332 98058 395344
rect 131298 395332 131304 395344
rect 98052 395304 131304 395332
rect 98052 395292 98058 395304
rect 131298 395292 131304 395304
rect 131356 395332 131362 395344
rect 322934 395332 322940 395344
rect 131356 395304 322940 395332
rect 131356 395292 131362 395304
rect 322934 395292 322940 395304
rect 322992 395292 322998 395344
rect 82814 394748 82820 394800
rect 82872 394788 82878 394800
rect 83090 394788 83096 394800
rect 82872 394760 83096 394788
rect 82872 394748 82878 394760
rect 83090 394748 83096 394760
rect 83148 394788 83154 394800
rect 139394 394788 139400 394800
rect 83148 394760 139400 394788
rect 83148 394748 83154 394760
rect 139394 394748 139400 394760
rect 139452 394748 139458 394800
rect 50982 394680 50988 394732
rect 51040 394720 51046 394732
rect 84194 394720 84200 394732
rect 51040 394692 84200 394720
rect 51040 394680 51046 394692
rect 84194 394680 84200 394692
rect 84252 394680 84258 394732
rect 103514 394680 103520 394732
rect 103572 394720 103578 394732
rect 104710 394720 104716 394732
rect 103572 394692 104716 394720
rect 103572 394680 103578 394692
rect 104710 394680 104716 394692
rect 104768 394720 104774 394732
rect 206278 394720 206284 394732
rect 104768 394692 206284 394720
rect 104768 394680 104774 394692
rect 206278 394680 206284 394692
rect 206336 394680 206342 394732
rect 109770 394612 109776 394664
rect 109828 394652 109834 394664
rect 111978 394652 111984 394664
rect 109828 394624 111984 394652
rect 109828 394612 109834 394624
rect 111978 394612 111984 394624
rect 112036 394612 112042 394664
rect 110874 394136 110880 394188
rect 110932 394176 110938 394188
rect 129734 394176 129740 394188
rect 110932 394148 129740 394176
rect 110932 394136 110938 394148
rect 129734 394136 129740 394148
rect 129792 394136 129798 394188
rect 93854 394068 93860 394120
rect 93912 394108 93918 394120
rect 128722 394108 128728 394120
rect 93912 394080 128728 394108
rect 93912 394068 93918 394080
rect 128722 394068 128728 394080
rect 128780 394068 128786 394120
rect 45370 394000 45376 394052
rect 45428 394040 45434 394052
rect 57606 394040 57612 394052
rect 45428 394012 57612 394040
rect 45428 394000 45434 394012
rect 57606 394000 57612 394012
rect 57664 394000 57670 394052
rect 96706 394000 96712 394052
rect 96764 394040 96770 394052
rect 131206 394040 131212 394052
rect 96764 394012 131212 394040
rect 96764 394000 96770 394012
rect 131206 394000 131212 394012
rect 131264 394040 131270 394052
rect 131264 394012 132494 394040
rect 131264 394000 131270 394012
rect 46566 393932 46572 393984
rect 46624 393972 46630 393984
rect 82906 393972 82912 393984
rect 46624 393944 82912 393972
rect 46624 393932 46630 393944
rect 82906 393932 82912 393944
rect 82964 393932 82970 393984
rect 88242 393932 88248 393984
rect 88300 393972 88306 393984
rect 124306 393972 124312 393984
rect 88300 393944 124312 393972
rect 88300 393932 88306 393944
rect 124306 393932 124312 393944
rect 124364 393932 124370 393984
rect 128722 393932 128728 393984
rect 128780 393972 128786 393984
rect 129734 393972 129740 393984
rect 128780 393944 129740 393972
rect 128780 393932 128786 393944
rect 129734 393932 129740 393944
rect 129792 393932 129798 393984
rect 132466 393972 132494 394012
rect 150434 393972 150440 393984
rect 132466 393944 150440 393972
rect 150434 393932 150440 393944
rect 150492 393932 150498 393984
rect 57606 393456 57612 393508
rect 57664 393496 57670 393508
rect 91094 393496 91100 393508
rect 57664 393468 91100 393496
rect 57664 393456 57670 393468
rect 91094 393456 91100 393468
rect 91152 393456 91158 393508
rect 39758 393388 39764 393440
rect 39816 393428 39822 393440
rect 110874 393428 110880 393440
rect 39816 393400 110880 393428
rect 39816 393388 39822 393400
rect 110874 393388 110880 393400
rect 110932 393388 110938 393440
rect 85114 393320 85120 393372
rect 85172 393360 85178 393372
rect 260098 393360 260104 393372
rect 85172 393332 260104 393360
rect 85172 393320 85178 393332
rect 260098 393320 260104 393332
rect 260156 393320 260162 393372
rect 105538 392776 105544 392828
rect 105596 392816 105602 392828
rect 117590 392816 117596 392828
rect 105596 392788 117596 392816
rect 105596 392776 105602 392788
rect 117590 392776 117596 392788
rect 117648 392776 117654 392828
rect 110322 392708 110328 392760
rect 110380 392748 110386 392760
rect 132494 392748 132500 392760
rect 110380 392720 132500 392748
rect 110380 392708 110386 392720
rect 132494 392708 132500 392720
rect 132552 392748 132558 392760
rect 136634 392748 136640 392760
rect 132552 392720 136640 392748
rect 132552 392708 132558 392720
rect 136634 392708 136640 392720
rect 136692 392708 136698 392760
rect 56410 392640 56416 392692
rect 56468 392680 56474 392692
rect 74534 392680 74540 392692
rect 56468 392652 74540 392680
rect 56468 392640 56474 392652
rect 74534 392640 74540 392652
rect 74592 392640 74598 392692
rect 96522 392640 96528 392692
rect 96580 392680 96586 392692
rect 123018 392680 123024 392692
rect 96580 392652 123024 392680
rect 96580 392640 96586 392652
rect 123018 392640 123024 392652
rect 123076 392640 123082 392692
rect 3418 392572 3424 392624
rect 3476 392612 3482 392624
rect 3476 392584 103514 392612
rect 3476 392572 3482 392584
rect 103486 392476 103514 392584
rect 116118 392476 116124 392488
rect 103486 392448 116124 392476
rect 116118 392436 116124 392448
rect 116176 392476 116182 392488
rect 118694 392476 118700 392488
rect 116176 392448 118700 392476
rect 116176 392436 116182 392448
rect 118694 392436 118700 392448
rect 118752 392436 118758 392488
rect 111058 392028 111064 392080
rect 111116 392068 111122 392080
rect 113634 392068 113640 392080
rect 111116 392040 113640 392068
rect 111116 392028 111122 392040
rect 113634 392028 113640 392040
rect 113692 392028 113698 392080
rect 67450 391960 67456 392012
rect 67508 392000 67514 392012
rect 298738 392000 298744 392012
rect 67508 391972 298744 392000
rect 67508 391960 67514 391972
rect 298738 391960 298744 391972
rect 298796 391960 298802 392012
rect 99282 391280 99288 391332
rect 99340 391320 99346 391332
rect 120166 391320 120172 391332
rect 99340 391292 120172 391320
rect 99340 391280 99346 391292
rect 120166 391280 120172 391292
rect 120224 391280 120230 391332
rect 53282 391212 53288 391264
rect 53340 391252 53346 391264
rect 75454 391252 75460 391264
rect 53340 391224 75460 391252
rect 53340 391212 53346 391224
rect 75454 391212 75460 391224
rect 75512 391212 75518 391264
rect 96522 391212 96528 391264
rect 96580 391252 96586 391264
rect 127158 391252 127164 391264
rect 96580 391224 127164 391252
rect 96580 391212 96586 391224
rect 127158 391212 127164 391224
rect 127216 391252 127222 391264
rect 142430 391252 142436 391264
rect 127216 391224 142436 391252
rect 127216 391212 127222 391224
rect 142430 391212 142436 391224
rect 142488 391212 142494 391264
rect 120074 390736 120080 390788
rect 120132 390776 120138 390788
rect 120718 390776 120724 390788
rect 120132 390748 120724 390776
rect 120132 390736 120138 390748
rect 120718 390736 120724 390748
rect 120776 390776 120782 390788
rect 127158 390776 127164 390788
rect 120776 390748 127164 390776
rect 120776 390736 120782 390748
rect 127158 390736 127164 390748
rect 127216 390736 127222 390788
rect 49602 390668 49608 390720
rect 49660 390708 49666 390720
rect 77938 390708 77944 390720
rect 49660 390680 77944 390708
rect 49660 390668 49666 390680
rect 77938 390668 77944 390680
rect 77996 390668 78002 390720
rect 81434 390668 81440 390720
rect 81492 390708 81498 390720
rect 82538 390708 82544 390720
rect 81492 390680 82544 390708
rect 81492 390668 81498 390680
rect 82538 390668 82544 390680
rect 82596 390708 82602 390720
rect 143718 390708 143724 390720
rect 82596 390680 143724 390708
rect 82596 390668 82602 390680
rect 143718 390668 143724 390680
rect 143776 390668 143782 390720
rect 75454 390600 75460 390652
rect 75512 390640 75518 390652
rect 140774 390640 140780 390652
rect 75512 390612 140780 390640
rect 75512 390600 75518 390612
rect 140774 390600 140780 390612
rect 140832 390600 140838 390652
rect 72418 390532 72424 390584
rect 72476 390572 72482 390584
rect 146570 390572 146576 390584
rect 72476 390544 146576 390572
rect 72476 390532 72482 390544
rect 146570 390532 146576 390544
rect 146628 390532 146634 390584
rect 58894 390056 58900 390108
rect 58952 390096 58958 390108
rect 104526 390096 104532 390108
rect 58952 390068 104532 390096
rect 58952 390056 58958 390068
rect 104526 390056 104532 390068
rect 104584 390056 104590 390108
rect 70302 389988 70308 390040
rect 70360 390028 70366 390040
rect 79318 390028 79324 390040
rect 70360 390000 79324 390028
rect 70360 389988 70366 390000
rect 79318 389988 79324 390000
rect 79376 389988 79382 390040
rect 69842 389920 69848 389972
rect 69900 389960 69906 389972
rect 85574 389960 85580 389972
rect 69900 389932 85580 389960
rect 69900 389920 69906 389932
rect 85574 389920 85580 389932
rect 85632 389920 85638 389972
rect 118786 389920 118792 389972
rect 118844 389960 118850 389972
rect 131206 389960 131212 389972
rect 118844 389932 131212 389960
rect 118844 389920 118850 389932
rect 131206 389920 131212 389932
rect 131264 389920 131270 389972
rect 57330 389852 57336 389904
rect 57388 389892 57394 389904
rect 120074 389892 120080 389904
rect 57388 389864 120080 389892
rect 57388 389852 57394 389864
rect 120074 389852 120080 389864
rect 120132 389852 120138 389904
rect 52178 389784 52184 389836
rect 52236 389824 52242 389836
rect 58894 389824 58900 389836
rect 52236 389796 58900 389824
rect 52236 389784 52242 389796
rect 58894 389784 58900 389796
rect 58952 389784 58958 389836
rect 99374 389784 99380 389836
rect 99432 389824 99438 389836
rect 111794 389824 111800 389836
rect 99432 389796 111800 389824
rect 99432 389784 99438 389796
rect 111794 389784 111800 389796
rect 111852 389824 111858 389836
rect 334710 389824 334716 389836
rect 111852 389796 334716 389824
rect 111852 389784 111858 389796
rect 334710 389784 334716 389796
rect 334768 389784 334774 389836
rect 111702 389580 111708 389632
rect 111760 389620 111766 389632
rect 114830 389620 114836 389632
rect 111760 389592 114836 389620
rect 111760 389580 111766 389592
rect 114830 389580 114836 389592
rect 114888 389580 114894 389632
rect 115566 389444 115572 389496
rect 115624 389484 115630 389496
rect 118786 389484 118792 389496
rect 115624 389456 118792 389484
rect 115624 389444 115630 389456
rect 118786 389444 118792 389456
rect 118844 389444 118850 389496
rect 101306 389308 101312 389360
rect 101364 389348 101370 389360
rect 133874 389348 133880 389360
rect 101364 389320 133880 389348
rect 101364 389308 101370 389320
rect 133874 389308 133880 389320
rect 133932 389308 133938 389360
rect 50798 389240 50804 389292
rect 50856 389280 50862 389292
rect 53742 389280 53748 389292
rect 50856 389252 53748 389280
rect 50856 389240 50862 389252
rect 53742 389240 53748 389252
rect 53800 389280 53806 389292
rect 79318 389280 79324 389292
rect 53800 389252 79324 389280
rect 53800 389240 53806 389252
rect 79318 389240 79324 389252
rect 79376 389240 79382 389292
rect 114278 389240 114284 389292
rect 114336 389280 114342 389292
rect 146478 389280 146484 389292
rect 114336 389252 146484 389280
rect 114336 389240 114342 389252
rect 146478 389240 146484 389252
rect 146536 389240 146542 389292
rect 42978 389172 42984 389224
rect 43036 389212 43042 389224
rect 43438 389212 43444 389224
rect 43036 389184 43444 389212
rect 43036 389172 43042 389184
rect 43438 389172 43444 389184
rect 43496 389212 43502 389224
rect 71774 389212 71780 389224
rect 43496 389184 71780 389212
rect 43496 389172 43502 389184
rect 71774 389172 71780 389184
rect 71832 389172 71838 389224
rect 113634 389172 113640 389224
rect 113692 389212 113698 389224
rect 262858 389212 262864 389224
rect 113692 389184 262864 389212
rect 113692 389172 113698 389184
rect 262858 389172 262864 389184
rect 262916 389172 262922 389224
rect 36630 389104 36636 389156
rect 36688 389144 36694 389156
rect 37090 389144 37096 389156
rect 36688 389116 37096 389144
rect 36688 389104 36694 389116
rect 37090 389104 37096 389116
rect 37148 389144 37154 389156
rect 72418 389144 72424 389156
rect 37148 389116 72424 389144
rect 37148 389104 37154 389116
rect 72418 389104 72424 389116
rect 72476 389104 72482 389156
rect 39942 389036 39948 389088
rect 40000 389076 40006 389088
rect 42978 389076 42984 389088
rect 40000 389048 42984 389076
rect 40000 389036 40006 389048
rect 42978 389036 42984 389048
rect 43036 389036 43042 389088
rect 90266 388560 90272 388612
rect 90324 388600 90330 388612
rect 99374 388600 99380 388612
rect 90324 388572 99380 388600
rect 90324 388560 90330 388572
rect 99374 388560 99380 388572
rect 99432 388560 99438 388612
rect 88242 388492 88248 388544
rect 88300 388532 88306 388544
rect 103514 388532 103520 388544
rect 88300 388504 103520 388532
rect 88300 388492 88306 388504
rect 103514 388492 103520 388504
rect 103572 388492 103578 388544
rect 107010 388492 107016 388544
rect 107068 388532 107074 388544
rect 135254 388532 135260 388544
rect 107068 388504 135260 388532
rect 107068 388492 107074 388504
rect 135254 388492 135260 388504
rect 135312 388532 135318 388544
rect 136542 388532 136548 388544
rect 135312 388504 136548 388532
rect 135312 388492 135318 388504
rect 136542 388492 136548 388504
rect 136600 388492 136606 388544
rect 4798 388424 4804 388476
rect 4856 388464 4862 388476
rect 36630 388464 36636 388476
rect 4856 388436 36636 388464
rect 4856 388424 4862 388436
rect 36630 388424 36636 388436
rect 36688 388424 36694 388476
rect 91002 388424 91008 388476
rect 91060 388464 91066 388476
rect 113082 388464 113088 388476
rect 91060 388436 113088 388464
rect 91060 388424 91066 388436
rect 113082 388424 113088 388436
rect 113140 388464 113146 388476
rect 313918 388464 313924 388476
rect 113140 388436 313924 388464
rect 113140 388424 113146 388436
rect 313918 388424 313924 388436
rect 313976 388424 313982 388476
rect 102594 388356 102600 388408
rect 102652 388396 102658 388408
rect 106182 388396 106188 388408
rect 102652 388368 106188 388396
rect 102652 388356 102658 388368
rect 106182 388356 106188 388368
rect 106240 388356 106246 388408
rect 73522 388084 73528 388136
rect 73580 388124 73586 388136
rect 73798 388124 73804 388136
rect 73580 388096 73804 388124
rect 73580 388084 73586 388096
rect 73798 388084 73804 388096
rect 73856 388124 73862 388136
rect 122190 388124 122196 388136
rect 73856 388096 122196 388124
rect 73856 388084 73862 388096
rect 122190 388084 122196 388096
rect 122248 388084 122254 388136
rect 109678 388016 109684 388068
rect 109736 388056 109742 388068
rect 119430 388056 119436 388068
rect 109736 388028 119436 388056
rect 109736 388016 109742 388028
rect 119430 388016 119436 388028
rect 119488 388016 119494 388068
rect 52270 387948 52276 388000
rect 52328 387988 52334 388000
rect 92934 387988 92940 388000
rect 52328 387960 92940 387988
rect 52328 387948 52334 387960
rect 92934 387948 92940 387960
rect 92992 387948 92998 388000
rect 101398 387948 101404 388000
rect 101456 387988 101462 388000
rect 119338 387988 119344 388000
rect 101456 387960 119344 387988
rect 101456 387948 101462 387960
rect 119338 387948 119344 387960
rect 119396 387948 119402 388000
rect 35526 387880 35532 387932
rect 35584 387920 35590 387932
rect 35710 387920 35716 387932
rect 35584 387892 35716 387920
rect 35584 387880 35590 387892
rect 35710 387880 35716 387892
rect 35768 387920 35774 387932
rect 80054 387920 80060 387932
rect 35768 387892 80060 387920
rect 35768 387880 35774 387892
rect 80054 387880 80060 387892
rect 80112 387880 80118 387932
rect 100018 387880 100024 387932
rect 100076 387920 100082 387932
rect 119522 387920 119528 387932
rect 100076 387892 119528 387920
rect 100076 387880 100082 387892
rect 119522 387880 119528 387892
rect 119580 387880 119586 387932
rect 58526 387812 58532 387864
rect 58584 387852 58590 387864
rect 70210 387852 70216 387864
rect 58584 387824 70216 387852
rect 58584 387812 58590 387824
rect 70210 387812 70216 387824
rect 70268 387812 70274 387864
rect 106182 387812 106188 387864
rect 106240 387852 106246 387864
rect 108758 387852 108764 387864
rect 106240 387824 108764 387852
rect 106240 387812 106246 387824
rect 108758 387812 108764 387824
rect 108816 387812 108822 387864
rect 69658 387336 69664 387388
rect 69716 387376 69722 387388
rect 78674 387376 78680 387388
rect 69716 387348 78680 387376
rect 69716 387336 69722 387348
rect 78674 387336 78680 387348
rect 78732 387336 78738 387388
rect 47946 387268 47952 387320
rect 48004 387308 48010 387320
rect 71866 387308 71872 387320
rect 48004 387280 71872 387308
rect 48004 387268 48010 387280
rect 71866 387268 71872 387280
rect 71924 387268 71930 387320
rect 52362 387200 52368 387252
rect 52420 387240 52426 387252
rect 80606 387240 80612 387252
rect 52420 387212 80612 387240
rect 52420 387200 52426 387212
rect 80606 387200 80612 387212
rect 80664 387200 80670 387252
rect 89622 387200 89628 387252
rect 89680 387240 89686 387252
rect 118694 387240 118700 387252
rect 89680 387212 118700 387240
rect 89680 387200 89686 387212
rect 118694 387200 118700 387212
rect 118752 387200 118758 387252
rect 59078 387132 59084 387184
rect 59136 387172 59142 387184
rect 90358 387172 90364 387184
rect 59136 387144 90364 387172
rect 59136 387132 59142 387144
rect 90358 387132 90364 387144
rect 90416 387132 90422 387184
rect 108298 387132 108304 387184
rect 108356 387172 108362 387184
rect 117406 387172 117412 387184
rect 108356 387144 117412 387172
rect 108356 387132 108362 387144
rect 117406 387132 117412 387144
rect 117464 387132 117470 387184
rect 60642 387064 60648 387116
rect 60700 387104 60706 387116
rect 95234 387104 95240 387116
rect 60700 387076 95240 387104
rect 60700 387064 60706 387076
rect 95234 387064 95240 387076
rect 95292 387064 95298 387116
rect 99282 387064 99288 387116
rect 99340 387104 99346 387116
rect 127342 387104 127348 387116
rect 99340 387076 127348 387104
rect 99340 387064 99346 387076
rect 127342 387064 127348 387076
rect 127400 387104 127406 387116
rect 127526 387104 127532 387116
rect 127400 387076 127532 387104
rect 127400 387064 127406 387076
rect 127526 387064 127532 387076
rect 127584 387064 127590 387116
rect 54938 386452 54944 386504
rect 54996 386492 55002 386504
rect 87046 386492 87052 386504
rect 54996 386464 87052 386492
rect 54996 386452 55002 386464
rect 87046 386452 87052 386464
rect 87104 386452 87110 386504
rect 103698 386452 103704 386504
rect 103756 386492 103762 386504
rect 104158 386492 104164 386504
rect 103756 386464 104164 386492
rect 103756 386452 103762 386464
rect 104158 386452 104164 386464
rect 104216 386492 104222 386504
rect 138198 386492 138204 386504
rect 104216 386464 138204 386492
rect 104216 386452 104222 386464
rect 138198 386452 138204 386464
rect 138256 386452 138262 386504
rect 76650 386384 76656 386436
rect 76708 386424 76714 386436
rect 327718 386424 327724 386436
rect 76708 386396 327724 386424
rect 76708 386384 76714 386396
rect 327718 386384 327724 386396
rect 327776 386384 327782 386436
rect 121362 386316 121368 386368
rect 121420 386356 121426 386368
rect 121546 386356 121552 386368
rect 121420 386328 121552 386356
rect 121420 386316 121426 386328
rect 121546 386316 121552 386328
rect 121604 386316 121610 386368
rect 66070 386248 66076 386300
rect 66128 386288 66134 386300
rect 68738 386288 68744 386300
rect 66128 386260 68744 386288
rect 66128 386248 66134 386260
rect 68738 386248 68744 386260
rect 68796 386248 68802 386300
rect 80146 386016 80152 386028
rect 64846 385988 80152 386016
rect 53558 385704 53564 385756
rect 53616 385744 53622 385756
rect 64846 385744 64874 385988
rect 80146 385976 80152 385988
rect 80204 385976 80210 386028
rect 53616 385716 64874 385744
rect 53616 385704 53622 385716
rect 105630 385704 105636 385756
rect 105688 385744 105694 385756
rect 131298 385744 131304 385756
rect 105688 385716 131304 385744
rect 105688 385704 105694 385716
rect 131298 385704 131304 385716
rect 131356 385704 131362 385756
rect 41322 385636 41328 385688
rect 41380 385676 41386 385688
rect 113358 385676 113364 385688
rect 41380 385648 113364 385676
rect 41380 385636 41386 385648
rect 113358 385636 113364 385648
rect 113416 385676 113422 385688
rect 117222 385676 117228 385688
rect 113416 385648 117228 385676
rect 113416 385636 113422 385648
rect 117222 385636 117228 385648
rect 117280 385636 117286 385688
rect 122282 385636 122288 385688
rect 122340 385676 122346 385688
rect 136910 385676 136916 385688
rect 122340 385648 136916 385676
rect 122340 385636 122346 385648
rect 136910 385636 136916 385648
rect 136968 385636 136974 385688
rect 112162 385364 112168 385416
rect 112220 385404 112226 385416
rect 112220 385376 122834 385404
rect 112220 385364 112226 385376
rect 107102 385336 107108 385348
rect 103486 385308 107108 385336
rect 52362 385024 52368 385076
rect 52420 385064 52426 385076
rect 103486 385064 103514 385308
rect 107102 385296 107108 385308
rect 107160 385296 107166 385348
rect 108942 385296 108948 385348
rect 109000 385336 109006 385348
rect 122098 385336 122104 385348
rect 109000 385308 122104 385336
rect 109000 385296 109006 385308
rect 122098 385296 122104 385308
rect 122156 385336 122162 385348
rect 122282 385336 122288 385348
rect 122156 385308 122288 385336
rect 122156 385296 122162 385308
rect 122282 385296 122288 385308
rect 122340 385296 122346 385348
rect 52420 385036 103514 385064
rect 122806 385064 122834 385376
rect 324958 385064 324964 385076
rect 122806 385036 324964 385064
rect 52420 385024 52426 385036
rect 324958 385024 324964 385036
rect 325016 385024 325022 385076
rect 116026 384344 116032 384396
rect 116084 384384 116090 384396
rect 122926 384384 122932 384396
rect 116084 384356 122932 384384
rect 116084 384344 116090 384356
rect 122926 384344 122932 384356
rect 122984 384344 122990 384396
rect 118602 384276 118608 384328
rect 118660 384316 118666 384328
rect 249058 384316 249064 384328
rect 118660 384288 249064 384316
rect 118660 384276 118666 384288
rect 249058 384276 249064 384288
rect 249116 384276 249122 384328
rect 34238 383664 34244 383716
rect 34296 383704 34302 383716
rect 68738 383704 68744 383716
rect 34296 383676 68744 383704
rect 34296 383664 34302 383676
rect 68738 383664 68744 383676
rect 68796 383664 68802 383716
rect 35802 382236 35808 382288
rect 35860 382276 35866 382288
rect 67634 382276 67640 382288
rect 35860 382248 67640 382276
rect 35860 382236 35866 382248
rect 67634 382236 67640 382248
rect 67692 382236 67698 382288
rect 116210 382236 116216 382288
rect 116268 382276 116274 382288
rect 145006 382276 145012 382288
rect 116268 382248 145012 382276
rect 116268 382236 116274 382248
rect 145006 382236 145012 382248
rect 145064 382236 145070 382288
rect 118602 382168 118608 382220
rect 118660 382208 118666 382220
rect 142338 382208 142344 382220
rect 118660 382180 142344 382208
rect 118660 382168 118666 382180
rect 142338 382168 142344 382180
rect 142396 382208 142402 382220
rect 143442 382208 143448 382220
rect 142396 382180 143448 382208
rect 142396 382168 142402 382180
rect 143442 382168 143448 382180
rect 143500 382168 143506 382220
rect 118602 381556 118608 381608
rect 118660 381596 118666 381608
rect 147674 381596 147680 381608
rect 118660 381568 147680 381596
rect 118660 381556 118666 381568
rect 147674 381556 147680 381568
rect 147732 381556 147738 381608
rect 143442 381488 143448 381540
rect 143500 381528 143506 381540
rect 204898 381528 204904 381540
rect 143500 381500 204904 381528
rect 143500 381488 143506 381500
rect 204898 381488 204904 381500
rect 204956 381488 204962 381540
rect 147674 380876 147680 380928
rect 147732 380916 147738 380928
rect 147950 380916 147956 380928
rect 147732 380888 147956 380916
rect 147732 380876 147738 380888
rect 147950 380876 147956 380888
rect 148008 380876 148014 380928
rect 42794 380808 42800 380860
rect 42852 380848 42858 380860
rect 44082 380848 44088 380860
rect 42852 380820 44088 380848
rect 42852 380808 42858 380820
rect 44082 380808 44088 380820
rect 44140 380848 44146 380860
rect 67634 380848 67640 380860
rect 44140 380820 67640 380848
rect 44140 380808 44146 380820
rect 67634 380808 67640 380820
rect 67692 380808 67698 380860
rect 60366 380740 60372 380792
rect 60424 380780 60430 380792
rect 68002 380780 68008 380792
rect 60424 380752 68008 380780
rect 60424 380740 60430 380752
rect 68002 380740 68008 380752
rect 68060 380740 68066 380792
rect 35618 380196 35624 380248
rect 35676 380236 35682 380248
rect 60182 380236 60188 380248
rect 35676 380208 60188 380236
rect 35676 380196 35682 380208
rect 60182 380196 60188 380208
rect 60240 380196 60246 380248
rect 18598 380128 18604 380180
rect 18656 380168 18662 380180
rect 42794 380168 42800 380180
rect 18656 380140 42800 380168
rect 18656 380128 18662 380140
rect 42794 380128 42800 380140
rect 42852 380128 42858 380180
rect 118602 379584 118608 379636
rect 118660 379624 118666 379636
rect 124490 379624 124496 379636
rect 118660 379596 124496 379624
rect 118660 379584 118666 379596
rect 124490 379584 124496 379596
rect 124548 379624 124554 379636
rect 128354 379624 128360 379636
rect 124548 379596 128360 379624
rect 124548 379584 124554 379596
rect 128354 379584 128360 379596
rect 128412 379584 128418 379636
rect 60182 379516 60188 379568
rect 60240 379556 60246 379568
rect 60458 379556 60464 379568
rect 60240 379528 60464 379556
rect 60240 379516 60246 379528
rect 60458 379516 60464 379528
rect 60516 379556 60522 379568
rect 67634 379556 67640 379568
rect 60516 379528 67640 379556
rect 60516 379516 60522 379528
rect 67634 379516 67640 379528
rect 67692 379516 67698 379568
rect 118510 379516 118516 379568
rect 118568 379556 118574 379568
rect 342898 379556 342904 379568
rect 118568 379528 342904 379556
rect 118568 379516 118574 379528
rect 342898 379516 342904 379528
rect 342956 379516 342962 379568
rect 118602 378836 118608 378888
rect 118660 378876 118666 378888
rect 123110 378876 123116 378888
rect 118660 378848 123116 378876
rect 118660 378836 118666 378848
rect 123110 378836 123116 378848
rect 123168 378836 123174 378888
rect 65150 378768 65156 378820
rect 65208 378808 65214 378820
rect 67634 378808 67640 378820
rect 65208 378780 67640 378808
rect 65208 378768 65214 378780
rect 67634 378768 67640 378780
rect 67692 378768 67698 378820
rect 119522 378768 119528 378820
rect 119580 378808 119586 378820
rect 346394 378808 346400 378820
rect 119580 378780 346400 378808
rect 119580 378768 119586 378780
rect 346394 378768 346400 378780
rect 346452 378768 346458 378820
rect 117866 378156 117872 378208
rect 117924 378196 117930 378208
rect 121546 378196 121552 378208
rect 117924 378168 121552 378196
rect 117924 378156 117930 378168
rect 121546 378156 121552 378168
rect 121604 378156 121610 378208
rect 121546 377544 121552 377596
rect 121604 377584 121610 377596
rect 125870 377584 125876 377596
rect 121604 377556 125876 377584
rect 121604 377544 121610 377556
rect 125870 377544 125876 377556
rect 125928 377544 125934 377596
rect 119522 377408 119528 377460
rect 119580 377448 119586 377460
rect 125686 377448 125692 377460
rect 119580 377420 125692 377448
rect 119580 377408 119586 377420
rect 125686 377408 125692 377420
rect 125744 377408 125750 377460
rect 118602 376796 118608 376848
rect 118660 376836 118666 376848
rect 119522 376836 119528 376848
rect 118660 376808 119528 376836
rect 118660 376796 118666 376808
rect 119522 376796 119528 376808
rect 119580 376796 119586 376848
rect 65518 376768 65524 376780
rect 64846 376740 65524 376768
rect 55030 376660 55036 376712
rect 55088 376700 55094 376712
rect 64846 376700 64874 376740
rect 65518 376728 65524 376740
rect 65576 376768 65582 376780
rect 67634 376768 67640 376780
rect 65576 376740 67640 376768
rect 65576 376728 65582 376740
rect 67634 376728 67640 376740
rect 67692 376728 67698 376780
rect 125870 376728 125876 376780
rect 125928 376768 125934 376780
rect 372614 376768 372620 376780
rect 125928 376740 372620 376768
rect 125928 376728 125934 376740
rect 372614 376728 372620 376740
rect 372672 376728 372678 376780
rect 55088 376672 64874 376700
rect 55088 376660 55094 376672
rect 149054 376660 149060 376712
rect 149112 376700 149118 376712
rect 150618 376700 150624 376712
rect 149112 376672 150624 376700
rect 149112 376660 149118 376672
rect 150618 376660 150624 376672
rect 150676 376660 150682 376712
rect 61930 376592 61936 376644
rect 61988 376632 61994 376644
rect 67634 376632 67640 376644
rect 61988 376604 67640 376632
rect 61988 376592 61994 376604
rect 67634 376592 67640 376604
rect 67692 376592 67698 376644
rect 55030 375980 55036 376032
rect 55088 376020 55094 376032
rect 70302 376020 70308 376032
rect 55088 375992 70308 376020
rect 55088 375980 55094 375992
rect 70302 375980 70308 375992
rect 70360 375980 70366 376032
rect 66990 375844 66996 375896
rect 67048 375884 67054 375896
rect 67634 375884 67640 375896
rect 67048 375856 67640 375884
rect 67048 375844 67054 375856
rect 67634 375844 67640 375856
rect 67692 375844 67698 375896
rect 118602 375368 118608 375420
rect 118660 375408 118666 375420
rect 149054 375408 149060 375420
rect 118660 375380 149060 375408
rect 118660 375368 118666 375380
rect 149054 375368 149060 375380
rect 149112 375368 149118 375420
rect 46658 375300 46664 375352
rect 46716 375340 46722 375352
rect 69106 375340 69112 375352
rect 46716 375312 69112 375340
rect 46716 375300 46722 375312
rect 69106 375300 69112 375312
rect 69164 375300 69170 375352
rect 118142 375300 118148 375352
rect 118200 375340 118206 375352
rect 147674 375340 147680 375352
rect 118200 375312 147680 375340
rect 118200 375300 118206 375312
rect 147674 375300 147680 375312
rect 147732 375340 147738 375352
rect 147858 375340 147864 375352
rect 147732 375312 147864 375340
rect 147732 375300 147738 375312
rect 147858 375300 147864 375312
rect 147916 375300 147922 375352
rect 63402 374620 63408 374672
rect 63460 374660 63466 374672
rect 67634 374660 67640 374672
rect 63460 374632 67640 374660
rect 63460 374620 63466 374632
rect 67634 374620 67640 374632
rect 67692 374620 67698 374672
rect 147674 374620 147680 374672
rect 147732 374660 147738 374672
rect 191098 374660 191104 374672
rect 147732 374632 191104 374660
rect 147732 374620 147738 374632
rect 191098 374620 191104 374632
rect 191156 374620 191162 374672
rect 58986 373940 58992 373992
rect 59044 373980 59050 373992
rect 67634 373980 67640 373992
rect 59044 373952 67640 373980
rect 59044 373940 59050 373952
rect 67634 373940 67640 373952
rect 67692 373940 67698 373992
rect 65978 373124 65984 373176
rect 66036 373164 66042 373176
rect 67634 373164 67640 373176
rect 66036 373136 67640 373164
rect 66036 373124 66042 373136
rect 67634 373124 67640 373136
rect 67692 373124 67698 373176
rect 118326 372648 118332 372700
rect 118384 372688 118390 372700
rect 120166 372688 120172 372700
rect 118384 372660 120172 372688
rect 118384 372648 118390 372660
rect 120166 372648 120172 372660
rect 120224 372648 120230 372700
rect 118510 372580 118516 372632
rect 118568 372620 118574 372632
rect 331858 372620 331864 372632
rect 118568 372592 331864 372620
rect 118568 372580 118574 372592
rect 331858 372580 331864 372592
rect 331916 372580 331922 372632
rect 3234 372512 3240 372564
rect 3292 372552 3298 372564
rect 57330 372552 57336 372564
rect 3292 372524 57336 372552
rect 3292 372512 3298 372524
rect 57330 372512 57336 372524
rect 57388 372512 57394 372564
rect 118142 371220 118148 371272
rect 118200 371260 118206 371272
rect 421558 371260 421564 371272
rect 118200 371232 421564 371260
rect 118200 371220 118206 371232
rect 421558 371220 421564 371232
rect 421616 371220 421622 371272
rect 120166 371152 120172 371204
rect 120224 371192 120230 371204
rect 151814 371192 151820 371204
rect 120224 371164 151820 371192
rect 120224 371152 120230 371164
rect 151814 371152 151820 371164
rect 151872 371192 151878 371204
rect 153102 371192 153108 371204
rect 151872 371164 153108 371192
rect 151872 371152 151878 371164
rect 153102 371152 153108 371164
rect 153160 371152 153166 371204
rect 64506 370608 64512 370660
rect 64564 370648 64570 370660
rect 67634 370648 67640 370660
rect 64564 370620 67640 370648
rect 64564 370608 64570 370620
rect 67634 370608 67640 370620
rect 67692 370608 67698 370660
rect 50338 370540 50344 370592
rect 50396 370580 50402 370592
rect 67266 370580 67272 370592
rect 50396 370552 67272 370580
rect 50396 370540 50402 370552
rect 67266 370540 67272 370552
rect 67324 370580 67330 370592
rect 67726 370580 67732 370592
rect 67324 370552 67732 370580
rect 67324 370540 67330 370552
rect 67726 370540 67732 370552
rect 67784 370540 67790 370592
rect 50798 370472 50804 370524
rect 50856 370512 50862 370524
rect 69750 370512 69756 370524
rect 50856 370484 69756 370512
rect 50856 370472 50862 370484
rect 69750 370472 69756 370484
rect 69808 370472 69814 370524
rect 115934 369928 115940 369980
rect 115992 369968 115998 369980
rect 120166 369968 120172 369980
rect 115992 369940 120172 369968
rect 115992 369928 115998 369940
rect 120166 369928 120172 369940
rect 120224 369928 120230 369980
rect 118142 369860 118148 369912
rect 118200 369900 118206 369912
rect 151814 369900 151820 369912
rect 118200 369872 151820 369900
rect 118200 369860 118206 369872
rect 151814 369860 151820 369872
rect 151872 369860 151878 369912
rect 57238 369112 57244 369164
rect 57296 369152 57302 369164
rect 67634 369152 67640 369164
rect 57296 369124 67640 369152
rect 57296 369112 57302 369124
rect 67634 369112 67640 369124
rect 67692 369112 67698 369164
rect 118602 368500 118608 368552
rect 118660 368540 118666 368552
rect 124398 368540 124404 368552
rect 118660 368512 124404 368540
rect 118660 368500 118666 368512
rect 124398 368500 124404 368512
rect 124456 368540 124462 368552
rect 128446 368540 128452 368552
rect 124456 368512 128452 368540
rect 124456 368500 124462 368512
rect 128446 368500 128452 368512
rect 128504 368500 128510 368552
rect 59170 367820 59176 367872
rect 59228 367860 59234 367872
rect 67910 367860 67916 367872
rect 59228 367832 67916 367860
rect 59228 367820 59234 367832
rect 67910 367820 67916 367832
rect 67968 367820 67974 367872
rect 118602 367820 118608 367872
rect 118660 367860 118666 367872
rect 121454 367860 121460 367872
rect 118660 367832 121460 367860
rect 118660 367820 118666 367832
rect 121454 367820 121460 367832
rect 121512 367860 121518 367872
rect 134518 367860 134524 367872
rect 121512 367832 134524 367860
rect 121512 367820 121518 367832
rect 134518 367820 134524 367832
rect 134576 367820 134582 367872
rect 58986 367752 58992 367804
rect 59044 367792 59050 367804
rect 69658 367792 69664 367804
rect 59044 367764 69664 367792
rect 59044 367752 59050 367764
rect 69658 367752 69664 367764
rect 69716 367752 69722 367804
rect 124122 367752 124128 367804
rect 124180 367792 124186 367804
rect 144914 367792 144920 367804
rect 124180 367764 144920 367792
rect 124180 367752 124186 367764
rect 144914 367752 144920 367764
rect 144972 367752 144978 367804
rect 479518 367752 479524 367804
rect 479576 367792 479582 367804
rect 579614 367792 579620 367804
rect 479576 367764 579620 367792
rect 479576 367752 479582 367764
rect 579614 367752 579620 367764
rect 579672 367752 579678 367804
rect 118602 367208 118608 367260
rect 118660 367248 118666 367260
rect 122926 367248 122932 367260
rect 118660 367220 122932 367248
rect 118660 367208 118666 367220
rect 122926 367208 122932 367220
rect 122984 367248 122990 367260
rect 124122 367248 124128 367260
rect 122984 367220 124128 367248
rect 122984 367208 122990 367220
rect 124122 367208 124128 367220
rect 124180 367208 124186 367260
rect 48222 367004 48228 367056
rect 48280 367044 48286 367056
rect 60182 367044 60188 367056
rect 48280 367016 60188 367044
rect 48280 367004 48286 367016
rect 60182 367004 60188 367016
rect 60240 367004 60246 367056
rect 120166 367004 120172 367056
rect 120224 367044 120230 367056
rect 137002 367044 137008 367056
rect 120224 367016 137008 367044
rect 120224 367004 120230 367016
rect 137002 367004 137008 367016
rect 137060 367044 137066 367056
rect 137186 367044 137192 367056
rect 137060 367016 137192 367044
rect 137060 367004 137066 367016
rect 137186 367004 137192 367016
rect 137244 367004 137250 367056
rect 64598 366392 64604 366444
rect 64656 366432 64662 366444
rect 68462 366432 68468 366444
rect 64656 366404 68468 366432
rect 64656 366392 64662 366404
rect 68462 366392 68468 366404
rect 68520 366392 68526 366444
rect 118602 366392 118608 366444
rect 118660 366432 118666 366444
rect 143534 366432 143540 366444
rect 118660 366404 143540 366432
rect 118660 366392 118666 366404
rect 143534 366392 143540 366404
rect 143592 366392 143598 366444
rect 60182 366324 60188 366376
rect 60240 366364 60246 366376
rect 67634 366364 67640 366376
rect 60240 366336 67640 366364
rect 60240 366324 60246 366336
rect 67634 366324 67640 366336
rect 67692 366324 67698 366376
rect 137186 366324 137192 366376
rect 137244 366364 137250 366376
rect 579614 366364 579620 366376
rect 137244 366336 579620 366364
rect 137244 366324 137250 366336
rect 579614 366324 579620 366336
rect 579672 366324 579678 366376
rect 60550 365752 60556 365764
rect 41248 365724 60556 365752
rect 37182 365644 37188 365696
rect 37240 365684 37246 365696
rect 40954 365684 40960 365696
rect 37240 365656 40960 365684
rect 37240 365644 37246 365656
rect 40954 365644 40960 365656
rect 41012 365684 41018 365696
rect 41248 365684 41276 365724
rect 60550 365712 60556 365724
rect 60608 365712 60614 365764
rect 41012 365656 41276 365684
rect 41012 365644 41018 365656
rect 120810 365644 120816 365696
rect 120868 365684 120874 365696
rect 121454 365684 121460 365696
rect 120868 365656 121460 365684
rect 120868 365644 120874 365656
rect 121454 365644 121460 365656
rect 121512 365644 121518 365696
rect 118602 365032 118608 365084
rect 118660 365072 118666 365084
rect 132586 365072 132592 365084
rect 118660 365044 132592 365072
rect 118660 365032 118666 365044
rect 132586 365032 132592 365044
rect 132644 365032 132650 365084
rect 63126 364964 63132 365016
rect 63184 365004 63190 365016
rect 68554 365004 68560 365016
rect 63184 364976 68560 365004
rect 63184 364964 63190 364976
rect 68554 364964 68560 364976
rect 68612 364964 68618 365016
rect 120718 364964 120724 365016
rect 120776 365004 120782 365016
rect 146294 365004 146300 365016
rect 120776 364976 146300 365004
rect 120776 364964 120782 364976
rect 146294 364964 146300 364976
rect 146352 364964 146358 365016
rect 118510 364352 118516 364404
rect 118568 364392 118574 364404
rect 120718 364392 120724 364404
rect 118568 364364 120724 364392
rect 118568 364352 118574 364364
rect 120718 364352 120724 364364
rect 120776 364352 120782 364404
rect 121454 364352 121460 364404
rect 121512 364392 121518 364404
rect 579798 364392 579804 364404
rect 121512 364364 579804 364392
rect 121512 364352 121518 364364
rect 579798 364352 579804 364364
rect 579856 364352 579862 364404
rect 60550 364284 60556 364336
rect 60608 364324 60614 364336
rect 67726 364324 67732 364336
rect 60608 364296 67732 364324
rect 60608 364284 60614 364296
rect 67726 364284 67732 364296
rect 67784 364284 67790 364336
rect 48038 363604 48044 363656
rect 48096 363644 48102 363656
rect 67634 363644 67640 363656
rect 48096 363616 67640 363644
rect 48096 363604 48102 363616
rect 67634 363604 67640 363616
rect 67692 363604 67698 363656
rect 117406 363604 117412 363656
rect 117464 363644 117470 363656
rect 282178 363644 282184 363656
rect 117464 363616 282184 363644
rect 117464 363604 117470 363616
rect 282178 363604 282184 363616
rect 282236 363604 282242 363656
rect 48038 363060 48044 363112
rect 48096 363100 48102 363112
rect 48222 363100 48228 363112
rect 48096 363072 48228 363100
rect 48096 363060 48102 363072
rect 48222 363060 48228 363072
rect 48280 363060 48286 363112
rect 118602 362856 118608 362908
rect 118660 362896 118666 362908
rect 143626 362896 143632 362908
rect 118660 362868 143632 362896
rect 118660 362856 118666 362868
rect 143626 362856 143632 362868
rect 143684 362896 143690 362908
rect 144822 362896 144828 362908
rect 143684 362868 144828 362896
rect 143684 362856 143690 362868
rect 144822 362856 144828 362868
rect 144880 362856 144886 362908
rect 118602 362176 118608 362228
rect 118660 362216 118666 362228
rect 119982 362216 119988 362228
rect 118660 362188 119988 362216
rect 118660 362176 118666 362188
rect 119982 362176 119988 362188
rect 120040 362216 120046 362228
rect 134058 362216 134064 362228
rect 120040 362188 134064 362216
rect 120040 362176 120046 362188
rect 134058 362176 134064 362188
rect 134116 362176 134122 362228
rect 144822 362176 144828 362228
rect 144880 362216 144886 362228
rect 202138 362216 202144 362228
rect 144880 362188 202144 362216
rect 144880 362176 144886 362188
rect 202138 362176 202144 362188
rect 202196 362176 202202 362228
rect 116578 361972 116584 362024
rect 116636 362012 116642 362024
rect 117314 362012 117320 362024
rect 116636 361984 117320 362012
rect 116636 361972 116642 361984
rect 117314 361972 117320 361984
rect 117372 361972 117378 362024
rect 36538 361604 36544 361616
rect 35866 361576 36544 361604
rect 32950 361496 32956 361548
rect 33008 361536 33014 361548
rect 35866 361536 35894 361576
rect 36538 361564 36544 361576
rect 36596 361604 36602 361616
rect 36596 361576 60780 361604
rect 36596 361564 36602 361576
rect 33008 361508 35894 361536
rect 60752 361536 60780 361576
rect 67634 361536 67640 361548
rect 60752 361508 67640 361536
rect 33008 361496 33014 361508
rect 67634 361496 67640 361508
rect 67692 361496 67698 361548
rect 44818 360816 44824 360868
rect 44876 360856 44882 360868
rect 45462 360856 45468 360868
rect 44876 360828 45468 360856
rect 44876 360816 44882 360828
rect 45462 360816 45468 360828
rect 45520 360856 45526 360868
rect 67634 360856 67640 360868
rect 45520 360828 67640 360856
rect 45520 360816 45526 360828
rect 67634 360816 67640 360828
rect 67692 360816 67698 360868
rect 125502 360272 125508 360324
rect 125560 360312 125566 360324
rect 128446 360312 128452 360324
rect 125560 360284 128452 360312
rect 125560 360272 125566 360284
rect 128446 360272 128452 360284
rect 128504 360272 128510 360324
rect 118050 360204 118056 360256
rect 118108 360244 118114 360256
rect 135898 360244 135904 360256
rect 118108 360216 135904 360244
rect 118108 360204 118114 360216
rect 135898 360204 135904 360216
rect 135956 360244 135962 360256
rect 139486 360244 139492 360256
rect 135956 360216 139492 360244
rect 135956 360204 135962 360216
rect 139486 360204 139492 360216
rect 139544 360204 139550 360256
rect 117958 360136 117964 360188
rect 118016 360176 118022 360188
rect 151998 360176 152004 360188
rect 118016 360148 152004 360176
rect 118016 360136 118022 360148
rect 151998 360136 152004 360148
rect 152056 360176 152062 360188
rect 153102 360176 153108 360188
rect 152056 360148 153108 360176
rect 152056 360136 152062 360148
rect 153102 360136 153108 360148
rect 153160 360136 153166 360188
rect 118602 360068 118608 360120
rect 118660 360108 118666 360120
rect 125502 360108 125508 360120
rect 118660 360080 125508 360108
rect 118660 360068 118666 360080
rect 125502 360068 125508 360080
rect 125560 360068 125566 360120
rect 68554 359524 68560 359576
rect 68612 359564 68618 359576
rect 68922 359564 68928 359576
rect 68612 359536 68928 359564
rect 68612 359524 68618 359536
rect 68922 359524 68928 359536
rect 68980 359524 68986 359576
rect 53190 359456 53196 359508
rect 53248 359496 53254 359508
rect 53650 359496 53656 359508
rect 53248 359468 53656 359496
rect 53248 359456 53254 359468
rect 53650 359456 53656 359468
rect 53708 359496 53714 359508
rect 67634 359496 67640 359508
rect 53708 359468 67640 359496
rect 53708 359456 53714 359468
rect 67634 359456 67640 359468
rect 67692 359456 67698 359508
rect 68462 359456 68468 359508
rect 68520 359496 68526 359508
rect 68830 359496 68836 359508
rect 68520 359468 68836 359496
rect 68520 359456 68526 359468
rect 68830 359456 68836 359468
rect 68888 359456 68894 359508
rect 153102 359456 153108 359508
rect 153160 359496 153166 359508
rect 188338 359496 188344 359508
rect 153160 359468 188344 359496
rect 153160 359456 153166 359468
rect 188338 359456 188344 359468
rect 188396 359456 188402 359508
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 36998 358748 37004 358760
rect 3384 358720 37004 358748
rect 3384 358708 3390 358720
rect 36998 358708 37004 358720
rect 37056 358748 37062 358760
rect 43530 358748 43536 358760
rect 37056 358720 43536 358748
rect 37056 358708 37062 358720
rect 43530 358708 43536 358720
rect 43588 358708 43594 358760
rect 56502 358708 56508 358760
rect 56560 358748 56566 358760
rect 59354 358748 59360 358760
rect 56560 358720 59360 358748
rect 56560 358708 56566 358720
rect 59354 358708 59360 358720
rect 59412 358708 59418 358760
rect 118602 358708 118608 358760
rect 118660 358748 118666 358760
rect 127158 358748 127164 358760
rect 118660 358720 127164 358748
rect 118660 358708 118666 358720
rect 127158 358708 127164 358720
rect 127216 358748 127222 358760
rect 129826 358748 129832 358760
rect 127216 358720 129832 358748
rect 127216 358708 127222 358720
rect 129826 358708 129832 358720
rect 129884 358708 129890 358760
rect 30282 358028 30288 358080
rect 30340 358068 30346 358080
rect 65978 358068 65984 358080
rect 30340 358040 65984 358068
rect 30340 358028 30346 358040
rect 65978 358028 65984 358040
rect 66036 358068 66042 358080
rect 67634 358068 67640 358080
rect 66036 358040 67640 358068
rect 66036 358028 66042 358040
rect 67634 358028 67640 358040
rect 67692 358028 67698 358080
rect 59354 357416 59360 357468
rect 59412 357456 59418 357468
rect 67634 357456 67640 357468
rect 59412 357428 67640 357456
rect 59412 357416 59418 357428
rect 67634 357416 67640 357428
rect 67692 357416 67698 357468
rect 115842 357348 115848 357400
rect 115900 357388 115906 357400
rect 117406 357388 117412 357400
rect 115900 357360 117412 357388
rect 115900 357348 115906 357360
rect 117406 357348 117412 357360
rect 117464 357348 117470 357400
rect 118602 357348 118608 357400
rect 118660 357388 118666 357400
rect 138106 357388 138112 357400
rect 118660 357360 138112 357388
rect 118660 357348 118666 357360
rect 138106 357348 138112 357360
rect 138164 357388 138170 357400
rect 140866 357388 140872 357400
rect 138164 357360 140872 357388
rect 138164 357348 138170 357360
rect 140866 357348 140872 357360
rect 140924 357348 140930 357400
rect 42702 356668 42708 356720
rect 42760 356708 42766 356720
rect 67634 356708 67640 356720
rect 42760 356680 67640 356708
rect 42760 356668 42766 356680
rect 67634 356668 67640 356680
rect 67692 356668 67698 356720
rect 118234 356668 118240 356720
rect 118292 356708 118298 356720
rect 340138 356708 340144 356720
rect 118292 356680 340144 356708
rect 118292 356668 118298 356680
rect 340138 356668 340144 356680
rect 340196 356668 340202 356720
rect 61488 356068 64874 356096
rect 61488 356040 61516 356068
rect 55122 355988 55128 356040
rect 55180 356028 55186 356040
rect 61470 356028 61476 356040
rect 55180 356000 61476 356028
rect 55180 355988 55186 356000
rect 61470 355988 61476 356000
rect 61528 355988 61534 356040
rect 64846 356028 64874 356068
rect 67634 356028 67640 356040
rect 64846 356000 67640 356028
rect 67634 355988 67640 356000
rect 67692 355988 67698 356040
rect 52086 355308 52092 355360
rect 52144 355348 52150 355360
rect 59170 355348 59176 355360
rect 52144 355320 59176 355348
rect 52144 355308 52150 355320
rect 59170 355308 59176 355320
rect 59228 355308 59234 355360
rect 119338 355308 119344 355360
rect 119396 355348 119402 355360
rect 580258 355348 580264 355360
rect 119396 355320 580264 355348
rect 119396 355308 119402 355320
rect 580258 355308 580264 355320
rect 580316 355308 580322 355360
rect 59170 354696 59176 354748
rect 59228 354736 59234 354748
rect 67634 354736 67640 354748
rect 59228 354708 67640 354736
rect 59228 354696 59234 354708
rect 67634 354696 67640 354708
rect 67692 354696 67698 354748
rect 118602 354628 118608 354680
rect 118660 354668 118666 354680
rect 140958 354668 140964 354680
rect 118660 354640 140964 354668
rect 118660 354628 118666 354640
rect 140958 354628 140964 354640
rect 141016 354628 141022 354680
rect 117498 354560 117504 354612
rect 117556 354600 117562 354612
rect 125594 354600 125600 354612
rect 117556 354572 125600 354600
rect 117556 354560 117562 354572
rect 125594 354560 125600 354572
rect 125652 354560 125658 354612
rect 140958 354016 140964 354068
rect 141016 354056 141022 354068
rect 147674 354056 147680 354068
rect 141016 354028 147680 354056
rect 141016 354016 141022 354028
rect 147674 354016 147680 354028
rect 147732 354016 147738 354068
rect 118786 353948 118792 354000
rect 118844 353988 118850 354000
rect 297358 353988 297364 354000
rect 118844 353960 297364 353988
rect 118844 353948 118850 353960
rect 297358 353948 297364 353960
rect 297416 353948 297422 354000
rect 125594 353268 125600 353320
rect 125652 353308 125658 353320
rect 126974 353308 126980 353320
rect 125652 353280 126980 353308
rect 125652 353268 125658 353280
rect 126974 353268 126980 353280
rect 127032 353268 127038 353320
rect 146294 353308 146300 353320
rect 135180 353280 146300 353308
rect 117498 353200 117504 353252
rect 117556 353240 117562 353252
rect 134058 353240 134064 353252
rect 117556 353212 134064 353240
rect 117556 353200 117562 353212
rect 134058 353200 134064 353212
rect 134116 353240 134122 353252
rect 135180 353240 135208 353280
rect 146294 353268 146300 353280
rect 146352 353268 146358 353320
rect 134116 353212 135208 353240
rect 134116 353200 134122 353212
rect 64782 352588 64788 352640
rect 64840 352628 64846 352640
rect 67634 352628 67640 352640
rect 64840 352600 67640 352628
rect 64840 352588 64846 352600
rect 67634 352588 67640 352600
rect 67692 352588 67698 352640
rect 7558 352520 7564 352572
rect 7616 352560 7622 352572
rect 68554 352560 68560 352572
rect 7616 352532 68560 352560
rect 7616 352520 7622 352532
rect 68554 352520 68560 352532
rect 68612 352520 68618 352572
rect 482278 352520 482284 352572
rect 482336 352560 482342 352572
rect 579614 352560 579620 352572
rect 482336 352532 579620 352560
rect 482336 352520 482342 352532
rect 579614 352520 579620 352532
rect 579672 352520 579678 352572
rect 118050 351840 118056 351892
rect 118108 351880 118114 351892
rect 138014 351880 138020 351892
rect 118108 351852 138020 351880
rect 118108 351840 118114 351852
rect 138014 351840 138020 351852
rect 138072 351840 138078 351892
rect 138014 351228 138020 351280
rect 138072 351268 138078 351280
rect 196618 351268 196624 351280
rect 138072 351240 196624 351268
rect 138072 351228 138078 351240
rect 196618 351228 196624 351240
rect 196676 351228 196682 351280
rect 64690 351160 64696 351212
rect 64748 351200 64754 351212
rect 68002 351200 68008 351212
rect 64748 351172 68008 351200
rect 64748 351160 64754 351172
rect 68002 351160 68008 351172
rect 68060 351160 68066 351212
rect 118602 351160 118608 351212
rect 118660 351200 118666 351212
rect 318058 351200 318064 351212
rect 118660 351172 318064 351200
rect 118660 351160 118666 351172
rect 318058 351160 318064 351172
rect 318116 351160 318122 351212
rect 49418 350548 49424 350600
rect 49476 350588 49482 350600
rect 53834 350588 53840 350600
rect 49476 350560 53840 350588
rect 49476 350548 49482 350560
rect 53834 350548 53840 350560
rect 53892 350548 53898 350600
rect 53834 349800 53840 349852
rect 53892 349840 53898 349852
rect 55122 349840 55128 349852
rect 53892 349812 55128 349840
rect 53892 349800 53898 349812
rect 55122 349800 55128 349812
rect 55180 349840 55186 349852
rect 67634 349840 67640 349852
rect 55180 349812 67640 349840
rect 55180 349800 55186 349812
rect 67634 349800 67640 349812
rect 67692 349800 67698 349852
rect 122190 349800 122196 349852
rect 122248 349840 122254 349852
rect 346486 349840 346492 349852
rect 122248 349812 346492 349840
rect 122248 349800 122254 349812
rect 346486 349800 346492 349812
rect 346544 349800 346550 349852
rect 61378 349120 61384 349172
rect 61436 349160 61442 349172
rect 64414 349160 64420 349172
rect 61436 349132 64420 349160
rect 61436 349120 61442 349132
rect 64414 349120 64420 349132
rect 64472 349160 64478 349172
rect 67634 349160 67640 349172
rect 64472 349132 67640 349160
rect 64472 349120 64478 349132
rect 67634 349120 67640 349132
rect 67692 349120 67698 349172
rect 117498 349120 117504 349172
rect 117556 349160 117562 349172
rect 119430 349160 119436 349172
rect 117556 349132 119436 349160
rect 117556 349120 117562 349132
rect 119430 349120 119436 349132
rect 119488 349120 119494 349172
rect 46842 349052 46848 349104
rect 46900 349092 46906 349104
rect 48130 349092 48136 349104
rect 46900 349064 48136 349092
rect 46900 349052 46906 349064
rect 48130 349052 48136 349064
rect 48188 349052 48194 349104
rect 63218 348440 63224 348492
rect 63276 348480 63282 348492
rect 67634 348480 67640 348492
rect 63276 348452 67640 348480
rect 63276 348440 63282 348452
rect 67634 348440 67640 348452
rect 67692 348440 67698 348492
rect 48130 348372 48136 348424
rect 48188 348412 48194 348424
rect 63494 348412 63500 348424
rect 48188 348384 63500 348412
rect 48188 348372 48194 348384
rect 63494 348372 63500 348384
rect 63552 348372 63558 348424
rect 118510 348372 118516 348424
rect 118568 348412 118574 348424
rect 320818 348412 320824 348424
rect 118568 348384 320824 348412
rect 118568 348372 118574 348384
rect 320818 348372 320824 348384
rect 320876 348372 320882 348424
rect 63494 347692 63500 347744
rect 63552 347732 63558 347744
rect 67634 347732 67640 347744
rect 63552 347704 67640 347732
rect 63552 347692 63558 347704
rect 67634 347692 67640 347704
rect 67692 347692 67698 347744
rect 118602 347692 118608 347744
rect 118660 347732 118666 347744
rect 151906 347732 151912 347744
rect 118660 347704 151912 347732
rect 118660 347692 118666 347704
rect 151906 347692 151912 347704
rect 151964 347732 151970 347744
rect 153102 347732 153108 347744
rect 151964 347704 153108 347732
rect 151964 347692 151970 347704
rect 153102 347692 153108 347704
rect 153160 347692 153166 347744
rect 153102 347012 153108 347064
rect 153160 347052 153166 347064
rect 184198 347052 184204 347064
rect 153160 347024 184204 347052
rect 153160 347012 153166 347024
rect 184198 347012 184204 347024
rect 184256 347012 184262 347064
rect 118602 346332 118608 346384
rect 118660 346372 118666 346384
rect 135346 346372 135352 346384
rect 118660 346344 135352 346372
rect 118660 346332 118666 346344
rect 135346 346332 135352 346344
rect 135404 346372 135410 346384
rect 136542 346372 136548 346384
rect 135404 346344 136548 346372
rect 135404 346332 135410 346344
rect 136542 346332 136548 346344
rect 136600 346332 136606 346384
rect 2774 346264 2780 346316
rect 2832 346304 2838 346316
rect 4798 346304 4804 346316
rect 2832 346276 4804 346304
rect 2832 346264 2838 346276
rect 4798 346264 4804 346276
rect 4856 346264 4862 346316
rect 118510 345720 118516 345772
rect 118568 345760 118574 345772
rect 142246 345760 142252 345772
rect 118568 345732 142252 345760
rect 118568 345720 118574 345732
rect 142246 345720 142252 345732
rect 142304 345720 142310 345772
rect 43530 345652 43536 345704
rect 43588 345692 43594 345704
rect 61930 345692 61936 345704
rect 43588 345664 61936 345692
rect 43588 345652 43594 345664
rect 61930 345652 61936 345664
rect 61988 345652 61994 345704
rect 136542 345652 136548 345704
rect 136600 345692 136606 345704
rect 186958 345692 186964 345704
rect 136600 345664 186964 345692
rect 136600 345652 136606 345664
rect 186958 345652 186964 345664
rect 187016 345652 187022 345704
rect 61930 345108 61936 345160
rect 61988 345148 61994 345160
rect 67634 345148 67640 345160
rect 61988 345120 67640 345148
rect 61988 345108 61994 345120
rect 67634 345108 67640 345120
rect 67692 345108 67698 345160
rect 56318 345040 56324 345092
rect 56376 345080 56382 345092
rect 67082 345080 67088 345092
rect 56376 345052 67088 345080
rect 56376 345040 56382 345052
rect 67082 345040 67088 345052
rect 67140 345080 67146 345092
rect 67140 345052 67634 345080
rect 67140 345040 67146 345052
rect 67606 345012 67634 345052
rect 68002 345012 68008 345024
rect 67606 344984 68008 345012
rect 68002 344972 68008 344984
rect 68060 344972 68066 345024
rect 117958 344972 117964 345024
rect 118016 345012 118022 345024
rect 149238 345012 149244 345024
rect 118016 344984 149244 345012
rect 118016 344972 118022 344984
rect 149238 344972 149244 344984
rect 149296 344972 149302 345024
rect 149238 344292 149244 344344
rect 149296 344332 149302 344344
rect 349890 344332 349896 344344
rect 149296 344304 349896 344332
rect 149296 344292 149302 344304
rect 349890 344292 349896 344304
rect 349948 344292 349954 344344
rect 62114 343612 62120 343664
rect 62172 343652 62178 343664
rect 67634 343652 67640 343664
rect 62172 343624 67640 343652
rect 62172 343612 62178 343624
rect 67634 343612 67640 343624
rect 67692 343612 67698 343664
rect 117866 343612 117872 343664
rect 117924 343652 117930 343664
rect 244918 343652 244924 343664
rect 117924 343624 244924 343652
rect 117924 343612 117930 343624
rect 244918 343612 244924 343624
rect 244976 343612 244982 343664
rect 34330 342864 34336 342916
rect 34388 342904 34394 342916
rect 41138 342904 41144 342916
rect 34388 342876 41144 342904
rect 34388 342864 34394 342876
rect 41138 342864 41144 342876
rect 41196 342904 41202 342916
rect 62114 342904 62120 342916
rect 41196 342876 62120 342904
rect 41196 342864 41202 342876
rect 62114 342864 62120 342876
rect 62172 342864 62178 342916
rect 118602 342864 118608 342916
rect 118660 342904 118666 342916
rect 130102 342904 130108 342916
rect 118660 342876 130108 342904
rect 118660 342864 118666 342876
rect 130102 342864 130108 342876
rect 130160 342864 130166 342916
rect 61838 342252 61844 342304
rect 61896 342292 61902 342304
rect 66070 342292 66076 342304
rect 61896 342264 66076 342292
rect 61896 342252 61902 342264
rect 66070 342252 66076 342264
rect 66128 342292 66134 342304
rect 67634 342292 67640 342304
rect 66128 342264 67640 342292
rect 66128 342252 66134 342264
rect 67634 342252 67640 342264
rect 67692 342252 67698 342304
rect 118602 342184 118608 342236
rect 118660 342224 118666 342236
rect 150526 342224 150532 342236
rect 118660 342196 150532 342224
rect 118660 342184 118666 342196
rect 150526 342184 150532 342196
rect 150584 342224 150590 342236
rect 150986 342224 150992 342236
rect 150584 342196 150992 342224
rect 150584 342184 150590 342196
rect 150986 342184 150992 342196
rect 151044 342184 151050 342236
rect 66162 341572 66168 341624
rect 66220 341612 66226 341624
rect 68646 341612 68652 341624
rect 66220 341584 68652 341612
rect 66220 341572 66226 341584
rect 68646 341572 68652 341584
rect 68704 341572 68710 341624
rect 150986 341504 150992 341556
rect 151044 341544 151050 341556
rect 348418 341544 348424 341556
rect 151044 341516 348424 341544
rect 151044 341504 151050 341516
rect 348418 341504 348424 341516
rect 348476 341504 348482 341556
rect 64138 340932 64144 340944
rect 63236 340904 64144 340932
rect 33042 340756 33048 340808
rect 33100 340796 33106 340808
rect 63236 340796 63264 340904
rect 64138 340892 64144 340904
rect 64196 340932 64202 340944
rect 67634 340932 67640 340944
rect 64196 340904 67640 340932
rect 64196 340892 64202 340904
rect 67634 340892 67640 340904
rect 67692 340892 67698 340944
rect 118050 340892 118056 340944
rect 118108 340932 118114 340944
rect 142246 340932 142252 340944
rect 118108 340904 142252 340932
rect 118108 340892 118114 340904
rect 142246 340892 142252 340904
rect 142304 340892 142310 340944
rect 63310 340824 63316 340876
rect 63368 340864 63374 340876
rect 68646 340864 68652 340876
rect 63368 340836 68652 340864
rect 63368 340824 63374 340836
rect 68646 340824 68652 340836
rect 68704 340824 68710 340876
rect 117958 340824 117964 340876
rect 118016 340864 118022 340876
rect 147766 340864 147772 340876
rect 118016 340836 147772 340864
rect 118016 340824 118022 340836
rect 147766 340824 147772 340836
rect 147824 340824 147830 340876
rect 33100 340768 63264 340796
rect 33100 340756 33106 340768
rect 118602 340756 118608 340808
rect 118660 340796 118666 340808
rect 135438 340796 135444 340808
rect 118660 340768 135444 340796
rect 118660 340756 118666 340768
rect 135438 340756 135444 340768
rect 135496 340796 135502 340808
rect 138014 340796 138020 340808
rect 135496 340768 138020 340796
rect 135496 340756 135502 340768
rect 138014 340756 138020 340768
rect 138072 340756 138078 340808
rect 147766 340144 147772 340196
rect 147824 340184 147830 340196
rect 338758 340184 338764 340196
rect 147824 340156 338764 340184
rect 147824 340144 147830 340156
rect 338758 340144 338764 340156
rect 338816 340144 338822 340196
rect 69014 340008 69020 340060
rect 69072 340048 69078 340060
rect 69750 340048 69756 340060
rect 69072 340020 69756 340048
rect 69072 340008 69078 340020
rect 69750 340008 69756 340020
rect 69808 340008 69814 340060
rect 71774 339872 71780 339924
rect 71832 339912 71838 339924
rect 72418 339912 72424 339924
rect 71832 339884 72424 339912
rect 71832 339872 71838 339884
rect 72418 339872 72424 339884
rect 72476 339872 72482 339924
rect 43898 339464 43904 339516
rect 43956 339504 43962 339516
rect 78398 339504 78404 339516
rect 43956 339476 78404 339504
rect 43956 339464 43962 339476
rect 78398 339464 78404 339476
rect 78456 339464 78462 339516
rect 97718 339464 97724 339516
rect 97776 339504 97782 339516
rect 129918 339504 129924 339516
rect 97776 339476 129924 339504
rect 97776 339464 97782 339476
rect 129918 339464 129924 339476
rect 129976 339464 129982 339516
rect 42518 339396 42524 339448
rect 42576 339436 42582 339448
rect 75178 339436 75184 339448
rect 42576 339408 75184 339436
rect 42576 339396 42582 339408
rect 75178 339396 75184 339408
rect 75236 339436 75242 339448
rect 75822 339436 75828 339448
rect 75236 339408 75828 339436
rect 75236 339396 75242 339408
rect 75822 339396 75828 339408
rect 75880 339396 75886 339448
rect 87414 339396 87420 339448
rect 87472 339436 87478 339448
rect 87690 339436 87696 339448
rect 87472 339408 87696 339436
rect 87472 339396 87478 339408
rect 87690 339396 87696 339408
rect 87748 339436 87754 339448
rect 121454 339436 121460 339448
rect 87748 339408 121460 339436
rect 87748 339396 87754 339408
rect 121454 339396 121460 339408
rect 121512 339396 121518 339448
rect 46750 339328 46756 339380
rect 46808 339368 46814 339380
rect 50706 339368 50712 339380
rect 46808 339340 50712 339368
rect 46808 339328 46814 339340
rect 50706 339328 50712 339340
rect 50764 339328 50770 339380
rect 99650 339328 99656 339380
rect 99708 339368 99714 339380
rect 100662 339368 100668 339380
rect 99708 339340 100668 339368
rect 99708 339328 99714 339340
rect 100662 339328 100668 339340
rect 100720 339368 100726 339380
rect 130010 339368 130016 339380
rect 100720 339340 130016 339368
rect 100720 339328 100726 339340
rect 130010 339328 130016 339340
rect 130068 339328 130074 339380
rect 67358 338852 67364 338904
rect 67416 338892 67422 338904
rect 77938 338892 77944 338904
rect 67416 338864 77944 338892
rect 67416 338852 67422 338864
rect 77938 338852 77944 338864
rect 77996 338852 78002 338904
rect 78398 338784 78404 338836
rect 78456 338824 78462 338836
rect 93118 338824 93124 338836
rect 78456 338796 93124 338824
rect 78456 338784 78462 338796
rect 93118 338784 93124 338796
rect 93176 338784 93182 338836
rect 64782 338716 64788 338768
rect 64840 338756 64846 338768
rect 87598 338756 87604 338768
rect 64840 338728 87604 338756
rect 64840 338716 64846 338728
rect 87598 338716 87604 338728
rect 87656 338716 87662 338768
rect 50706 338104 50712 338156
rect 50764 338144 50770 338156
rect 50764 338116 80100 338144
rect 50764 338104 50770 338116
rect 43990 338036 43996 338088
rect 44048 338076 44054 338088
rect 79042 338076 79048 338088
rect 44048 338048 79048 338076
rect 44048 338036 44054 338048
rect 79042 338036 79048 338048
rect 79100 338036 79106 338088
rect 80072 338076 80100 338116
rect 82262 338076 82268 338088
rect 80072 338048 82268 338076
rect 82262 338036 82268 338048
rect 82320 338036 82326 338088
rect 106182 338036 106188 338088
rect 106240 338076 106246 338088
rect 131114 338076 131120 338088
rect 106240 338048 131120 338076
rect 106240 338036 106246 338048
rect 131114 338036 131120 338048
rect 131172 338036 131178 338088
rect 57882 337968 57888 338020
rect 57940 338008 57946 338020
rect 84194 338008 84200 338020
rect 57940 337980 84200 338008
rect 57940 337968 57946 337980
rect 84194 337968 84200 337980
rect 84252 337968 84258 338020
rect 100294 337968 100300 338020
rect 100352 338008 100358 338020
rect 123018 338008 123024 338020
rect 100352 337980 123024 338008
rect 100352 337968 100358 337980
rect 123018 337968 123024 337980
rect 123076 337968 123082 338020
rect 56410 337900 56416 337952
rect 56468 337940 56474 337952
rect 76466 337940 76472 337952
rect 56468 337912 76472 337940
rect 56468 337900 56474 337912
rect 76466 337900 76472 337912
rect 76524 337900 76530 337952
rect 113818 337900 113824 337952
rect 113876 337940 113882 337952
rect 127066 337940 127072 337952
rect 113876 337912 127072 337940
rect 113876 337900 113882 337912
rect 127066 337900 127072 337912
rect 127124 337900 127130 337952
rect 55858 337832 55864 337884
rect 55916 337872 55922 337884
rect 74534 337872 74540 337884
rect 55916 337844 74540 337872
rect 55916 337832 55922 337844
rect 74534 337832 74540 337844
rect 74592 337872 74598 337884
rect 75270 337872 75276 337884
rect 74592 337844 75276 337872
rect 74592 337832 74598 337844
rect 75270 337832 75276 337844
rect 75328 337832 75334 337884
rect 103514 337560 103520 337612
rect 103572 337600 103578 337612
rect 114462 337600 114468 337612
rect 103572 337572 114468 337600
rect 103572 337560 103578 337572
rect 114462 337560 114468 337572
rect 114520 337560 114526 337612
rect 84838 337532 84844 337544
rect 64846 337504 84844 337532
rect 50890 337356 50896 337408
rect 50948 337396 50954 337408
rect 60550 337396 60556 337408
rect 50948 337368 60556 337396
rect 50948 337356 50954 337368
rect 60550 337356 60556 337368
rect 60608 337396 60614 337408
rect 64846 337396 64874 337504
rect 84838 337492 84844 337504
rect 84896 337492 84902 337544
rect 93946 337492 93952 337544
rect 94004 337532 94010 337544
rect 123110 337532 123116 337544
rect 94004 337504 123116 337532
rect 94004 337492 94010 337504
rect 123110 337492 123116 337504
rect 123168 337492 123174 337544
rect 79042 337424 79048 337476
rect 79100 337464 79106 337476
rect 220078 337464 220084 337476
rect 79100 337436 220084 337464
rect 79100 337424 79106 337436
rect 220078 337424 220084 337436
rect 220136 337424 220142 337476
rect 60608 337368 64874 337396
rect 60608 337356 60614 337368
rect 68554 337356 68560 337408
rect 68612 337396 68618 337408
rect 322198 337396 322204 337408
rect 68612 337368 322204 337396
rect 68612 337356 68618 337368
rect 322198 337356 322204 337368
rect 322256 337356 322262 337408
rect 59078 336676 59084 336728
rect 59136 336716 59142 336728
rect 92474 336716 92480 336728
rect 59136 336688 92480 336716
rect 59136 336676 59142 336688
rect 92474 336676 92480 336688
rect 92532 336676 92538 336728
rect 108022 336676 108028 336728
rect 108080 336716 108086 336728
rect 139578 336716 139584 336728
rect 108080 336688 139584 336716
rect 108080 336676 108086 336688
rect 139578 336676 139584 336688
rect 139636 336676 139642 336728
rect 39666 336608 39672 336660
rect 39724 336648 39730 336660
rect 71958 336648 71964 336660
rect 39724 336620 71964 336648
rect 39724 336608 39730 336620
rect 71958 336608 71964 336620
rect 72016 336648 72022 336660
rect 72510 336648 72516 336660
rect 72016 336620 72516 336648
rect 72016 336608 72022 336620
rect 72510 336608 72516 336620
rect 72568 336608 72574 336660
rect 115106 336608 115112 336660
rect 115164 336648 115170 336660
rect 115290 336648 115296 336660
rect 115164 336620 115296 336648
rect 115164 336608 115170 336620
rect 115290 336608 115296 336620
rect 115348 336608 115354 336660
rect 119430 336608 119436 336660
rect 119488 336648 119494 336660
rect 133966 336648 133972 336660
rect 119488 336620 133972 336648
rect 119488 336608 119494 336620
rect 133966 336608 133972 336620
rect 134024 336648 134030 336660
rect 135162 336648 135168 336660
rect 134024 336620 135168 336648
rect 134024 336608 134030 336620
rect 135162 336608 135168 336620
rect 135220 336608 135226 336660
rect 55030 336540 55036 336592
rect 55088 336580 55094 336592
rect 83458 336580 83464 336592
rect 55088 336552 83464 336580
rect 55088 336540 55094 336552
rect 83458 336540 83464 336552
rect 83516 336540 83522 336592
rect 115308 336580 115336 336608
rect 122834 336580 122840 336592
rect 115308 336552 122840 336580
rect 122834 336540 122840 336552
rect 122892 336540 122898 336592
rect 123478 336540 123484 336592
rect 123536 336580 123542 336592
rect 124214 336580 124220 336592
rect 123536 336552 124220 336580
rect 123536 336540 123542 336552
rect 124214 336540 124220 336552
rect 124272 336540 124278 336592
rect 53558 336472 53564 336524
rect 53616 336512 53622 336524
rect 79318 336512 79324 336524
rect 53616 336484 79324 336512
rect 53616 336472 53622 336484
rect 79318 336472 79324 336484
rect 79376 336472 79382 336524
rect 47946 336404 47952 336456
rect 48004 336444 48010 336456
rect 73338 336444 73344 336456
rect 48004 336416 73344 336444
rect 48004 336404 48010 336416
rect 73338 336404 73344 336416
rect 73396 336404 73402 336456
rect 92474 335996 92480 336048
rect 92532 336036 92538 336048
rect 93210 336036 93216 336048
rect 92532 336008 93216 336036
rect 92532 335996 92538 336008
rect 93210 335996 93216 336008
rect 93268 336036 93274 336048
rect 104158 336036 104164 336048
rect 93268 336008 104164 336036
rect 93268 335996 93274 336008
rect 104158 335996 104164 336008
rect 104216 335996 104222 336048
rect 114462 335996 114468 336048
rect 114520 336036 114526 336048
rect 123478 336036 123484 336048
rect 114520 336008 123484 336036
rect 114520 335996 114526 336008
rect 123478 335996 123484 336008
rect 123536 335996 123542 336048
rect 135162 335996 135168 336048
rect 135220 336036 135226 336048
rect 269758 336036 269764 336048
rect 135220 336008 269764 336036
rect 135220 335996 135226 336008
rect 269758 335996 269764 336008
rect 269816 335996 269822 336048
rect 46566 335248 46572 335300
rect 46624 335288 46630 335300
rect 81618 335288 81624 335300
rect 46624 335260 81624 335288
rect 46624 335248 46630 335260
rect 81618 335248 81624 335260
rect 81676 335248 81682 335300
rect 115198 335248 115204 335300
rect 115256 335288 115262 335300
rect 149146 335288 149152 335300
rect 115256 335260 149152 335288
rect 115256 335248 115262 335260
rect 149146 335248 149152 335260
rect 149204 335248 149210 335300
rect 50798 335180 50804 335232
rect 50856 335220 50862 335232
rect 86770 335220 86776 335232
rect 50856 335192 86776 335220
rect 50856 335180 50862 335192
rect 86770 335180 86776 335192
rect 86828 335180 86834 335232
rect 109954 335180 109960 335232
rect 110012 335220 110018 335232
rect 128814 335220 128820 335232
rect 110012 335192 128820 335220
rect 110012 335180 110018 335192
rect 128814 335180 128820 335192
rect 128872 335220 128878 335232
rect 133966 335220 133972 335232
rect 128872 335192 133972 335220
rect 128872 335180 128878 335192
rect 133966 335180 133972 335192
rect 134024 335180 134030 335232
rect 60642 335112 60648 335164
rect 60700 335152 60706 335164
rect 94498 335152 94504 335164
rect 60700 335124 94504 335152
rect 60700 335112 60706 335124
rect 94498 335112 94504 335124
rect 94556 335112 94562 335164
rect 102870 335112 102876 335164
rect 102928 335152 102934 335164
rect 103422 335152 103428 335164
rect 102928 335124 103428 335152
rect 102928 335112 102934 335124
rect 103422 335112 103428 335124
rect 103480 335152 103486 335164
rect 120074 335152 120080 335164
rect 103480 335124 120080 335152
rect 103480 335112 103486 335124
rect 120074 335112 120080 335124
rect 120132 335112 120138 335164
rect 58986 335044 58992 335096
rect 59044 335084 59050 335096
rect 80974 335084 80980 335096
rect 59044 335056 80980 335084
rect 59044 335044 59050 335056
rect 80974 335044 80980 335056
rect 81032 335044 81038 335096
rect 86310 334636 86316 334688
rect 86368 334676 86374 334688
rect 86770 334676 86776 334688
rect 86368 334648 86776 334676
rect 86368 334636 86374 334648
rect 86770 334636 86776 334648
rect 86828 334636 86834 334688
rect 100018 334636 100024 334688
rect 100076 334676 100082 334688
rect 124398 334676 124404 334688
rect 100076 334648 124404 334676
rect 100076 334636 100082 334648
rect 124398 334636 124404 334648
rect 124456 334636 124462 334688
rect 56502 334568 56508 334620
rect 56560 334608 56566 334620
rect 119430 334608 119436 334620
rect 56560 334580 119436 334608
rect 56560 334568 56566 334580
rect 119430 334568 119436 334580
rect 119488 334568 119494 334620
rect 81618 333956 81624 334008
rect 81676 333996 81682 334008
rect 82078 333996 82084 334008
rect 81676 333968 82084 333996
rect 81676 333956 81682 333968
rect 82078 333956 82084 333968
rect 82136 333956 82142 334008
rect 49510 333888 49516 333940
rect 49568 333928 49574 333940
rect 86218 333928 86224 333940
rect 49568 333900 86224 333928
rect 49568 333888 49574 333900
rect 86218 333888 86224 333900
rect 86276 333888 86282 333940
rect 97074 333888 97080 333940
rect 97132 333928 97138 333940
rect 127250 333928 127256 333940
rect 97132 333900 127256 333928
rect 97132 333888 97138 333900
rect 127250 333888 127256 333900
rect 127308 333888 127314 333940
rect 57698 333276 57704 333328
rect 57756 333316 57762 333328
rect 87690 333316 87696 333328
rect 57756 333288 87696 333316
rect 57756 333276 57762 333288
rect 87690 333276 87696 333288
rect 87748 333276 87754 333328
rect 95142 333276 95148 333328
rect 95200 333316 95206 333328
rect 113818 333316 113824 333328
rect 95200 333288 113824 333316
rect 95200 333276 95206 333288
rect 113818 333276 113824 333288
rect 113876 333276 113882 333328
rect 68738 333208 68744 333260
rect 68796 333248 68802 333260
rect 309778 333248 309784 333260
rect 68796 333220 309784 333248
rect 68796 333208 68802 333220
rect 309778 333208 309784 333220
rect 309836 333208 309842 333260
rect 97074 332732 97080 332784
rect 97132 332772 97138 332784
rect 97902 332772 97908 332784
rect 97132 332744 97908 332772
rect 97132 332732 97138 332744
rect 97902 332732 97908 332744
rect 97960 332732 97966 332784
rect 108298 332528 108304 332580
rect 108356 332568 108362 332580
rect 142154 332568 142160 332580
rect 108356 332540 142160 332568
rect 108356 332528 108362 332540
rect 142154 332528 142160 332540
rect 142212 332568 142218 332580
rect 143442 332568 143448 332580
rect 142212 332540 143448 332568
rect 142212 332528 142218 332540
rect 143442 332528 143448 332540
rect 143500 332528 143506 332580
rect 61930 331916 61936 331968
rect 61988 331956 61994 331968
rect 98638 331956 98644 331968
rect 61988 331928 98644 331956
rect 61988 331916 61994 331928
rect 98638 331916 98644 331928
rect 98696 331916 98702 331968
rect 64138 331848 64144 331900
rect 64196 331888 64202 331900
rect 124214 331888 124220 331900
rect 64196 331860 124220 331888
rect 64196 331848 64202 331860
rect 124214 331848 124220 331860
rect 124272 331848 124278 331900
rect 143442 331848 143448 331900
rect 143500 331888 143506 331900
rect 409874 331888 409880 331900
rect 143500 331860 409880 331888
rect 143500 331848 143506 331860
rect 409874 331848 409880 331860
rect 409932 331848 409938 331900
rect 59262 331168 59268 331220
rect 59320 331208 59326 331220
rect 88978 331208 88984 331220
rect 59320 331180 88984 331208
rect 59320 331168 59326 331180
rect 88978 331168 88984 331180
rect 89036 331168 89042 331220
rect 105446 331168 105452 331220
rect 105504 331208 105510 331220
rect 136818 331208 136824 331220
rect 105504 331180 136824 331208
rect 105504 331168 105510 331180
rect 136818 331168 136824 331180
rect 136876 331208 136882 331220
rect 137094 331208 137100 331220
rect 136876 331180 137100 331208
rect 136876 331168 136882 331180
rect 137094 331168 137100 331180
rect 137152 331168 137158 331220
rect 60458 330488 60464 330540
rect 60516 330528 60522 330540
rect 115198 330528 115204 330540
rect 60516 330500 115204 330528
rect 60516 330488 60522 330500
rect 115198 330488 115204 330500
rect 115256 330488 115262 330540
rect 137094 330488 137100 330540
rect 137152 330528 137158 330540
rect 425698 330528 425704 330540
rect 137152 330500 425704 330528
rect 137152 330488 137158 330500
rect 425698 330488 425704 330500
rect 425756 330488 425762 330540
rect 88702 329740 88708 329792
rect 88760 329780 88766 329792
rect 122006 329780 122012 329792
rect 88760 329752 122012 329780
rect 88760 329740 88766 329752
rect 122006 329740 122012 329752
rect 122064 329740 122070 329792
rect 92566 329672 92572 329724
rect 92624 329712 92630 329724
rect 125962 329712 125968 329724
rect 92624 329684 125968 329712
rect 92624 329672 92630 329684
rect 125962 329672 125968 329684
rect 126020 329712 126026 329724
rect 126882 329712 126888 329724
rect 126020 329684 126888 329712
rect 126020 329672 126026 329684
rect 126882 329672 126888 329684
rect 126940 329672 126946 329724
rect 69198 329128 69204 329180
rect 69256 329168 69262 329180
rect 121454 329168 121460 329180
rect 69256 329140 121460 329168
rect 69256 329128 69262 329140
rect 121454 329128 121460 329140
rect 121512 329128 121518 329180
rect 48130 329060 48136 329112
rect 48188 329100 48194 329112
rect 108022 329100 108028 329112
rect 48188 329072 108028 329100
rect 48188 329060 48194 329072
rect 108022 329060 108028 329072
rect 108080 329060 108086 329112
rect 126882 329060 126888 329112
rect 126940 329100 126946 329112
rect 295978 329100 295984 329112
rect 126940 329072 295984 329100
rect 126940 329060 126946 329072
rect 295978 329060 295984 329072
rect 296036 329060 296042 329112
rect 4798 328448 4804 328500
rect 4856 328488 4862 328500
rect 48130 328488 48136 328500
rect 4856 328460 48136 328488
rect 4856 328448 4862 328460
rect 48130 328448 48136 328460
rect 48188 328448 48194 328500
rect 122006 328448 122012 328500
rect 122064 328488 122070 328500
rect 216030 328488 216036 328500
rect 122064 328460 216036 328488
rect 122064 328448 122070 328460
rect 216030 328448 216036 328460
rect 216088 328448 216094 328500
rect 106090 327904 106096 327956
rect 106148 327944 106154 327956
rect 116026 327944 116032 327956
rect 106148 327916 116032 327944
rect 106148 327904 106154 327916
rect 116026 327904 116032 327916
rect 116084 327904 116090 327956
rect 91922 327836 91928 327888
rect 91980 327876 91986 327888
rect 125594 327876 125600 327888
rect 91980 327848 125600 327876
rect 91980 327836 91986 327848
rect 125594 327836 125600 327848
rect 125652 327836 125658 327888
rect 66070 327768 66076 327820
rect 66128 327808 66134 327820
rect 269850 327808 269856 327820
rect 66128 327780 269856 327808
rect 66128 327768 66134 327780
rect 269850 327768 269856 327780
rect 269908 327768 269914 327820
rect 78030 327700 78036 327752
rect 78088 327740 78094 327752
rect 358078 327740 358084 327752
rect 78088 327712 358084 327740
rect 78088 327700 78094 327712
rect 358078 327700 358084 327712
rect 358136 327700 358142 327752
rect 112530 327020 112536 327072
rect 112588 327060 112594 327072
rect 146386 327060 146392 327072
rect 112588 327032 146392 327060
rect 112588 327020 112594 327032
rect 146386 327020 146392 327032
rect 146444 327060 146450 327072
rect 146754 327060 146760 327072
rect 146444 327032 146760 327060
rect 146444 327020 146450 327032
rect 146754 327020 146760 327032
rect 146812 327020 146818 327072
rect 76558 326476 76564 326528
rect 76616 326516 76622 326528
rect 122190 326516 122196 326528
rect 76616 326488 122196 326516
rect 76616 326476 76622 326488
rect 122190 326476 122196 326488
rect 122248 326476 122254 326528
rect 214558 326448 214564 326460
rect 122806 326420 214564 326448
rect 71038 326340 71044 326392
rect 71096 326380 71102 326392
rect 122098 326380 122104 326392
rect 71096 326352 122104 326380
rect 71096 326340 71102 326352
rect 122098 326340 122104 326352
rect 122156 326380 122162 326392
rect 122806 326380 122834 326420
rect 214558 326408 214564 326420
rect 214616 326408 214622 326460
rect 122156 326352 122834 326380
rect 122156 326340 122162 326352
rect 146754 326340 146760 326392
rect 146812 326380 146818 326392
rect 254578 326380 254584 326392
rect 146812 326352 254584 326380
rect 146812 326340 146818 326352
rect 254578 326340 254584 326352
rect 254636 326340 254642 326392
rect 63218 325048 63224 325100
rect 63276 325088 63282 325100
rect 177298 325088 177304 325100
rect 63276 325060 177304 325088
rect 63276 325048 63282 325060
rect 177298 325048 177304 325060
rect 177356 325048 177362 325100
rect 82078 324980 82084 325032
rect 82136 325020 82142 325032
rect 268378 325020 268384 325032
rect 82136 324992 268384 325020
rect 82136 324980 82142 324992
rect 268378 324980 268384 324992
rect 268436 324980 268442 325032
rect 72510 324912 72516 324964
rect 72568 324952 72574 324964
rect 300118 324952 300124 324964
rect 72568 324924 300124 324952
rect 72568 324912 72574 324924
rect 300118 324912 300124 324924
rect 300176 324912 300182 324964
rect 95786 324232 95792 324284
rect 95844 324272 95850 324284
rect 128630 324272 128636 324284
rect 95844 324244 128636 324272
rect 95844 324232 95850 324244
rect 128630 324232 128636 324244
rect 128688 324232 128694 324284
rect 73154 323552 73160 323604
rect 73212 323592 73218 323604
rect 115934 323592 115940 323604
rect 73212 323564 115940 323592
rect 73212 323552 73218 323564
rect 115934 323552 115940 323564
rect 115992 323552 115998 323604
rect 128630 323552 128636 323604
rect 128688 323592 128694 323604
rect 395338 323592 395344 323604
rect 128688 323564 395344 323592
rect 128688 323552 128694 323564
rect 395338 323552 395344 323564
rect 395396 323552 395402 323604
rect 110598 322872 110604 322924
rect 110656 322912 110662 322924
rect 140958 322912 140964 322924
rect 110656 322884 140964 322912
rect 110656 322872 110662 322884
rect 140958 322872 140964 322884
rect 141016 322872 141022 322924
rect 140958 322260 140964 322312
rect 141016 322300 141022 322312
rect 302878 322300 302884 322312
rect 141016 322272 302884 322300
rect 141016 322260 141022 322272
rect 302878 322260 302884 322272
rect 302936 322260 302942 322312
rect 86310 322192 86316 322244
rect 86368 322232 86374 322244
rect 399478 322232 399484 322244
rect 86368 322204 399484 322232
rect 86368 322192 86374 322204
rect 399478 322192 399484 322204
rect 399536 322192 399542 322244
rect 89990 321512 89996 321564
rect 90048 321552 90054 321564
rect 124306 321552 124312 321564
rect 90048 321524 124312 321552
rect 90048 321512 90054 321524
rect 124306 321512 124312 321524
rect 124364 321552 124370 321564
rect 125502 321552 125508 321564
rect 124364 321524 125508 321552
rect 124364 321512 124370 321524
rect 125502 321512 125508 321524
rect 125560 321512 125566 321564
rect 67542 320900 67548 320952
rect 67600 320940 67606 320952
rect 116118 320940 116124 320952
rect 67600 320912 116124 320940
rect 67600 320900 67606 320912
rect 116118 320900 116124 320912
rect 116176 320900 116182 320952
rect 125502 320900 125508 320952
rect 125560 320940 125566 320952
rect 266998 320940 267004 320952
rect 125560 320912 267004 320940
rect 125560 320900 125566 320912
rect 266998 320900 267004 320912
rect 267056 320900 267062 320952
rect 68830 320832 68836 320884
rect 68888 320872 68894 320884
rect 336090 320872 336096 320884
rect 68888 320844 336096 320872
rect 68888 320832 68894 320844
rect 336090 320832 336096 320844
rect 336148 320832 336154 320884
rect 100938 320084 100944 320136
rect 100996 320124 101002 320136
rect 132770 320124 132776 320136
rect 100996 320096 132776 320124
rect 100996 320084 101002 320096
rect 132770 320084 132776 320096
rect 132828 320124 132834 320136
rect 133782 320124 133788 320136
rect 132828 320096 133788 320124
rect 132828 320084 132834 320096
rect 133782 320084 133788 320096
rect 133840 320084 133846 320136
rect 93762 319540 93768 319592
rect 93820 319580 93826 319592
rect 115290 319580 115296 319592
rect 93820 319552 115296 319580
rect 93820 319540 93826 319552
rect 115290 319540 115296 319552
rect 115348 319540 115354 319592
rect 3234 319472 3240 319524
rect 3292 319512 3298 319524
rect 18598 319512 18604 319524
rect 3292 319484 18604 319512
rect 3292 319472 3298 319484
rect 18598 319472 18604 319484
rect 18656 319512 18662 319524
rect 101398 319512 101404 319524
rect 18656 319484 101404 319512
rect 18656 319472 18662 319484
rect 101398 319472 101404 319484
rect 101456 319472 101462 319524
rect 133782 319472 133788 319524
rect 133840 319512 133846 319524
rect 216122 319512 216128 319524
rect 133840 319484 216128 319512
rect 133840 319472 133846 319484
rect 216122 319472 216128 319484
rect 216180 319472 216186 319524
rect 68922 319404 68928 319456
rect 68980 319444 68986 319456
rect 343634 319444 343640 319456
rect 68980 319416 343640 319444
rect 68980 319404 68986 319416
rect 343634 319404 343640 319416
rect 343692 319404 343698 319456
rect 91278 318724 91284 318776
rect 91336 318764 91342 318776
rect 118694 318764 118700 318776
rect 91336 318736 118700 318764
rect 91336 318724 91342 318736
rect 118694 318724 118700 318736
rect 118752 318724 118758 318776
rect 111242 318656 111248 318708
rect 111300 318696 111306 318708
rect 131298 318696 131304 318708
rect 111300 318668 131304 318696
rect 111300 318656 111306 318668
rect 131298 318656 131304 318668
rect 131356 318696 131362 318708
rect 131666 318696 131672 318708
rect 131356 318668 131672 318696
rect 131356 318656 131362 318668
rect 131666 318656 131672 318668
rect 131724 318656 131730 318708
rect 131666 318112 131672 318164
rect 131724 318152 131730 318164
rect 265618 318152 265624 318164
rect 131724 318124 265624 318152
rect 131724 318112 131730 318124
rect 265618 318112 265624 318124
rect 265676 318112 265682 318164
rect 75270 318044 75276 318096
rect 75328 318084 75334 318096
rect 115290 318084 115296 318096
rect 75328 318056 115296 318084
rect 75328 318044 75334 318056
rect 115290 318044 115296 318056
rect 115348 318044 115354 318096
rect 118694 318044 118700 318096
rect 118752 318084 118758 318096
rect 267090 318084 267096 318096
rect 118752 318056 267096 318084
rect 118752 318044 118758 318056
rect 267090 318044 267096 318056
rect 267148 318044 267154 318096
rect 102226 317364 102232 317416
rect 102284 317404 102290 317416
rect 132678 317404 132684 317416
rect 102284 317376 132684 317404
rect 102284 317364 102290 317376
rect 132678 317364 132684 317376
rect 132736 317404 132742 317416
rect 133782 317404 133788 317416
rect 132736 317376 133788 317404
rect 132736 317364 132742 317376
rect 133782 317364 133788 317376
rect 133840 317364 133846 317416
rect 72510 316684 72516 316736
rect 72568 316724 72574 316736
rect 108298 316724 108304 316736
rect 72568 316696 108304 316724
rect 72568 316684 72574 316696
rect 108298 316684 108304 316696
rect 108356 316684 108362 316736
rect 133782 316684 133788 316736
rect 133840 316724 133846 316736
rect 345014 316724 345020 316736
rect 133840 316696 345020 316724
rect 133840 316684 133846 316696
rect 345014 316684 345020 316696
rect 345072 316684 345078 316736
rect 84286 316072 84292 316124
rect 84344 316112 84350 316124
rect 113174 316112 113180 316124
rect 84344 316084 113180 316112
rect 84344 316072 84350 316084
rect 113174 316072 113180 316084
rect 113232 316072 113238 316124
rect 69198 316004 69204 316056
rect 69256 316044 69262 316056
rect 104250 316044 104256 316056
rect 69256 316016 104256 316044
rect 69256 316004 69262 316016
rect 104250 316004 104256 316016
rect 104308 316004 104314 316056
rect 72418 315256 72424 315308
rect 72476 315296 72482 315308
rect 159358 315296 159364 315308
rect 72476 315268 159364 315296
rect 72476 315256 72482 315268
rect 159358 315256 159364 315268
rect 159416 315256 159422 315308
rect 91094 314644 91100 314696
rect 91152 314684 91158 314696
rect 231118 314684 231124 314696
rect 91152 314656 231124 314684
rect 91152 314644 91158 314656
rect 231118 314644 231124 314656
rect 231176 314644 231182 314696
rect 57606 313964 57612 314016
rect 57664 314004 57670 314016
rect 80054 314004 80060 314016
rect 57664 313976 80060 314004
rect 57664 313964 57670 313976
rect 80054 313964 80060 313976
rect 80112 314004 80118 314016
rect 91094 314004 91100 314016
rect 80112 313976 91100 314004
rect 80112 313964 80118 313976
rect 91094 313964 91100 313976
rect 91152 313964 91158 314016
rect 93118 313964 93124 314016
rect 93176 314004 93182 314016
rect 151078 314004 151084 314016
rect 93176 313976 151084 314004
rect 93176 313964 93182 313976
rect 151078 313964 151084 313976
rect 151136 313964 151142 314016
rect 67450 313896 67456 313948
rect 67508 313936 67514 313948
rect 125870 313936 125876 313948
rect 67508 313908 125876 313936
rect 67508 313896 67514 313908
rect 125870 313896 125876 313908
rect 125928 313896 125934 313948
rect 81434 313284 81440 313336
rect 81492 313324 81498 313336
rect 226978 313324 226984 313336
rect 81492 313296 226984 313324
rect 81492 313284 81498 313296
rect 226978 313284 226984 313296
rect 227036 313284 227042 313336
rect 65518 311856 65524 311908
rect 65576 311896 65582 311908
rect 66162 311896 66168 311908
rect 65576 311868 66168 311896
rect 65576 311856 65582 311868
rect 66162 311856 66168 311868
rect 66220 311896 66226 311908
rect 264238 311896 264244 311908
rect 66220 311868 264244 311896
rect 66220 311856 66226 311868
rect 264238 311856 264244 311868
rect 264296 311856 264302 311908
rect 453298 311856 453304 311908
rect 453356 311896 453362 311908
rect 579982 311896 579988 311908
rect 453356 311868 579988 311896
rect 453356 311856 453362 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 101398 311244 101404 311296
rect 101456 311284 101462 311296
rect 116578 311284 116584 311296
rect 101456 311256 116584 311284
rect 101456 311244 101462 311256
rect 116578 311244 116584 311256
rect 116636 311244 116642 311296
rect 87598 311176 87604 311228
rect 87656 311216 87662 311228
rect 162118 311216 162124 311228
rect 87656 311188 162124 311216
rect 87656 311176 87662 311188
rect 162118 311176 162124 311188
rect 162176 311176 162182 311228
rect 115842 311108 115848 311160
rect 115900 311148 115906 311160
rect 135898 311148 135904 311160
rect 115900 311120 135904 311148
rect 115900 311108 115906 311120
rect 135898 311108 135904 311120
rect 135956 311148 135962 311160
rect 271138 311148 271144 311160
rect 135956 311120 271144 311148
rect 135956 311108 135962 311120
rect 271138 311108 271144 311120
rect 271196 311108 271202 311160
rect 84378 309884 84384 309936
rect 84436 309924 84442 309936
rect 115842 309924 115848 309936
rect 84436 309896 115848 309924
rect 84436 309884 84442 309896
rect 115842 309884 115848 309896
rect 115900 309884 115906 309936
rect 104894 309816 104900 309868
rect 104952 309856 104958 309868
rect 145006 309856 145012 309868
rect 104952 309828 145012 309856
rect 104952 309816 104958 309828
rect 145006 309816 145012 309828
rect 145064 309856 145070 309868
rect 445754 309856 445760 309868
rect 145064 309828 445760 309856
rect 145064 309816 145070 309828
rect 445754 309816 445760 309828
rect 445812 309816 445818 309868
rect 113174 309748 113180 309800
rect 113232 309788 113238 309800
rect 433334 309788 433340 309800
rect 113232 309760 433340 309788
rect 113232 309748 113238 309760
rect 433334 309748 433340 309760
rect 433392 309748 433398 309800
rect 75914 309136 75920 309188
rect 75972 309176 75978 309188
rect 155310 309176 155316 309188
rect 75972 309148 155316 309176
rect 75972 309136 75978 309148
rect 155310 309136 155316 309148
rect 155368 309136 155374 309188
rect 104250 309068 104256 309120
rect 104308 309108 104314 309120
rect 138198 309108 138204 309120
rect 104308 309080 138204 309108
rect 104308 309068 104314 309080
rect 138198 309068 138204 309080
rect 138256 309108 138262 309120
rect 138658 309108 138664 309120
rect 138256 309080 138664 309108
rect 138256 309068 138262 309080
rect 138658 309068 138664 309080
rect 138716 309068 138722 309120
rect 74442 308456 74448 308508
rect 74500 308496 74506 308508
rect 121546 308496 121552 308508
rect 74500 308468 121552 308496
rect 74500 308456 74506 308468
rect 121546 308456 121552 308468
rect 121604 308456 121610 308508
rect 138658 308456 138664 308508
rect 138716 308496 138722 308508
rect 262950 308496 262956 308508
rect 138716 308468 262956 308496
rect 138716 308456 138722 308468
rect 262950 308456 262956 308468
rect 263008 308456 263014 308508
rect 83458 308388 83464 308440
rect 83516 308428 83522 308440
rect 345658 308428 345664 308440
rect 83516 308400 345664 308428
rect 83516 308388 83522 308400
rect 345658 308388 345664 308400
rect 345716 308388 345722 308440
rect 88334 307776 88340 307828
rect 88392 307816 88398 307828
rect 153838 307816 153844 307828
rect 88392 307788 153844 307816
rect 88392 307776 88398 307788
rect 153838 307776 153844 307788
rect 153896 307776 153902 307828
rect 94222 307708 94228 307760
rect 94280 307748 94286 307760
rect 94590 307748 94596 307760
rect 94280 307720 94596 307748
rect 94280 307708 94286 307720
rect 94590 307708 94596 307720
rect 94648 307748 94654 307760
rect 128538 307748 128544 307760
rect 94648 307720 128544 307748
rect 94648 307708 94654 307720
rect 128538 307708 128544 307720
rect 128596 307748 128602 307760
rect 128722 307748 128728 307760
rect 128596 307720 128728 307748
rect 128596 307708 128602 307720
rect 128722 307708 128728 307720
rect 128780 307708 128786 307760
rect 128722 307164 128728 307216
rect 128780 307204 128786 307216
rect 155218 307204 155224 307216
rect 128780 307176 155224 307204
rect 128780 307164 128786 307176
rect 155218 307164 155224 307176
rect 155276 307164 155282 307216
rect 97902 307096 97908 307148
rect 97960 307136 97966 307148
rect 334618 307136 334624 307148
rect 97960 307108 334624 307136
rect 97960 307096 97966 307108
rect 334618 307096 334624 307108
rect 334676 307096 334682 307148
rect 106182 307028 106188 307080
rect 106240 307068 106246 307080
rect 113818 307068 113824 307080
rect 106240 307040 113824 307068
rect 106240 307028 106246 307040
rect 113818 307028 113824 307040
rect 113876 307028 113882 307080
rect 118694 307028 118700 307080
rect 118752 307068 118758 307080
rect 146570 307068 146576 307080
rect 118752 307040 146576 307068
rect 118752 307028 118758 307040
rect 146570 307028 146576 307040
rect 146628 307068 146634 307080
rect 403618 307068 403624 307080
rect 146628 307040 403624 307068
rect 146628 307028 146634 307040
rect 403618 307028 403624 307040
rect 403676 307028 403682 307080
rect 74534 306348 74540 306400
rect 74592 306388 74598 306400
rect 167638 306388 167644 306400
rect 74592 306360 167644 306388
rect 74592 306348 74598 306360
rect 167638 306348 167644 306360
rect 167696 306348 167702 306400
rect 98362 306280 98368 306332
rect 98420 306320 98426 306332
rect 125778 306320 125784 306332
rect 98420 306292 125784 306320
rect 98420 306280 98426 306292
rect 125778 306280 125784 306292
rect 125836 306280 125842 306332
rect 143626 306280 143632 306332
rect 143684 306320 143690 306332
rect 580258 306320 580264 306332
rect 143684 306292 580264 306320
rect 143684 306280 143690 306292
rect 580258 306280 580264 306292
rect 580316 306280 580322 306332
rect 3418 306212 3424 306264
rect 3476 306252 3482 306264
rect 7558 306252 7564 306264
rect 3476 306224 7564 306252
rect 3476 306212 3482 306224
rect 7558 306212 7564 306224
rect 7616 306212 7622 306264
rect 121270 305668 121276 305720
rect 121328 305708 121334 305720
rect 143626 305708 143632 305720
rect 121328 305680 143632 305708
rect 121328 305668 121334 305680
rect 143626 305668 143632 305680
rect 143684 305668 143690 305720
rect 97718 305600 97724 305652
rect 97776 305640 97782 305652
rect 341610 305640 341616 305652
rect 97776 305612 341616 305640
rect 97776 305600 97782 305612
rect 341610 305600 341616 305612
rect 341668 305600 341674 305652
rect 125778 305124 125784 305176
rect 125836 305164 125842 305176
rect 128538 305164 128544 305176
rect 125836 305136 128544 305164
rect 125836 305124 125842 305136
rect 128538 305124 128544 305136
rect 128596 305124 128602 305176
rect 85574 305056 85580 305108
rect 85632 305096 85638 305108
rect 214650 305096 214656 305108
rect 85632 305068 214656 305096
rect 85632 305056 85638 305068
rect 214650 305056 214656 305068
rect 214708 305056 214714 305108
rect 114554 304988 114560 305040
rect 114612 305028 114618 305040
rect 115290 305028 115296 305040
rect 114612 305000 115296 305028
rect 114612 304988 114618 305000
rect 115290 304988 115296 305000
rect 115348 305028 115354 305040
rect 245010 305028 245016 305040
rect 115348 305000 245016 305028
rect 115348 304988 115354 305000
rect 245010 304988 245016 305000
rect 245068 304988 245074 305040
rect 100662 304580 100668 304632
rect 100720 304620 100726 304632
rect 104250 304620 104256 304632
rect 100720 304592 104256 304620
rect 100720 304580 100726 304592
rect 104250 304580 104256 304592
rect 104308 304580 104314 304632
rect 57514 304240 57520 304292
rect 57572 304280 57578 304292
rect 126238 304280 126244 304292
rect 57572 304252 126244 304280
rect 57572 304240 57578 304252
rect 126238 304240 126244 304252
rect 126296 304240 126302 304292
rect 98638 303900 98644 303952
rect 98696 303940 98702 303952
rect 180058 303940 180064 303952
rect 98696 303912 180064 303940
rect 98696 303900 98702 303912
rect 180058 303900 180064 303912
rect 180116 303900 180122 303952
rect 92658 303832 92664 303884
rect 92716 303872 92722 303884
rect 210418 303872 210424 303884
rect 92716 303844 210424 303872
rect 92716 303832 92722 303844
rect 210418 303832 210424 303844
rect 210476 303832 210482 303884
rect 73246 303764 73252 303816
rect 73304 303804 73310 303816
rect 228450 303804 228456 303816
rect 73304 303776 228456 303804
rect 73304 303764 73310 303776
rect 228450 303764 228456 303776
rect 228508 303764 228514 303816
rect 95160 303708 103514 303736
rect 95160 303680 95188 303708
rect 94038 303628 94044 303680
rect 94096 303668 94102 303680
rect 95142 303668 95148 303680
rect 94096 303640 95148 303668
rect 94096 303628 94102 303640
rect 95142 303628 95148 303640
rect 95200 303628 95206 303680
rect 97994 303628 98000 303680
rect 98052 303668 98058 303680
rect 98638 303668 98644 303680
rect 98052 303640 98644 303668
rect 98052 303628 98058 303640
rect 98638 303628 98644 303640
rect 98696 303628 98702 303680
rect 103486 303668 103514 303708
rect 115934 303696 115940 303748
rect 115992 303736 115998 303748
rect 116578 303736 116584 303748
rect 115992 303708 116584 303736
rect 115992 303696 115998 303708
rect 116578 303696 116584 303708
rect 116636 303736 116642 303748
rect 326338 303736 326344 303748
rect 116636 303708 326344 303736
rect 116636 303696 116642 303708
rect 326338 303696 326344 303708
rect 326396 303696 326402 303748
rect 416774 303668 416780 303680
rect 103486 303640 416780 303668
rect 416774 303628 416780 303640
rect 416832 303628 416838 303680
rect 106826 303016 106832 303068
rect 106884 303056 106890 303068
rect 132586 303056 132592 303068
rect 106884 303028 132592 303056
rect 106884 303016 106890 303028
rect 132586 303016 132592 303028
rect 132644 303056 132650 303068
rect 173158 303056 173164 303068
rect 132644 303028 173164 303056
rect 132644 303016 132650 303028
rect 173158 303016 173164 303028
rect 173216 303016 173222 303068
rect 75270 302948 75276 303000
rect 75328 302988 75334 303000
rect 131206 302988 131212 303000
rect 75328 302960 131212 302988
rect 75328 302948 75334 302960
rect 131206 302948 131212 302960
rect 131264 302988 131270 303000
rect 353938 302988 353944 303000
rect 131264 302960 353944 302988
rect 131264 302948 131270 302960
rect 353938 302948 353944 302960
rect 353996 302948 354002 303000
rect 75178 302880 75184 302932
rect 75236 302920 75242 302932
rect 331950 302920 331956 302932
rect 75236 302892 331956 302920
rect 75236 302880 75242 302892
rect 331950 302880 331956 302892
rect 332008 302880 332014 302932
rect 87506 302268 87512 302320
rect 87564 302308 87570 302320
rect 240778 302308 240784 302320
rect 87564 302280 240784 302308
rect 87564 302268 87570 302280
rect 240778 302268 240784 302280
rect 240836 302268 240842 302320
rect 86310 302200 86316 302252
rect 86368 302240 86374 302252
rect 276658 302240 276664 302252
rect 86368 302212 276664 302240
rect 86368 302200 86374 302212
rect 276658 302200 276664 302212
rect 276716 302200 276722 302252
rect 104986 301316 104992 301368
rect 105044 301356 105050 301368
rect 106090 301356 106096 301368
rect 105044 301328 106096 301356
rect 105044 301316 105050 301328
rect 106090 301316 106096 301328
rect 106148 301316 106154 301368
rect 90266 301180 90272 301232
rect 90324 301220 90330 301232
rect 220170 301220 220176 301232
rect 90324 301192 220176 301220
rect 90324 301180 90330 301192
rect 220170 301180 220176 301192
rect 220228 301180 220234 301232
rect 81526 301112 81532 301164
rect 81584 301152 81590 301164
rect 251818 301152 251824 301164
rect 81584 301124 251824 301152
rect 81584 301112 81590 301124
rect 251818 301112 251824 301124
rect 251876 301112 251882 301164
rect 98638 301044 98644 301096
rect 98696 301084 98702 301096
rect 283006 301084 283012 301096
rect 98696 301056 283012 301084
rect 98696 301044 98702 301056
rect 283006 301044 283012 301056
rect 283064 301044 283070 301096
rect 109034 300976 109040 301028
rect 109092 301016 109098 301028
rect 298094 301016 298100 301028
rect 109092 300988 298100 301016
rect 109092 300976 109098 300988
rect 298094 300976 298100 300988
rect 298152 300976 298158 301028
rect 71774 300908 71780 300960
rect 71832 300948 71838 300960
rect 306374 300948 306380 300960
rect 71832 300920 306380 300948
rect 71832 300908 71838 300920
rect 306374 300908 306380 300920
rect 306432 300908 306438 300960
rect 106090 300840 106096 300892
rect 106148 300880 106154 300892
rect 450538 300880 450544 300892
rect 106148 300852 450544 300880
rect 106148 300840 106154 300852
rect 450538 300840 450544 300852
rect 450596 300840 450602 300892
rect 86218 300160 86224 300212
rect 86276 300200 86282 300212
rect 132586 300200 132592 300212
rect 86276 300172 132592 300200
rect 86276 300160 86282 300172
rect 132586 300160 132592 300172
rect 132644 300160 132650 300212
rect 69014 300092 69020 300144
rect 69072 300132 69078 300144
rect 342254 300132 342260 300144
rect 69072 300104 342260 300132
rect 69072 300092 69078 300104
rect 342254 300092 342260 300104
rect 342312 300092 342318 300144
rect 112438 299684 112444 299736
rect 112496 299724 112502 299736
rect 227070 299724 227076 299736
rect 112496 299696 227076 299724
rect 112496 299684 112502 299696
rect 227070 299684 227076 299696
rect 227128 299684 227134 299736
rect 100846 299616 100852 299668
rect 100904 299656 100910 299668
rect 256694 299656 256700 299668
rect 100904 299628 256700 299656
rect 100904 299616 100910 299628
rect 256694 299616 256700 299628
rect 256752 299616 256758 299668
rect 97350 299548 97356 299600
rect 97408 299588 97414 299600
rect 279418 299588 279424 299600
rect 97408 299560 279424 299588
rect 97408 299548 97414 299560
rect 279418 299548 279424 299560
rect 279476 299548 279482 299600
rect 88978 299480 88984 299532
rect 89036 299520 89042 299532
rect 303614 299520 303620 299532
rect 89036 299492 303620 299520
rect 89036 299480 89042 299492
rect 303614 299480 303620 299492
rect 303672 299480 303678 299532
rect 59170 298732 59176 298784
rect 59228 298772 59234 298784
rect 124858 298772 124864 298784
rect 59228 298744 124864 298772
rect 59228 298732 59234 298744
rect 124858 298732 124864 298744
rect 124916 298732 124922 298784
rect 113818 298392 113824 298444
rect 113876 298432 113882 298444
rect 169018 298432 169024 298444
rect 113876 298404 169024 298432
rect 113876 298392 113882 298404
rect 169018 298392 169024 298404
rect 169076 298392 169082 298444
rect 87414 298324 87420 298376
rect 87472 298364 87478 298376
rect 211798 298364 211804 298376
rect 87472 298336 211804 298364
rect 87472 298324 87478 298336
rect 211798 298324 211804 298336
rect 211856 298324 211862 298376
rect 66070 298256 66076 298308
rect 66128 298296 66134 298308
rect 203518 298296 203524 298308
rect 66128 298268 203524 298296
rect 66128 298256 66134 298268
rect 203518 298256 203524 298268
rect 203576 298256 203582 298308
rect 106734 298188 106740 298240
rect 106792 298228 106798 298240
rect 269942 298228 269948 298240
rect 106792 298200 269948 298228
rect 106792 298188 106798 298200
rect 269942 298188 269948 298200
rect 270000 298188 270006 298240
rect 111242 298120 111248 298172
rect 111300 298160 111306 298172
rect 278038 298160 278044 298172
rect 111300 298132 278044 298160
rect 111300 298120 111306 298132
rect 278038 298120 278044 298132
rect 278096 298120 278102 298172
rect 439498 298120 439504 298172
rect 439556 298160 439562 298172
rect 580166 298160 580172 298172
rect 439556 298132 580172 298160
rect 439556 298120 439562 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 107562 297440 107568 297492
rect 107620 297480 107626 297492
rect 127066 297480 127072 297492
rect 107620 297452 127072 297480
rect 107620 297440 107626 297452
rect 127066 297440 127072 297452
rect 127124 297440 127130 297492
rect 104158 297372 104164 297424
rect 104216 297412 104222 297424
rect 125686 297412 125692 297424
rect 104216 297384 125692 297412
rect 104216 297372 104222 297384
rect 125686 297372 125692 297384
rect 125744 297372 125750 297424
rect 83550 296896 83556 296948
rect 83608 296936 83614 296948
rect 133138 296936 133144 296948
rect 83608 296908 133144 296936
rect 83608 296896 83614 296908
rect 133138 296896 133144 296908
rect 133196 296896 133202 296948
rect 57882 296828 57888 296880
rect 57940 296868 57946 296880
rect 100018 296868 100024 296880
rect 57940 296840 100024 296868
rect 57940 296828 57946 296840
rect 100018 296828 100024 296840
rect 100076 296828 100082 296880
rect 110598 296828 110604 296880
rect 110656 296868 110662 296880
rect 249794 296868 249800 296880
rect 110656 296840 249800 296868
rect 110656 296828 110662 296840
rect 249794 296828 249800 296840
rect 249852 296828 249858 296880
rect 99650 296760 99656 296812
rect 99708 296800 99714 296812
rect 258074 296800 258080 296812
rect 99708 296772 258080 296800
rect 99708 296760 99714 296772
rect 258074 296760 258080 296772
rect 258132 296760 258138 296812
rect 70670 296692 70676 296744
rect 70728 296732 70734 296744
rect 300946 296732 300952 296744
rect 70728 296704 300952 296732
rect 70728 296692 70734 296704
rect 300946 296692 300952 296704
rect 301004 296692 301010 296744
rect 103422 295944 103428 295996
rect 103480 295984 103486 295996
rect 323578 295984 323584 295996
rect 103480 295956 323584 295984
rect 103480 295944 103486 295956
rect 323578 295944 323584 295956
rect 323636 295944 323642 295996
rect 82906 295604 82912 295656
rect 82964 295644 82970 295656
rect 135898 295644 135904 295656
rect 82964 295616 135904 295644
rect 82964 295604 82970 295616
rect 135898 295604 135904 295616
rect 135956 295604 135962 295656
rect 104250 295536 104256 295588
rect 104308 295576 104314 295588
rect 104802 295576 104808 295588
rect 104308 295548 104808 295576
rect 104308 295536 104314 295548
rect 104802 295536 104808 295548
rect 104860 295576 104866 295588
rect 160738 295576 160744 295588
rect 104860 295548 160744 295576
rect 104860 295536 104866 295548
rect 160738 295536 160744 295548
rect 160796 295536 160802 295588
rect 91922 295468 91928 295520
rect 91980 295508 91986 295520
rect 213270 295508 213276 295520
rect 91980 295480 213276 295508
rect 91980 295468 91986 295480
rect 213270 295468 213276 295480
rect 213328 295468 213334 295520
rect 102226 295400 102232 295452
rect 102284 295440 102290 295452
rect 234614 295440 234620 295452
rect 102284 295412 234620 295440
rect 102284 295400 102290 295412
rect 234614 295400 234620 295412
rect 234672 295400 234678 295452
rect 117038 295332 117044 295384
rect 117096 295372 117102 295384
rect 311894 295372 311900 295384
rect 117096 295344 311900 295372
rect 117096 295332 117102 295344
rect 311894 295332 311900 295344
rect 311952 295332 311958 295384
rect 72602 295264 72608 295316
rect 72660 295304 72666 295316
rect 75270 295304 75276 295316
rect 72660 295276 75276 295304
rect 72660 295264 72666 295276
rect 75270 295264 75276 295276
rect 75328 295264 75334 295316
rect 54938 294720 54944 294772
rect 54996 294760 55002 294772
rect 91278 294760 91284 294772
rect 54996 294732 91284 294760
rect 54996 294720 55002 294732
rect 91278 294720 91284 294732
rect 91336 294720 91342 294772
rect 70026 294652 70032 294704
rect 70084 294692 70090 294704
rect 112438 294692 112444 294704
rect 70084 294664 112444 294692
rect 70084 294652 70090 294664
rect 112438 294652 112444 294664
rect 112496 294652 112502 294704
rect 77110 294584 77116 294636
rect 77168 294624 77174 294636
rect 146478 294624 146484 294636
rect 77168 294596 146484 294624
rect 77168 294584 77174 294596
rect 146478 294584 146484 294596
rect 146536 294624 146542 294636
rect 428458 294624 428464 294636
rect 146536 294596 428464 294624
rect 146536 294584 146542 294596
rect 428458 294584 428464 294596
rect 428516 294584 428522 294636
rect 71314 294312 71320 294364
rect 71372 294352 71378 294364
rect 72510 294352 72516 294364
rect 71372 294324 72516 294352
rect 71372 294312 71378 294324
rect 72510 294312 72516 294324
rect 72568 294312 72574 294364
rect 73154 294312 73160 294364
rect 73212 294352 73218 294364
rect 73614 294352 73620 294364
rect 73212 294324 73620 294352
rect 73212 294312 73218 294324
rect 73614 294312 73620 294324
rect 73672 294312 73678 294364
rect 84286 294312 84292 294364
rect 84344 294352 84350 294364
rect 85206 294352 85212 294364
rect 84344 294324 85212 294352
rect 84344 294312 84350 294324
rect 85206 294312 85212 294324
rect 85264 294312 85270 294364
rect 93946 294312 93952 294364
rect 94004 294352 94010 294364
rect 94774 294352 94780 294364
rect 94004 294324 94780 294352
rect 94004 294312 94010 294324
rect 94774 294312 94780 294324
rect 94832 294312 94838 294364
rect 100018 294312 100024 294364
rect 100076 294352 100082 294364
rect 101582 294352 101588 294364
rect 100076 294324 101588 294352
rect 100076 294312 100082 294324
rect 101582 294312 101588 294324
rect 101640 294312 101646 294364
rect 104894 294312 104900 294364
rect 104952 294352 104958 294364
rect 105814 294352 105820 294364
rect 104952 294324 105820 294352
rect 104952 294312 104958 294324
rect 105814 294312 105820 294324
rect 105872 294312 105878 294364
rect 109954 294244 109960 294296
rect 110012 294284 110018 294296
rect 122926 294284 122932 294296
rect 110012 294256 122932 294284
rect 110012 294244 110018 294256
rect 122926 294244 122932 294256
rect 122984 294284 122990 294296
rect 123662 294284 123668 294296
rect 122984 294256 123668 294284
rect 122984 294244 122990 294256
rect 123662 294244 123668 294256
rect 123720 294244 123726 294296
rect 102870 294176 102876 294228
rect 102928 294216 102934 294228
rect 144178 294216 144184 294228
rect 102928 294188 144184 294216
rect 102928 294176 102934 294188
rect 144178 294176 144184 294188
rect 144236 294176 144242 294228
rect 97074 294108 97080 294160
rect 97132 294148 97138 294160
rect 159450 294148 159456 294160
rect 97132 294120 159456 294148
rect 97132 294108 97138 294120
rect 159450 294108 159456 294120
rect 159508 294108 159514 294160
rect 65518 294040 65524 294092
rect 65576 294080 65582 294092
rect 79042 294080 79048 294092
rect 65576 294052 79048 294080
rect 65576 294040 65582 294052
rect 79042 294040 79048 294052
rect 79100 294040 79106 294092
rect 108022 294040 108028 294092
rect 108080 294080 108086 294092
rect 222838 294080 222844 294092
rect 108080 294052 222844 294080
rect 108080 294040 108086 294052
rect 222838 294040 222844 294052
rect 222896 294040 222902 294092
rect 34330 293972 34336 294024
rect 34388 294012 34394 294024
rect 96430 294012 96436 294024
rect 34388 293984 96436 294012
rect 34388 293972 34394 293984
rect 96430 293972 96436 293984
rect 96488 293972 96494 294024
rect 113818 293972 113824 294024
rect 113876 294012 113882 294024
rect 314654 294012 314660 294024
rect 113876 293984 314660 294012
rect 113876 293972 113882 293984
rect 314654 293972 314660 293984
rect 314712 293972 314718 294024
rect 2774 293156 2780 293208
rect 2832 293196 2838 293208
rect 4798 293196 4804 293208
rect 2832 293168 4804 293196
rect 2832 293156 2838 293168
rect 4798 293156 4804 293168
rect 4856 293156 4862 293208
rect 118602 293020 118608 293072
rect 118660 293060 118666 293072
rect 120074 293060 120080 293072
rect 118660 293032 120080 293060
rect 118660 293020 118666 293032
rect 120074 293020 120080 293032
rect 120132 293020 120138 293072
rect 93854 292816 93860 292868
rect 93912 292856 93918 292868
rect 142798 292856 142804 292868
rect 93912 292828 142804 292856
rect 93912 292816 93918 292828
rect 142798 292816 142804 292828
rect 142856 292816 142862 292868
rect 69106 292748 69112 292800
rect 69164 292788 69170 292800
rect 199378 292788 199384 292800
rect 69164 292760 199384 292788
rect 69164 292748 69170 292760
rect 199378 292748 199384 292760
rect 199436 292748 199442 292800
rect 75178 292680 75184 292732
rect 75236 292720 75242 292732
rect 218698 292720 218704 292732
rect 75236 292692 218704 292720
rect 75236 292680 75242 292692
rect 218698 292680 218704 292692
rect 218756 292680 218762 292732
rect 51166 292612 51172 292664
rect 51224 292652 51230 292664
rect 97074 292652 97080 292664
rect 51224 292624 97080 292652
rect 51224 292612 51230 292624
rect 97074 292612 97080 292624
rect 97132 292612 97138 292664
rect 103514 292612 103520 292664
rect 103572 292652 103578 292664
rect 273898 292652 273904 292664
rect 103572 292624 273904 292652
rect 103572 292612 103578 292624
rect 273898 292612 273904 292624
rect 273956 292612 273962 292664
rect 11698 292544 11704 292596
rect 11756 292584 11762 292596
rect 92566 292584 92572 292596
rect 11756 292556 92572 292584
rect 11756 292544 11762 292556
rect 92566 292544 92572 292556
rect 92624 292584 92630 292596
rect 93762 292584 93768 292596
rect 92624 292556 93768 292584
rect 92624 292544 92630 292556
rect 93762 292544 93768 292556
rect 93820 292584 93826 292596
rect 352558 292584 352564 292596
rect 93820 292556 352564 292584
rect 93820 292544 93826 292556
rect 352558 292544 352564 292556
rect 352616 292544 352622 292596
rect 51074 292476 51080 292528
rect 51132 292516 51138 292528
rect 52178 292516 52184 292528
rect 51132 292488 52184 292516
rect 51132 292476 51138 292488
rect 52178 292476 52184 292488
rect 52236 292516 52242 292528
rect 65518 292516 65524 292528
rect 52236 292488 65524 292516
rect 52236 292476 52242 292488
rect 65518 292476 65524 292488
rect 65576 292476 65582 292528
rect 84286 291864 84292 291916
rect 84344 291904 84350 291916
rect 84344 291876 93854 291904
rect 84344 291864 84350 291876
rect 4062 291796 4068 291848
rect 4120 291836 4126 291848
rect 51074 291836 51080 291848
rect 4120 291808 51080 291836
rect 4120 291796 4126 291808
rect 51074 291796 51080 291808
rect 51132 291796 51138 291848
rect 93826 291360 93854 291876
rect 104434 291864 104440 291916
rect 104492 291864 104498 291916
rect 112806 291864 112812 291916
rect 112864 291904 112870 291916
rect 119706 291904 119712 291916
rect 112864 291876 119712 291904
rect 112864 291864 112870 291876
rect 119706 291864 119712 291876
rect 119764 291864 119770 291916
rect 104452 291428 104480 291864
rect 121546 291796 121552 291848
rect 121604 291836 121610 291848
rect 124122 291836 124128 291848
rect 121604 291808 124128 291836
rect 121604 291796 121610 291808
rect 124122 291796 124128 291808
rect 124180 291836 124186 291848
rect 129642 291836 129648 291848
rect 124180 291808 129648 291836
rect 124180 291796 124186 291808
rect 129642 291796 129648 291808
rect 129700 291796 129706 291848
rect 273990 291428 273996 291440
rect 104452 291400 273996 291428
rect 273990 291388 273996 291400
rect 274048 291388 274054 291440
rect 178770 291360 178776 291372
rect 93826 291332 178776 291360
rect 178770 291320 178776 291332
rect 178828 291320 178834 291372
rect 119706 291252 119712 291304
rect 119764 291292 119770 291304
rect 260834 291292 260840 291304
rect 119764 291264 260840 291292
rect 119764 291252 119770 291264
rect 260834 291252 260840 291264
rect 260892 291252 260898 291304
rect 22738 290436 22744 290488
rect 22796 290476 22802 290488
rect 67634 290476 67640 290488
rect 22796 290448 67640 290476
rect 22796 290436 22802 290448
rect 67634 290436 67640 290448
rect 67692 290436 67698 290488
rect 121546 289892 121552 289944
rect 121604 289932 121610 289944
rect 225598 289932 225604 289944
rect 121604 289904 225604 289932
rect 121604 289892 121610 289904
rect 225598 289892 225604 289904
rect 225656 289892 225662 289944
rect 121638 289824 121644 289876
rect 121696 289864 121702 289876
rect 253934 289864 253940 289876
rect 121696 289836 253940 289864
rect 121696 289824 121702 289836
rect 253934 289824 253940 289836
rect 253992 289824 253998 289876
rect 121730 289144 121736 289196
rect 121788 289184 121794 289196
rect 198090 289184 198096 289196
rect 121788 289156 198096 289184
rect 121788 289144 121794 289156
rect 198090 289144 198096 289156
rect 198148 289144 198154 289196
rect 121822 289076 121828 289128
rect 121880 289116 121886 289128
rect 122006 289116 122012 289128
rect 121880 289088 122012 289116
rect 121880 289076 121886 289088
rect 122006 289076 122012 289088
rect 122064 289116 122070 289128
rect 452654 289116 452660 289128
rect 122064 289088 452660 289116
rect 122064 289076 122070 289088
rect 452654 289076 452660 289088
rect 452712 289116 452718 289128
rect 453298 289116 453304 289128
rect 452712 289088 453304 289116
rect 452712 289076 452718 289088
rect 453298 289076 453304 289088
rect 453356 289076 453362 289128
rect 50982 288396 50988 288448
rect 51040 288436 51046 288448
rect 67634 288436 67640 288448
rect 51040 288408 67640 288436
rect 51040 288396 51046 288408
rect 67634 288396 67640 288408
rect 67692 288396 67698 288448
rect 121638 288396 121644 288448
rect 121696 288436 121702 288448
rect 233878 288436 233884 288448
rect 121696 288408 233884 288436
rect 121696 288396 121702 288408
rect 233878 288396 233884 288408
rect 233936 288396 233942 288448
rect 66162 288328 66168 288380
rect 66220 288368 66226 288380
rect 67726 288368 67732 288380
rect 66220 288340 67732 288368
rect 66220 288328 66226 288340
rect 67726 288328 67732 288340
rect 67784 288328 67790 288380
rect 121546 288328 121552 288380
rect 121604 288368 121610 288380
rect 142430 288368 142436 288380
rect 121604 288340 142436 288368
rect 121604 288328 121610 288340
rect 142430 288328 142436 288340
rect 142488 288368 142494 288380
rect 143442 288368 143448 288380
rect 142488 288340 143448 288368
rect 142488 288328 142494 288340
rect 143442 288328 143448 288340
rect 143500 288328 143506 288380
rect 66070 288260 66076 288312
rect 66128 288300 66134 288312
rect 68186 288300 68192 288312
rect 66128 288272 68192 288300
rect 66128 288260 66134 288272
rect 68186 288260 68192 288272
rect 68244 288260 68250 288312
rect 129734 287716 129740 287768
rect 129792 287756 129798 287768
rect 282270 287756 282276 287768
rect 129792 287728 282276 287756
rect 129792 287716 129798 287728
rect 282270 287716 282276 287728
rect 282328 287716 282334 287768
rect 143442 287648 143448 287700
rect 143500 287688 143506 287700
rect 360838 287688 360844 287700
rect 143500 287660 360844 287688
rect 143500 287648 143506 287660
rect 360838 287648 360844 287660
rect 360896 287648 360902 287700
rect 121454 286628 121460 286680
rect 121512 286668 121518 286680
rect 121638 286668 121644 286680
rect 121512 286640 121644 286668
rect 121512 286628 121518 286640
rect 121638 286628 121644 286640
rect 121696 286628 121702 286680
rect 121454 286492 121460 286544
rect 121512 286532 121518 286544
rect 125686 286532 125692 286544
rect 121512 286504 125692 286532
rect 121512 286492 121518 286504
rect 125686 286492 125692 286504
rect 125744 286492 125750 286544
rect 121546 286424 121552 286476
rect 121604 286464 121610 286476
rect 128446 286464 128452 286476
rect 121604 286436 128452 286464
rect 121604 286424 121610 286436
rect 128446 286424 128452 286436
rect 128504 286424 128510 286476
rect 121638 286356 121644 286408
rect 121696 286396 121702 286408
rect 130378 286396 130384 286408
rect 121696 286368 130384 286396
rect 121696 286356 121702 286368
rect 130378 286356 130384 286368
rect 130436 286356 130442 286408
rect 122282 286288 122288 286340
rect 122340 286328 122346 286340
rect 287330 286328 287336 286340
rect 122340 286300 287336 286328
rect 122340 286288 122346 286300
rect 287330 286288 287336 286300
rect 287388 286288 287394 286340
rect 125686 284928 125692 284980
rect 125744 284968 125750 284980
rect 305638 284968 305644 284980
rect 125744 284940 305644 284968
rect 125744 284928 125750 284940
rect 305638 284928 305644 284940
rect 305696 284928 305702 284980
rect 121454 284384 121460 284436
rect 121512 284424 121518 284436
rect 293954 284424 293960 284436
rect 121512 284396 293960 284424
rect 121512 284384 121518 284396
rect 293954 284384 293960 284396
rect 294012 284384 294018 284436
rect 49418 284316 49424 284368
rect 49476 284356 49482 284368
rect 67634 284356 67640 284368
rect 49476 284328 67640 284356
rect 49476 284316 49482 284328
rect 67634 284316 67640 284328
rect 67692 284316 67698 284368
rect 120902 284316 120908 284368
rect 120960 284356 120966 284368
rect 414658 284356 414664 284368
rect 120960 284328 414664 284356
rect 120960 284316 120966 284328
rect 414658 284316 414664 284328
rect 414716 284316 414722 284368
rect 49602 284248 49608 284300
rect 49660 284288 49666 284300
rect 67726 284288 67732 284300
rect 49660 284260 67732 284288
rect 49660 284248 49666 284260
rect 67726 284248 67732 284260
rect 67784 284248 67790 284300
rect 148318 283568 148324 283620
rect 148376 283608 148382 283620
rect 365714 283608 365720 283620
rect 148376 283580 365720 283608
rect 148376 283568 148382 283580
rect 365714 283568 365720 283580
rect 365772 283568 365778 283620
rect 121454 282888 121460 282940
rect 121512 282928 121518 282940
rect 272518 282928 272524 282940
rect 121512 282900 272524 282928
rect 121512 282888 121518 282900
rect 272518 282888 272524 282900
rect 272576 282888 272582 282940
rect 121454 281528 121460 281580
rect 121512 281568 121518 281580
rect 224218 281568 224224 281580
rect 121512 281540 224224 281568
rect 121512 281528 121518 281540
rect 224218 281528 224224 281540
rect 224276 281528 224282 281580
rect 59170 280236 59176 280288
rect 59228 280276 59234 280288
rect 67634 280276 67640 280288
rect 59228 280248 67640 280276
rect 59228 280236 59234 280248
rect 67634 280236 67640 280248
rect 67692 280236 67698 280288
rect 45370 280168 45376 280220
rect 45428 280208 45434 280220
rect 67726 280208 67732 280220
rect 45428 280180 67732 280208
rect 45428 280168 45434 280180
rect 67726 280168 67732 280180
rect 67784 280168 67790 280220
rect 121454 280168 121460 280220
rect 121512 280208 121518 280220
rect 251174 280208 251180 280220
rect 121512 280180 251180 280208
rect 121512 280168 121518 280180
rect 251174 280168 251180 280180
rect 251232 280168 251238 280220
rect 15838 279420 15844 279472
rect 15896 279460 15902 279472
rect 42702 279460 42708 279472
rect 15896 279432 42708 279460
rect 15896 279420 15902 279432
rect 42702 279420 42708 279432
rect 42760 279460 42766 279472
rect 56410 279460 56416 279472
rect 42760 279432 56416 279460
rect 42760 279420 42766 279432
rect 56410 279420 56416 279432
rect 56468 279420 56474 279472
rect 128446 279420 128452 279472
rect 128504 279460 128510 279472
rect 316678 279460 316684 279472
rect 128504 279432 316684 279460
rect 128504 279420 128510 279432
rect 316678 279420 316684 279432
rect 316736 279420 316742 279472
rect 121546 278808 121552 278860
rect 121604 278848 121610 278860
rect 206370 278848 206376 278860
rect 121604 278820 206376 278848
rect 121604 278808 121610 278820
rect 206370 278808 206376 278820
rect 206428 278808 206434 278860
rect 56410 278740 56416 278792
rect 56468 278780 56474 278792
rect 67634 278780 67640 278792
rect 56468 278752 67640 278780
rect 56468 278740 56474 278752
rect 67634 278740 67640 278752
rect 67692 278740 67698 278792
rect 121454 278740 121460 278792
rect 121512 278780 121518 278792
rect 228358 278780 228364 278792
rect 121512 278752 228364 278780
rect 121512 278740 121518 278752
rect 228358 278740 228364 278752
rect 228416 278740 228422 278792
rect 126330 277992 126336 278044
rect 126388 278032 126394 278044
rect 224310 278032 224316 278044
rect 126388 278004 224316 278032
rect 126388 277992 126394 278004
rect 224310 277992 224316 278004
rect 224368 277992 224374 278044
rect 121454 277448 121460 277500
rect 121512 277488 121518 277500
rect 278130 277488 278136 277500
rect 121512 277460 278136 277488
rect 121512 277448 121518 277460
rect 278130 277448 278136 277460
rect 278188 277448 278194 277500
rect 48038 277380 48044 277432
rect 48096 277420 48102 277432
rect 67634 277420 67640 277432
rect 48096 277392 67640 277420
rect 48096 277380 48102 277392
rect 67634 277380 67640 277392
rect 67692 277380 67698 277432
rect 121546 277380 121552 277432
rect 121604 277420 121610 277432
rect 280890 277420 280896 277432
rect 121604 277392 280896 277420
rect 121604 277380 121610 277392
rect 280890 277380 280896 277392
rect 280948 277380 280954 277432
rect 60642 276088 60648 276140
rect 60700 276128 60706 276140
rect 67634 276128 67640 276140
rect 60700 276100 67640 276128
rect 60700 276088 60706 276100
rect 67634 276088 67640 276100
rect 67692 276088 67698 276140
rect 121454 276088 121460 276140
rect 121512 276128 121518 276140
rect 311986 276128 311992 276140
rect 121512 276100 311992 276128
rect 121512 276088 121518 276100
rect 311986 276088 311992 276100
rect 312044 276088 312050 276140
rect 53558 276020 53564 276072
rect 53616 276060 53622 276072
rect 67726 276060 67732 276072
rect 53616 276032 67732 276060
rect 53616 276020 53622 276032
rect 67726 276020 67732 276032
rect 67784 276020 67790 276072
rect 121546 276020 121552 276072
rect 121604 276060 121610 276072
rect 122282 276060 122288 276072
rect 121604 276032 122288 276060
rect 121604 276020 121610 276032
rect 122282 276020 122288 276032
rect 122340 276060 122346 276072
rect 418798 276060 418804 276072
rect 122340 276032 418804 276060
rect 122340 276020 122346 276032
rect 418798 276020 418804 276032
rect 418856 276020 418862 276072
rect 124122 275272 124128 275324
rect 124180 275312 124186 275324
rect 419534 275312 419540 275324
rect 124180 275284 419540 275312
rect 124180 275272 124186 275284
rect 419534 275272 419540 275284
rect 419592 275272 419598 275324
rect 49510 274728 49516 274780
rect 49568 274768 49574 274780
rect 67634 274768 67640 274780
rect 49568 274740 67640 274768
rect 49568 274728 49574 274740
rect 67634 274728 67640 274740
rect 67692 274728 67698 274780
rect 123570 274728 123576 274780
rect 123628 274768 123634 274780
rect 129826 274768 129832 274780
rect 123628 274740 129832 274768
rect 123628 274728 123634 274740
rect 129826 274728 129832 274740
rect 129884 274728 129890 274780
rect 41230 274660 41236 274712
rect 41288 274700 41294 274712
rect 67726 274700 67732 274712
rect 41288 274672 67732 274700
rect 41288 274660 41294 274672
rect 67726 274660 67732 274672
rect 67784 274660 67790 274712
rect 121454 274660 121460 274712
rect 121512 274700 121518 274712
rect 234706 274700 234712 274712
rect 121512 274672 234712 274700
rect 121512 274660 121518 274672
rect 234706 274660 234712 274672
rect 234764 274660 234770 274712
rect 282178 273912 282184 273964
rect 282236 273952 282242 273964
rect 308398 273952 308404 273964
rect 282236 273924 308404 273952
rect 282236 273912 282242 273924
rect 308398 273912 308404 273924
rect 308456 273912 308462 273964
rect 64598 273232 64604 273284
rect 64656 273272 64662 273284
rect 67634 273272 67640 273284
rect 64656 273244 67640 273272
rect 64656 273232 64662 273244
rect 67634 273232 67640 273244
rect 67692 273232 67698 273284
rect 121454 273232 121460 273284
rect 121512 273272 121518 273284
rect 200850 273272 200856 273284
rect 121512 273244 200856 273272
rect 121512 273232 121518 273244
rect 200850 273232 200856 273244
rect 200908 273232 200914 273284
rect 121454 272484 121460 272536
rect 121512 272524 121518 272536
rect 123478 272524 123484 272536
rect 121512 272496 123484 272524
rect 121512 272484 121518 272496
rect 123478 272484 123484 272496
rect 123536 272524 123542 272536
rect 448514 272524 448520 272536
rect 123536 272496 448520 272524
rect 123536 272484 123542 272496
rect 448514 272484 448520 272496
rect 448572 272484 448578 272536
rect 65978 271940 65984 271992
rect 66036 271980 66042 271992
rect 68094 271980 68100 271992
rect 66036 271952 68100 271980
rect 66036 271940 66042 271952
rect 68094 271940 68100 271952
rect 68152 271940 68158 271992
rect 64690 271872 64696 271924
rect 64748 271912 64754 271924
rect 67634 271912 67640 271924
rect 64748 271884 67640 271912
rect 64748 271872 64754 271884
rect 67634 271872 67640 271884
rect 67692 271872 67698 271924
rect 121454 271872 121460 271924
rect 121512 271912 121518 271924
rect 173894 271912 173900 271924
rect 121512 271884 173900 271912
rect 121512 271872 121518 271884
rect 173894 271872 173900 271884
rect 173952 271872 173958 271924
rect 59262 271124 59268 271176
rect 59320 271164 59326 271176
rect 67634 271164 67640 271176
rect 59320 271136 67640 271164
rect 59320 271124 59326 271136
rect 67634 271124 67640 271136
rect 67692 271124 67698 271176
rect 123662 271124 123668 271176
rect 123720 271164 123726 271176
rect 430942 271164 430948 271176
rect 123720 271136 430948 271164
rect 123720 271124 123726 271136
rect 430942 271124 430948 271136
rect 431000 271124 431006 271176
rect 57606 270512 57612 270564
rect 57664 270552 57670 270564
rect 67726 270552 67732 270564
rect 57664 270524 67732 270552
rect 57664 270512 57670 270524
rect 67726 270512 67732 270524
rect 67784 270512 67790 270564
rect 121454 270512 121460 270564
rect 121512 270552 121518 270564
rect 221458 270552 221464 270564
rect 121512 270524 221464 270552
rect 121512 270512 121518 270524
rect 221458 270512 221464 270524
rect 221516 270512 221522 270564
rect 55030 269152 55036 269204
rect 55088 269192 55094 269204
rect 67726 269192 67732 269204
rect 55088 269164 67732 269192
rect 55088 269152 55094 269164
rect 67726 269152 67732 269164
rect 67784 269152 67790 269204
rect 121454 269152 121460 269204
rect 121512 269192 121518 269204
rect 231946 269192 231952 269204
rect 121512 269164 231952 269192
rect 121512 269152 121518 269164
rect 231946 269152 231952 269164
rect 232004 269152 232010 269204
rect 39942 269084 39948 269136
rect 40000 269124 40006 269136
rect 67634 269124 67640 269136
rect 40000 269096 67640 269124
rect 40000 269084 40006 269096
rect 67634 269084 67640 269096
rect 67692 269084 67698 269136
rect 121546 269084 121552 269136
rect 121604 269124 121610 269136
rect 232130 269124 232136 269136
rect 121604 269096 232136 269124
rect 121604 269084 121610 269096
rect 232130 269084 232136 269096
rect 232188 269084 232194 269136
rect 39850 269016 39856 269068
rect 39908 269056 39914 269068
rect 67726 269056 67732 269068
rect 39908 269028 67732 269056
rect 39908 269016 39914 269028
rect 67726 269016 67732 269028
rect 67784 269016 67790 269068
rect 121454 269016 121460 269068
rect 121512 269056 121518 269068
rect 150434 269056 150440 269068
rect 121512 269028 150440 269056
rect 121512 269016 121518 269028
rect 150434 269016 150440 269028
rect 150492 269016 150498 269068
rect 22002 268336 22008 268388
rect 22060 268376 22066 268388
rect 39850 268376 39856 268388
rect 22060 268348 39856 268376
rect 22060 268336 22066 268348
rect 39850 268336 39856 268348
rect 39908 268336 39914 268388
rect 150434 268336 150440 268388
rect 150492 268376 150498 268388
rect 231210 268376 231216 268388
rect 150492 268348 231216 268376
rect 150492 268336 150498 268348
rect 231210 268336 231216 268348
rect 231268 268336 231274 268388
rect 121546 267724 121552 267776
rect 121604 267764 121610 267776
rect 257338 267764 257344 267776
rect 121604 267736 257344 267764
rect 121604 267724 121610 267736
rect 257338 267724 257344 267736
rect 257396 267724 257402 267776
rect 41138 266976 41144 267028
rect 41196 267016 41202 267028
rect 60182 267016 60188 267028
rect 41196 266988 60188 267016
rect 41196 266976 41202 266988
rect 60182 266976 60188 266988
rect 60240 266976 60246 267028
rect 60734 266500 60740 266552
rect 60792 266540 60798 266552
rect 61378 266540 61384 266552
rect 60792 266512 61384 266540
rect 60792 266500 60798 266512
rect 61378 266500 61384 266512
rect 61436 266540 61442 266552
rect 67634 266540 67640 266552
rect 61436 266512 67640 266540
rect 61436 266500 61442 266512
rect 67634 266500 67640 266512
rect 67692 266500 67698 266552
rect 121638 266432 121644 266484
rect 121696 266472 121702 266484
rect 255958 266472 255964 266484
rect 121696 266444 255964 266472
rect 121696 266432 121702 266444
rect 255958 266432 255964 266444
rect 256016 266432 256022 266484
rect 60182 266364 60188 266416
rect 60240 266404 60246 266416
rect 60458 266404 60464 266416
rect 60240 266376 60464 266404
rect 60240 266364 60246 266376
rect 60458 266364 60464 266376
rect 60516 266404 60522 266416
rect 67726 266404 67732 266416
rect 60516 266376 64644 266404
rect 60516 266364 60522 266376
rect 52270 266296 52276 266348
rect 52328 266336 52334 266348
rect 60734 266336 60740 266348
rect 52328 266308 60740 266336
rect 52328 266296 52334 266308
rect 60734 266296 60740 266308
rect 60792 266296 60798 266348
rect 64616 266336 64644 266376
rect 64846 266376 67732 266404
rect 64846 266336 64874 266376
rect 67726 266364 67732 266376
rect 67784 266364 67790 266416
rect 121546 266364 121552 266416
rect 121604 266404 121610 266416
rect 300854 266404 300860 266416
rect 121604 266376 300860 266404
rect 121604 266364 121610 266376
rect 300854 266364 300860 266376
rect 300912 266364 300918 266416
rect 64616 266308 64874 266336
rect 62022 265616 62028 265668
rect 62080 265656 62086 265668
rect 67634 265656 67640 265668
rect 62080 265628 67640 265656
rect 62080 265616 62086 265628
rect 67634 265616 67640 265628
rect 67692 265616 67698 265668
rect 121546 265004 121552 265056
rect 121604 265044 121610 265056
rect 195330 265044 195336 265056
rect 121604 265016 195336 265044
rect 121604 265004 121610 265016
rect 195330 265004 195336 265016
rect 195388 265004 195394 265056
rect 52178 264936 52184 264988
rect 52236 264976 52242 264988
rect 67726 264976 67732 264988
rect 52236 264948 67732 264976
rect 52236 264936 52242 264948
rect 67726 264936 67732 264948
rect 67784 264936 67790 264988
rect 121638 264936 121644 264988
rect 121696 264976 121702 264988
rect 287146 264976 287152 264988
rect 121696 264948 287152 264976
rect 121696 264936 121702 264948
rect 287146 264936 287152 264948
rect 287204 264936 287210 264988
rect 48222 264868 48228 264920
rect 48280 264908 48286 264920
rect 67634 264908 67640 264920
rect 48280 264880 67640 264908
rect 48280 264868 48286 264880
rect 67634 264868 67640 264880
rect 67692 264868 67698 264920
rect 7558 264188 7564 264240
rect 7616 264228 7622 264240
rect 48222 264228 48228 264240
rect 7616 264200 48228 264228
rect 7616 264188 7622 264200
rect 48222 264188 48228 264200
rect 48280 264188 48286 264240
rect 130378 264188 130384 264240
rect 130436 264228 130442 264240
rect 379514 264228 379520 264240
rect 130436 264200 379520 264228
rect 130436 264188 130442 264200
rect 379514 264188 379520 264200
rect 379572 264188 379578 264240
rect 121638 263576 121644 263628
rect 121696 263616 121702 263628
rect 239030 263616 239036 263628
rect 121696 263588 239036 263616
rect 121696 263576 121702 263588
rect 239030 263576 239036 263588
rect 239088 263576 239094 263628
rect 121546 263508 121552 263560
rect 121604 263548 121610 263560
rect 123018 263548 123024 263560
rect 121604 263520 123024 263548
rect 121604 263508 121610 263520
rect 123018 263508 123024 263520
rect 123076 263548 123082 263560
rect 124122 263548 124128 263560
rect 123076 263520 124128 263548
rect 123076 263508 123082 263520
rect 124122 263508 124128 263520
rect 124180 263508 124186 263560
rect 41322 262964 41328 263016
rect 41380 263004 41386 263016
rect 53834 263004 53840 263016
rect 41380 262976 53840 263004
rect 41380 262964 41386 262976
rect 53834 262964 53840 262976
rect 53892 262964 53898 263016
rect 41322 262828 41328 262880
rect 41380 262868 41386 262880
rect 66898 262868 66904 262880
rect 41380 262840 66904 262868
rect 41380 262828 41386 262840
rect 66898 262828 66904 262840
rect 66956 262828 66962 262880
rect 53834 262284 53840 262336
rect 53892 262324 53898 262336
rect 54846 262324 54852 262336
rect 53892 262296 54852 262324
rect 53892 262284 53898 262296
rect 54846 262284 54852 262296
rect 54904 262324 54910 262336
rect 67726 262324 67732 262336
rect 54904 262296 67732 262324
rect 54904 262284 54910 262296
rect 67726 262284 67732 262296
rect 67784 262284 67790 262336
rect 121546 262284 121552 262336
rect 121604 262324 121610 262336
rect 284294 262324 284300 262336
rect 121604 262296 284300 262324
rect 121604 262284 121610 262296
rect 284294 262284 284300 262296
rect 284352 262284 284358 262336
rect 50798 262216 50804 262268
rect 50856 262256 50862 262268
rect 67634 262256 67640 262268
rect 50856 262228 67640 262256
rect 50856 262216 50862 262228
rect 67634 262216 67640 262228
rect 67692 262216 67698 262268
rect 134702 262216 134708 262268
rect 134760 262256 134766 262268
rect 454034 262256 454040 262268
rect 134760 262228 454040 262256
rect 134760 262216 134766 262228
rect 454034 262216 454040 262228
rect 454092 262216 454098 262268
rect 121546 262148 121552 262200
rect 121604 262188 121610 262200
rect 140774 262188 140780 262200
rect 121604 262160 140780 262188
rect 121604 262148 121610 262160
rect 140774 262148 140780 262160
rect 140832 262148 140838 262200
rect 140774 261468 140780 261520
rect 140832 261508 140838 261520
rect 371878 261508 371884 261520
rect 140832 261480 371884 261508
rect 140832 261468 140838 261480
rect 371878 261468 371884 261480
rect 371936 261468 371942 261520
rect 48222 260856 48228 260908
rect 48280 260896 48286 260908
rect 67726 260896 67732 260908
rect 48280 260868 67732 260896
rect 48280 260856 48286 260868
rect 67726 260856 67732 260868
rect 67784 260856 67790 260908
rect 121638 260856 121644 260908
rect 121696 260896 121702 260908
rect 304994 260896 305000 260908
rect 121696 260868 305000 260896
rect 121696 260856 121702 260868
rect 304994 260856 305000 260868
rect 305052 260856 305058 260908
rect 56502 260788 56508 260840
rect 56560 260828 56566 260840
rect 67634 260828 67640 260840
rect 56560 260800 67640 260828
rect 56560 260788 56566 260800
rect 67634 260788 67640 260800
rect 67692 260788 67698 260840
rect 121546 260788 121552 260840
rect 121604 260828 121610 260840
rect 134702 260828 134708 260840
rect 121604 260800 134708 260828
rect 121604 260788 121610 260800
rect 134702 260788 134708 260800
rect 134760 260788 134766 260840
rect 124122 260108 124128 260160
rect 124180 260148 124186 260160
rect 432138 260148 432144 260160
rect 124180 260120 432144 260148
rect 124180 260108 124186 260120
rect 432138 260108 432144 260120
rect 432196 260108 432202 260160
rect 121546 259496 121552 259548
rect 121604 259536 121610 259548
rect 248414 259536 248420 259548
rect 121604 259508 248420 259536
rect 121604 259496 121610 259508
rect 248414 259496 248420 259508
rect 248472 259496 248478 259548
rect 63126 259428 63132 259480
rect 63184 259468 63190 259480
rect 67634 259468 67640 259480
rect 63184 259440 67640 259468
rect 63184 259428 63190 259440
rect 67634 259428 67640 259440
rect 67692 259428 67698 259480
rect 137278 259468 137284 259480
rect 137191 259440 137284 259468
rect 137278 259428 137284 259440
rect 137336 259468 137342 259480
rect 370498 259468 370504 259480
rect 137336 259440 370504 259468
rect 137336 259428 137342 259440
rect 370498 259428 370504 259440
rect 370556 259428 370562 259480
rect 121546 259360 121552 259412
rect 121604 259400 121610 259412
rect 137296 259400 137324 259428
rect 121604 259372 137324 259400
rect 121604 259360 121610 259372
rect 119982 259292 119988 259344
rect 120040 259332 120046 259344
rect 121638 259332 121644 259344
rect 120040 259304 121644 259332
rect 120040 259292 120046 259304
rect 121638 259292 121644 259304
rect 121696 259292 121702 259344
rect 63310 258136 63316 258188
rect 63368 258176 63374 258188
rect 67634 258176 67640 258188
rect 63368 258148 67640 258176
rect 63368 258136 63374 258148
rect 67634 258136 67640 258148
rect 67692 258136 67698 258188
rect 52270 258068 52276 258120
rect 52328 258108 52334 258120
rect 67726 258108 67732 258120
rect 52328 258080 67732 258108
rect 52328 258068 52334 258080
rect 67726 258068 67732 258080
rect 67784 258068 67790 258120
rect 121730 258068 121736 258120
rect 121788 258108 121794 258120
rect 280798 258108 280804 258120
rect 121788 258080 280804 258108
rect 121788 258068 121794 258080
rect 280798 258068 280804 258080
rect 280856 258068 280862 258120
rect 485038 258068 485044 258120
rect 485096 258108 485102 258120
rect 580166 258108 580172 258120
rect 485096 258080 580172 258108
rect 485096 258068 485102 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 121454 257864 121460 257916
rect 121512 257904 121518 257916
rect 121730 257904 121736 257916
rect 121512 257876 121736 257904
rect 121512 257864 121518 257876
rect 121730 257864 121736 257876
rect 121788 257864 121794 257916
rect 17218 257320 17224 257372
rect 17276 257360 17282 257372
rect 35710 257360 35716 257372
rect 17276 257332 35716 257360
rect 17276 257320 17282 257332
rect 35710 257320 35716 257332
rect 35768 257360 35774 257372
rect 52454 257360 52460 257372
rect 35768 257332 52460 257360
rect 35768 257320 35774 257332
rect 52454 257320 52460 257332
rect 52512 257320 52518 257372
rect 162210 257320 162216 257372
rect 162268 257360 162274 257372
rect 460934 257360 460940 257372
rect 162268 257332 460940 257360
rect 162268 257320 162274 257332
rect 460934 257320 460940 257332
rect 460992 257320 460998 257372
rect 121270 257048 121276 257100
rect 121328 257088 121334 257100
rect 121638 257088 121644 257100
rect 121328 257060 121644 257088
rect 121328 257048 121334 257060
rect 121638 257048 121644 257060
rect 121696 257048 121702 257100
rect 61838 256776 61844 256828
rect 61896 256816 61902 256828
rect 67634 256816 67640 256828
rect 61896 256788 67640 256816
rect 61896 256776 61902 256788
rect 67634 256776 67640 256788
rect 67692 256776 67698 256828
rect 52454 256708 52460 256760
rect 52512 256748 52518 256760
rect 53466 256748 53472 256760
rect 52512 256720 53472 256748
rect 52512 256708 52518 256720
rect 53466 256708 53472 256720
rect 53524 256748 53530 256760
rect 67726 256748 67732 256760
rect 53524 256720 67732 256748
rect 53524 256708 53530 256720
rect 67726 256708 67732 256720
rect 67784 256708 67790 256760
rect 121454 256708 121460 256760
rect 121512 256748 121518 256760
rect 227162 256748 227168 256760
rect 121512 256720 227168 256748
rect 121512 256708 121518 256720
rect 227162 256708 227168 256720
rect 227220 256708 227226 256760
rect 121638 255960 121644 256012
rect 121696 256000 121702 256012
rect 315298 256000 315304 256012
rect 121696 255972 315304 256000
rect 121696 255960 121702 255972
rect 315298 255960 315304 255972
rect 315356 255960 315362 256012
rect 122834 255756 122840 255808
rect 122892 255796 122898 255808
rect 125594 255796 125600 255808
rect 122892 255768 125600 255796
rect 122892 255756 122898 255768
rect 125594 255756 125600 255768
rect 125652 255756 125658 255808
rect 56318 255348 56324 255400
rect 56376 255388 56382 255400
rect 67634 255388 67640 255400
rect 56376 255360 67640 255388
rect 56376 255348 56382 255360
rect 67634 255348 67640 255360
rect 67692 255348 67698 255400
rect 44082 255280 44088 255332
rect 44140 255320 44146 255332
rect 67726 255320 67732 255332
rect 44140 255292 67732 255320
rect 44140 255280 44146 255292
rect 67726 255280 67732 255292
rect 67784 255280 67790 255332
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 33318 255252 33324 255264
rect 3200 255224 33324 255252
rect 3200 255212 3206 255224
rect 33318 255212 33324 255224
rect 33376 255212 33382 255264
rect 53742 255212 53748 255264
rect 53800 255252 53806 255264
rect 67634 255252 67640 255264
rect 53800 255224 67640 255252
rect 53800 255212 53806 255224
rect 67634 255212 67640 255224
rect 67692 255212 67698 255264
rect 121454 255212 121460 255264
rect 121512 255252 121518 255264
rect 131114 255252 131120 255264
rect 121512 255224 131120 255252
rect 121512 255212 121518 255224
rect 131114 255212 131120 255224
rect 131172 255252 131178 255264
rect 131482 255252 131488 255264
rect 131172 255224 131488 255252
rect 131172 255212 131178 255224
rect 131482 255212 131488 255224
rect 131540 255212 131546 255264
rect 33318 254532 33324 254584
rect 33376 254572 33382 254584
rect 34238 254572 34244 254584
rect 33376 254544 34244 254572
rect 33376 254532 33382 254544
rect 34238 254532 34244 254544
rect 34296 254572 34302 254584
rect 59998 254572 60004 254584
rect 34296 254544 60004 254572
rect 34296 254532 34302 254544
rect 59998 254532 60004 254544
rect 60056 254532 60062 254584
rect 60550 254532 60556 254584
rect 60608 254572 60614 254584
rect 67634 254572 67640 254584
rect 60608 254544 67640 254572
rect 60608 254532 60614 254544
rect 67634 254532 67640 254544
rect 67692 254532 67698 254584
rect 131482 254532 131488 254584
rect 131540 254572 131546 254584
rect 330478 254572 330484 254584
rect 131540 254544 330484 254572
rect 131540 254532 131546 254544
rect 330478 254532 330484 254544
rect 330536 254532 330542 254584
rect 121638 253988 121644 254040
rect 121696 254028 121702 254040
rect 250438 254028 250444 254040
rect 121696 254000 250444 254028
rect 121696 253988 121702 254000
rect 250438 253988 250444 254000
rect 250496 253988 250502 254040
rect 121454 253920 121460 253972
rect 121512 253960 121518 253972
rect 259454 253960 259460 253972
rect 121512 253932 259460 253960
rect 121512 253920 121518 253932
rect 259454 253920 259460 253932
rect 259512 253920 259518 253972
rect 45462 253852 45468 253904
rect 45520 253892 45526 253904
rect 47302 253892 47308 253904
rect 45520 253864 47308 253892
rect 45520 253852 45526 253864
rect 47302 253852 47308 253864
rect 47360 253852 47366 253904
rect 125594 253172 125600 253224
rect 125652 253212 125658 253224
rect 356054 253212 356060 253224
rect 125652 253184 356060 253212
rect 125652 253172 125658 253184
rect 356054 253172 356060 253184
rect 356112 253172 356118 253224
rect 121638 252628 121644 252680
rect 121696 252668 121702 252680
rect 220262 252668 220268 252680
rect 121696 252640 220268 252668
rect 121696 252628 121702 252640
rect 220262 252628 220268 252640
rect 220320 252628 220326 252680
rect 46934 252560 46940 252612
rect 46992 252600 46998 252612
rect 47302 252600 47308 252612
rect 46992 252572 47308 252600
rect 46992 252560 46998 252572
rect 47302 252560 47308 252572
rect 47360 252600 47366 252612
rect 69014 252600 69020 252612
rect 47360 252572 69020 252600
rect 47360 252560 47366 252572
rect 69014 252560 69020 252572
rect 69072 252560 69078 252612
rect 121454 252560 121460 252612
rect 121512 252600 121518 252612
rect 283098 252600 283104 252612
rect 121512 252572 283104 252600
rect 121512 252560 121518 252572
rect 283098 252560 283104 252572
rect 283156 252560 283162 252612
rect 178678 251880 178684 251932
rect 178736 251920 178742 251932
rect 271230 251920 271236 251932
rect 178736 251892 271236 251920
rect 178736 251880 178742 251892
rect 271230 251880 271236 251892
rect 271288 251880 271294 251932
rect 121730 251812 121736 251864
rect 121788 251852 121794 251864
rect 407758 251852 407764 251864
rect 121788 251824 407764 251852
rect 121788 251812 121794 251824
rect 407758 251812 407764 251824
rect 407816 251812 407822 251864
rect 54938 251200 54944 251252
rect 54996 251240 55002 251252
rect 67634 251240 67640 251252
rect 54996 251212 67640 251240
rect 54996 251200 55002 251212
rect 67634 251200 67640 251212
rect 67692 251200 67698 251252
rect 121454 251200 121460 251252
rect 121512 251240 121518 251252
rect 310514 251240 310520 251252
rect 121512 251212 310520 251240
rect 121512 251200 121518 251212
rect 310514 251200 310520 251212
rect 310572 251200 310578 251252
rect 169018 250520 169024 250572
rect 169076 250560 169082 250572
rect 264330 250560 264336 250572
rect 169076 250532 264336 250560
rect 169076 250520 169082 250532
rect 264330 250520 264336 250532
rect 264388 250520 264394 250572
rect 135898 250452 135904 250504
rect 135956 250492 135962 250504
rect 238846 250492 238852 250504
rect 135956 250464 238852 250492
rect 135956 250452 135962 250464
rect 238846 250452 238852 250464
rect 238904 250452 238910 250504
rect 53742 249840 53748 249892
rect 53800 249880 53806 249892
rect 67726 249880 67732 249892
rect 53800 249852 67732 249880
rect 53800 249840 53806 249852
rect 67726 249840 67732 249852
rect 67784 249840 67790 249892
rect 120074 249840 120080 249892
rect 120132 249880 120138 249892
rect 122834 249880 122840 249892
rect 120132 249852 122840 249880
rect 120132 249840 120138 249852
rect 122834 249840 122840 249852
rect 122892 249840 122898 249892
rect 50890 249772 50896 249824
rect 50948 249812 50954 249824
rect 67634 249812 67640 249824
rect 50948 249784 67640 249812
rect 50948 249772 50954 249784
rect 67634 249772 67640 249784
rect 67692 249772 67698 249824
rect 121454 249772 121460 249824
rect 121512 249812 121518 249824
rect 221550 249812 221556 249824
rect 121512 249784 221556 249812
rect 121512 249772 121518 249784
rect 221550 249772 221556 249784
rect 221608 249772 221614 249824
rect 121638 249364 121644 249416
rect 121696 249404 121702 249416
rect 122742 249404 122748 249416
rect 121696 249376 122748 249404
rect 121696 249364 121702 249376
rect 122742 249364 122748 249376
rect 122800 249404 122806 249416
rect 124214 249404 124220 249416
rect 122800 249376 124220 249404
rect 122800 249364 122806 249376
rect 124214 249364 124220 249376
rect 124272 249364 124278 249416
rect 56502 249092 56508 249144
rect 56560 249132 56566 249144
rect 68278 249132 68284 249144
rect 56560 249104 68284 249132
rect 56560 249092 56566 249104
rect 68278 249092 68284 249104
rect 68336 249092 68342 249144
rect 43438 249024 43444 249076
rect 43496 249064 43502 249076
rect 59078 249064 59084 249076
rect 43496 249036 59084 249064
rect 43496 249024 43502 249036
rect 59078 249024 59084 249036
rect 59136 249024 59142 249076
rect 65886 249024 65892 249076
rect 65944 249064 65950 249076
rect 68094 249064 68100 249076
rect 65944 249036 68100 249064
rect 65944 249024 65950 249036
rect 68094 249024 68100 249036
rect 68152 249024 68158 249076
rect 173158 249024 173164 249076
rect 173216 249064 173222 249076
rect 400858 249064 400864 249076
rect 173216 249036 400864 249064
rect 173216 249024 173222 249036
rect 400858 249024 400864 249036
rect 400916 249024 400922 249076
rect 64506 248480 64512 248532
rect 64564 248520 64570 248532
rect 67634 248520 67640 248532
rect 64564 248492 67640 248520
rect 64564 248480 64570 248492
rect 67634 248480 67640 248492
rect 67692 248480 67698 248532
rect 59078 248412 59084 248464
rect 59136 248452 59142 248464
rect 67726 248452 67732 248464
rect 59136 248424 67732 248452
rect 59136 248412 59142 248424
rect 67726 248412 67732 248424
rect 67784 248412 67790 248464
rect 121454 248412 121460 248464
rect 121512 248452 121518 248464
rect 196710 248452 196716 248464
rect 121512 248424 196716 248452
rect 121512 248412 121518 248424
rect 196710 248412 196716 248424
rect 196768 248412 196774 248464
rect 159450 247732 159456 247784
rect 159508 247772 159514 247784
rect 367094 247772 367100 247784
rect 159508 247744 367100 247772
rect 159508 247732 159514 247744
rect 367094 247732 367100 247744
rect 367152 247732 367158 247784
rect 122834 247664 122840 247716
rect 122892 247704 122898 247716
rect 375374 247704 375380 247716
rect 122892 247676 375380 247704
rect 122892 247664 122898 247676
rect 375374 247664 375380 247676
rect 375432 247664 375438 247716
rect 63218 247120 63224 247172
rect 63276 247160 63282 247172
rect 67726 247160 67732 247172
rect 63276 247132 67732 247160
rect 63276 247120 63282 247132
rect 67726 247120 67732 247132
rect 67784 247120 67790 247172
rect 61930 247052 61936 247104
rect 61988 247092 61994 247104
rect 67634 247092 67640 247104
rect 61988 247064 67640 247092
rect 61988 247052 61994 247064
rect 67634 247052 67640 247064
rect 67692 247052 67698 247104
rect 121454 247052 121460 247104
rect 121512 247092 121518 247104
rect 240134 247092 240140 247104
rect 121512 247064 240140 247092
rect 121512 247052 121518 247064
rect 240134 247052 240140 247064
rect 240192 247052 240198 247104
rect 121454 246304 121460 246356
rect 121512 246344 121518 246356
rect 431954 246344 431960 246356
rect 121512 246316 431960 246344
rect 121512 246304 121518 246316
rect 431954 246304 431960 246316
rect 432012 246304 432018 246356
rect 121546 245692 121552 245744
rect 121604 245732 121610 245744
rect 234798 245732 234804 245744
rect 121604 245704 234804 245732
rect 121604 245692 121610 245704
rect 234798 245692 234804 245704
rect 234856 245692 234862 245744
rect 121454 245624 121460 245676
rect 121512 245664 121518 245676
rect 242894 245664 242900 245676
rect 121512 245636 242900 245664
rect 121512 245624 121518 245636
rect 242894 245624 242900 245636
rect 242952 245624 242958 245676
rect 121546 244332 121552 244384
rect 121604 244372 121610 244384
rect 258718 244372 258724 244384
rect 121604 244344 258724 244372
rect 121604 244332 121610 244344
rect 258718 244332 258724 244344
rect 258776 244332 258782 244384
rect 64782 244264 64788 244316
rect 64840 244304 64846 244316
rect 67634 244304 67640 244316
rect 64840 244276 67640 244304
rect 64840 244264 64846 244276
rect 67634 244264 67640 244276
rect 67692 244264 67698 244316
rect 126238 244264 126244 244316
rect 126296 244304 126302 244316
rect 579614 244304 579620 244316
rect 126296 244276 579620 244304
rect 126296 244264 126302 244276
rect 579614 244264 579620 244276
rect 579672 244304 579678 244316
rect 579982 244304 579988 244316
rect 579672 244276 579988 244304
rect 579672 244264 579678 244276
rect 579982 244264 579988 244276
rect 580040 244264 580046 244316
rect 121454 244196 121460 244248
rect 121512 244236 121518 244248
rect 142246 244236 142252 244248
rect 121512 244208 142252 244236
rect 121512 244196 121518 244208
rect 142246 244196 142252 244208
rect 142304 244236 142310 244248
rect 143442 244236 143448 244248
rect 142304 244208 143448 244236
rect 142304 244196 142310 244208
rect 143442 244196 143448 244208
rect 143500 244196 143506 244248
rect 143442 243516 143448 243568
rect 143500 243556 143506 243568
rect 311158 243556 311164 243568
rect 143500 243528 311164 243556
rect 143500 243516 143506 243528
rect 311158 243516 311164 243528
rect 311216 243516 311222 243568
rect 66162 242972 66168 243024
rect 66220 243012 66226 243024
rect 67726 243012 67732 243024
rect 66220 242984 67732 243012
rect 66220 242972 66226 242984
rect 67726 242972 67732 242984
rect 67784 242972 67790 243024
rect 121546 242972 121552 243024
rect 121604 243012 121610 243024
rect 279510 243012 279516 243024
rect 121604 242984 279516 243012
rect 121604 242972 121610 242984
rect 279510 242972 279516 242984
rect 279568 242972 279574 243024
rect 67634 242944 67640 242956
rect 59280 242916 67640 242944
rect 48130 242836 48136 242888
rect 48188 242876 48194 242888
rect 58618 242876 58624 242888
rect 48188 242848 58624 242876
rect 48188 242836 48194 242848
rect 58618 242836 58624 242848
rect 58676 242876 58682 242888
rect 59280 242876 59308 242916
rect 67634 242904 67640 242916
rect 67692 242904 67698 242956
rect 124858 242904 124864 242956
rect 124916 242944 124922 242956
rect 413278 242944 413284 242956
rect 124916 242916 413284 242944
rect 124916 242904 124922 242916
rect 413278 242904 413284 242916
rect 413336 242904 413342 242956
rect 58676 242848 59308 242876
rect 58676 242836 58682 242848
rect 121546 242836 121552 242888
rect 121604 242876 121610 242888
rect 128354 242876 128360 242888
rect 121604 242848 128360 242876
rect 121604 242836 121610 242848
rect 128354 242836 128360 242848
rect 128412 242836 128418 242888
rect 121454 242768 121460 242820
rect 121512 242808 121518 242820
rect 126238 242808 126244 242820
rect 121512 242780 126244 242808
rect 121512 242768 121518 242780
rect 126238 242768 126244 242780
rect 126296 242768 126302 242820
rect 122098 242156 122104 242208
rect 122156 242196 122162 242208
rect 433518 242196 433524 242208
rect 122156 242168 433524 242196
rect 122156 242156 122162 242168
rect 433518 242156 433524 242168
rect 433576 242156 433582 242208
rect 66070 241476 66076 241528
rect 66128 241516 66134 241528
rect 68186 241516 68192 241528
rect 66128 241488 68192 241516
rect 66128 241476 66134 241488
rect 68186 241476 68192 241488
rect 68244 241476 68250 241528
rect 121638 240728 121644 240780
rect 121696 240768 121702 240780
rect 182174 240768 182180 240780
rect 121696 240740 182180 240768
rect 121696 240728 121702 240740
rect 182174 240728 182180 240740
rect 182232 240728 182238 240780
rect 121454 240116 121460 240168
rect 121512 240156 121518 240168
rect 241790 240156 241796 240168
rect 121512 240128 241796 240156
rect 121512 240116 121518 240128
rect 241790 240116 241796 240128
rect 241848 240116 241854 240168
rect 3142 240048 3148 240100
rect 3200 240088 3206 240100
rect 37182 240088 37188 240100
rect 3200 240060 37188 240088
rect 3200 240048 3206 240060
rect 37182 240048 37188 240060
rect 37240 240048 37246 240100
rect 69842 240048 69848 240100
rect 69900 240088 69906 240100
rect 133966 240088 133972 240100
rect 69900 240060 133972 240088
rect 69900 240048 69906 240060
rect 133966 240048 133972 240060
rect 134024 240088 134030 240100
rect 134518 240088 134524 240100
rect 134024 240060 134524 240088
rect 134024 240048 134030 240060
rect 134518 240048 134524 240060
rect 134576 240048 134582 240100
rect 117682 239912 117688 239964
rect 117740 239952 117746 239964
rect 124858 239952 124864 239964
rect 117740 239924 124864 239952
rect 117740 239912 117746 239924
rect 124858 239912 124864 239924
rect 124916 239912 124922 239964
rect 75914 239776 75920 239828
rect 75972 239816 75978 239828
rect 77098 239816 77104 239828
rect 75972 239788 77104 239816
rect 75972 239776 75978 239788
rect 77098 239776 77104 239788
rect 77156 239776 77162 239828
rect 77294 239776 77300 239828
rect 77352 239816 77358 239828
rect 78386 239816 78392 239828
rect 77352 239788 78392 239816
rect 77352 239776 77358 239788
rect 78386 239776 78392 239788
rect 78444 239776 78450 239828
rect 80054 239776 80060 239828
rect 80112 239816 80118 239828
rect 80962 239816 80968 239828
rect 80112 239788 80968 239816
rect 80112 239776 80118 239788
rect 80962 239776 80968 239788
rect 81020 239776 81026 239828
rect 86954 239776 86960 239828
rect 87012 239816 87018 239828
rect 88046 239816 88052 239828
rect 87012 239788 88052 239816
rect 87012 239776 87018 239788
rect 88046 239776 88052 239788
rect 88104 239776 88110 239828
rect 89714 239776 89720 239828
rect 89772 239816 89778 239828
rect 90622 239816 90628 239828
rect 89772 239788 90628 239816
rect 89772 239776 89778 239788
rect 90622 239776 90628 239788
rect 90680 239776 90686 239828
rect 95234 239776 95240 239828
rect 95292 239816 95298 239828
rect 96418 239816 96424 239828
rect 95292 239788 96424 239816
rect 95292 239776 95298 239788
rect 96418 239776 96424 239788
rect 96476 239776 96482 239828
rect 96614 239776 96620 239828
rect 96672 239816 96678 239828
rect 97706 239816 97712 239828
rect 96672 239788 97712 239816
rect 96672 239776 96678 239788
rect 97706 239776 97712 239788
rect 97764 239776 97770 239828
rect 104894 239776 104900 239828
rect 104952 239816 104958 239828
rect 106078 239816 106084 239828
rect 104952 239788 106084 239816
rect 104952 239776 104958 239788
rect 106078 239776 106084 239788
rect 106136 239776 106142 239828
rect 114554 239776 114560 239828
rect 114612 239816 114618 239828
rect 115738 239816 115744 239828
rect 114612 239788 115744 239816
rect 114612 239776 114618 239788
rect 115738 239776 115744 239788
rect 115796 239776 115802 239828
rect 64782 239436 64788 239488
rect 64840 239476 64846 239488
rect 78306 239476 78312 239488
rect 64840 239448 78312 239476
rect 64840 239436 64846 239448
rect 78306 239436 78312 239448
rect 78364 239436 78370 239488
rect 37182 239368 37188 239420
rect 37240 239408 37246 239420
rect 88242 239408 88248 239420
rect 37240 239380 88248 239408
rect 37240 239368 37246 239380
rect 88242 239368 88248 239380
rect 88300 239368 88306 239420
rect 231210 239368 231216 239420
rect 231268 239408 231274 239420
rect 411254 239408 411260 239420
rect 231268 239380 411260 239408
rect 231268 239368 231274 239380
rect 411254 239368 411260 239380
rect 411312 239368 411318 239420
rect 74626 239300 74632 239352
rect 74684 239340 74690 239352
rect 75822 239340 75828 239352
rect 74684 239312 75828 239340
rect 74684 239300 74690 239312
rect 75822 239300 75828 239312
rect 75880 239300 75886 239352
rect 93946 239300 93952 239352
rect 94004 239340 94010 239352
rect 95142 239340 95148 239352
rect 94004 239312 95148 239340
rect 94004 239300 94010 239312
rect 95142 239300 95148 239312
rect 95200 239300 95206 239352
rect 59998 238756 60004 238808
rect 60056 238796 60062 238808
rect 111886 238796 111892 238808
rect 60056 238768 111892 238796
rect 60056 238756 60062 238768
rect 111886 238756 111892 238768
rect 111944 238796 111950 238808
rect 112530 238796 112536 238808
rect 111944 238768 112536 238796
rect 111944 238756 111950 238768
rect 112530 238756 112536 238768
rect 112588 238756 112594 238808
rect 116026 238756 116032 238808
rect 116084 238796 116090 238808
rect 117038 238796 117044 238808
rect 116084 238768 117044 238796
rect 116084 238756 116090 238768
rect 117038 238756 117044 238768
rect 117096 238796 117102 238808
rect 127066 238796 127072 238808
rect 117096 238768 127072 238796
rect 117096 238756 117102 238768
rect 127066 238756 127072 238768
rect 127124 238756 127130 238808
rect 3418 238688 3424 238740
rect 3476 238728 3482 238740
rect 86770 238728 86776 238740
rect 3476 238700 86776 238728
rect 3476 238688 3482 238700
rect 86770 238688 86776 238700
rect 86828 238688 86834 238740
rect 88242 238688 88248 238740
rect 88300 238728 88306 238740
rect 103514 238728 103520 238740
rect 88300 238700 103520 238728
rect 88300 238688 88306 238700
rect 103514 238688 103520 238700
rect 103572 238688 103578 238740
rect 114462 238688 114468 238740
rect 114520 238728 114526 238740
rect 132586 238728 132592 238740
rect 114520 238700 132592 238728
rect 114520 238688 114526 238700
rect 132586 238688 132592 238700
rect 132644 238728 132650 238740
rect 133782 238728 133788 238740
rect 132644 238700 133788 238728
rect 132644 238688 132650 238700
rect 133782 238688 133788 238700
rect 133840 238688 133846 238740
rect 57790 238620 57796 238672
rect 57848 238660 57854 238672
rect 86126 238660 86132 238672
rect 57848 238632 86132 238660
rect 57848 238620 57854 238632
rect 86126 238620 86132 238632
rect 86184 238620 86190 238672
rect 57698 238552 57704 238604
rect 57756 238592 57762 238604
rect 72602 238592 72608 238604
rect 57756 238564 72608 238592
rect 57756 238552 57762 238564
rect 72602 238552 72608 238564
rect 72660 238552 72666 238604
rect 86770 238280 86776 238332
rect 86828 238320 86834 238332
rect 98822 238320 98828 238332
rect 86828 238292 98828 238320
rect 86828 238280 86834 238292
rect 98822 238280 98828 238292
rect 98880 238280 98886 238332
rect 105446 238280 105452 238332
rect 105504 238320 105510 238332
rect 178678 238320 178684 238332
rect 105504 238292 178684 238320
rect 105504 238280 105510 238292
rect 178678 238280 178684 238292
rect 178736 238280 178742 238332
rect 100294 238212 100300 238264
rect 100352 238252 100358 238264
rect 233234 238252 233240 238264
rect 100352 238224 233240 238252
rect 100352 238212 100358 238224
rect 233234 238212 233240 238224
rect 233292 238212 233298 238264
rect 69934 238144 69940 238196
rect 69992 238184 69998 238196
rect 288526 238184 288532 238196
rect 69992 238156 288532 238184
rect 69992 238144 69998 238156
rect 288526 238144 288532 238156
rect 288584 238144 288590 238196
rect 70670 238076 70676 238128
rect 70728 238116 70734 238128
rect 313274 238116 313280 238128
rect 70728 238088 313280 238116
rect 70728 238076 70734 238088
rect 313274 238076 313280 238088
rect 313332 238076 313338 238128
rect 72602 238008 72608 238060
rect 72660 238048 72666 238060
rect 86310 238048 86316 238060
rect 72660 238020 86316 238048
rect 72660 238008 72666 238020
rect 86310 238008 86316 238020
rect 86368 238008 86374 238060
rect 98822 238008 98828 238060
rect 98880 238048 98886 238060
rect 99190 238048 99196 238060
rect 98880 238020 99196 238048
rect 98880 238008 98886 238020
rect 99190 238008 99196 238020
rect 99248 238048 99254 238060
rect 128538 238048 128544 238060
rect 99248 238020 128544 238048
rect 99248 238008 99254 238020
rect 128538 238008 128544 238020
rect 128596 238008 128602 238060
rect 133782 238008 133788 238060
rect 133840 238048 133846 238060
rect 434714 238048 434720 238060
rect 133840 238020 434720 238048
rect 133840 238008 133846 238020
rect 434714 238008 434720 238020
rect 434772 238008 434778 238060
rect 103514 237464 103520 237516
rect 103572 237504 103578 237516
rect 104158 237504 104164 237516
rect 103572 237476 104164 237504
rect 103572 237464 103578 237476
rect 104158 237464 104164 237476
rect 104216 237464 104222 237516
rect 85482 237396 85488 237448
rect 85540 237436 85546 237448
rect 86218 237436 86224 237448
rect 85540 237408 86224 237436
rect 85540 237396 85546 237408
rect 86218 237396 86224 237408
rect 86276 237396 86282 237448
rect 102870 237396 102876 237448
rect 102928 237436 102934 237448
rect 105538 237436 105544 237448
rect 102928 237408 105544 237436
rect 102928 237396 102934 237408
rect 105538 237396 105544 237408
rect 105596 237396 105602 237448
rect 69198 237328 69204 237380
rect 69256 237368 69262 237380
rect 138014 237368 138020 237380
rect 69256 237340 138020 237368
rect 69256 237328 69262 237340
rect 138014 237328 138020 237340
rect 138072 237328 138078 237380
rect 52362 237260 52368 237312
rect 52420 237300 52426 237312
rect 81618 237300 81624 237312
rect 52420 237272 81624 237300
rect 52420 237260 52426 237272
rect 81618 237260 81624 237272
rect 81676 237260 81682 237312
rect 99282 237260 99288 237312
rect 99340 237300 99346 237312
rect 123570 237300 123576 237312
rect 99340 237272 123576 237300
rect 99340 237260 99346 237272
rect 123570 237260 123576 237272
rect 123628 237260 123634 237312
rect 66162 236716 66168 236768
rect 66220 236756 66226 236768
rect 276750 236756 276756 236768
rect 66220 236728 276756 236756
rect 66220 236716 66226 236728
rect 276750 236716 276756 236728
rect 276808 236716 276814 236768
rect 138014 236648 138020 236700
rect 138072 236688 138078 236700
rect 385034 236688 385040 236700
rect 138072 236660 385040 236688
rect 138072 236648 138078 236660
rect 385034 236648 385040 236660
rect 385092 236648 385098 236700
rect 81618 235968 81624 236020
rect 81676 236008 81682 236020
rect 82078 236008 82084 236020
rect 81676 235980 82084 236008
rect 81676 235968 81682 235980
rect 82078 235968 82084 235980
rect 82136 235968 82142 236020
rect 110598 235900 110604 235952
rect 110656 235940 110662 235952
rect 111058 235940 111064 235952
rect 110656 235912 111064 235940
rect 110656 235900 110662 235912
rect 111058 235900 111064 235912
rect 111116 235940 111122 235952
rect 136634 235940 136640 235952
rect 111116 235912 136640 235940
rect 111116 235900 111122 235912
rect 136634 235900 136640 235912
rect 136692 235900 136698 235952
rect 61930 235356 61936 235408
rect 61988 235396 61994 235408
rect 245654 235396 245660 235408
rect 61988 235368 245660 235396
rect 61988 235356 61994 235368
rect 245654 235356 245660 235368
rect 245712 235356 245718 235408
rect 231118 235288 231124 235340
rect 231176 235328 231182 235340
rect 446398 235328 446404 235340
rect 231176 235300 446404 235328
rect 231176 235288 231182 235300
rect 446398 235288 446404 235300
rect 446456 235288 446462 235340
rect 57606 235220 57612 235272
rect 57664 235260 57670 235272
rect 290090 235260 290096 235272
rect 57664 235232 290096 235260
rect 57664 235220 57670 235232
rect 290090 235220 290096 235232
rect 290148 235220 290154 235272
rect 46842 234540 46848 234592
rect 46900 234580 46906 234592
rect 118970 234580 118976 234592
rect 46900 234552 118976 234580
rect 46900 234540 46906 234552
rect 118970 234540 118976 234552
rect 119028 234540 119034 234592
rect 53650 234472 53656 234524
rect 53708 234512 53714 234524
rect 91738 234512 91744 234524
rect 53708 234484 91744 234512
rect 53708 234472 53714 234484
rect 91738 234472 91744 234484
rect 91796 234472 91802 234524
rect 118970 234132 118976 234184
rect 119028 234172 119034 234184
rect 119338 234172 119344 234184
rect 119028 234144 119344 234172
rect 119028 234132 119034 234144
rect 119338 234132 119344 234144
rect 119396 234132 119402 234184
rect 108022 233860 108028 233912
rect 108080 233900 108086 233912
rect 284386 233900 284392 233912
rect 108080 233872 284392 233900
rect 108080 233860 108086 233872
rect 284386 233860 284392 233872
rect 284444 233860 284450 233912
rect 84194 233792 84200 233844
rect 84252 233832 84258 233844
rect 84252 233804 84332 233832
rect 84252 233792 84258 233804
rect 84304 233640 84332 233804
rect 84286 233588 84292 233640
rect 84344 233588 84350 233640
rect 55122 233180 55128 233232
rect 55180 233220 55186 233232
rect 109678 233220 109684 233232
rect 55180 233192 109684 233220
rect 55180 233180 55186 233192
rect 109678 233180 109684 233192
rect 109736 233180 109742 233232
rect 52178 232704 52184 232756
rect 52236 232744 52242 232756
rect 157978 232744 157984 232756
rect 52236 232716 157984 232744
rect 52236 232704 52242 232716
rect 157978 232704 157984 232716
rect 158036 232704 158042 232756
rect 78306 232636 78312 232688
rect 78364 232676 78370 232688
rect 222930 232676 222936 232688
rect 78364 232648 222936 232676
rect 78364 232636 78370 232648
rect 222930 232636 222936 232648
rect 222988 232636 222994 232688
rect 69106 232568 69112 232620
rect 69164 232608 69170 232620
rect 281718 232608 281724 232620
rect 69164 232580 281724 232608
rect 69164 232568 69170 232580
rect 281718 232568 281724 232580
rect 281776 232568 281782 232620
rect 107378 232500 107384 232552
rect 107436 232540 107442 232552
rect 411898 232540 411904 232552
rect 107436 232512 411904 232540
rect 107436 232500 107442 232512
rect 411898 232500 411904 232512
rect 411956 232500 411962 232552
rect 74442 231820 74448 231872
rect 74500 231860 74506 231872
rect 75178 231860 75184 231872
rect 74500 231832 75184 231860
rect 74500 231820 74506 231832
rect 75178 231820 75184 231832
rect 75236 231820 75242 231872
rect 93762 231820 93768 231872
rect 93820 231860 93826 231872
rect 94498 231860 94504 231872
rect 93820 231832 94504 231860
rect 93820 231820 93826 231832
rect 94498 231820 94504 231832
rect 94556 231820 94562 231872
rect 349062 231820 349068 231872
rect 349120 231860 349126 231872
rect 580166 231860 580172 231872
rect 349120 231832 580172 231860
rect 349120 231820 349126 231832
rect 580166 231820 580172 231832
rect 580224 231820 580230 231872
rect 101490 231140 101496 231192
rect 101548 231180 101554 231192
rect 229278 231180 229284 231192
rect 101548 231152 229284 231180
rect 101548 231140 101554 231152
rect 229278 231140 229284 231152
rect 229336 231140 229342 231192
rect 134518 231072 134524 231124
rect 134576 231112 134582 231124
rect 442994 231112 443000 231124
rect 134576 231084 443000 231112
rect 134576 231072 134582 231084
rect 442994 231072 443000 231084
rect 443052 231072 443058 231124
rect 82906 230392 82912 230444
rect 82964 230432 82970 230444
rect 83458 230432 83464 230444
rect 82964 230404 83464 230432
rect 82964 230392 82970 230404
rect 83458 230392 83464 230404
rect 83516 230432 83522 230444
rect 149054 230432 149060 230444
rect 83516 230404 149060 230432
rect 83516 230392 83522 230404
rect 149054 230392 149060 230404
rect 149112 230392 149118 230444
rect 89254 230324 89260 230376
rect 89312 230364 89318 230376
rect 126974 230364 126980 230376
rect 89312 230336 126980 230364
rect 89312 230324 89318 230336
rect 126974 230324 126980 230336
rect 127032 230364 127038 230376
rect 127434 230364 127440 230376
rect 127032 230336 127440 230364
rect 127032 230324 127038 230336
rect 127434 230324 127440 230336
rect 127492 230324 127498 230376
rect 67450 229848 67456 229900
rect 67508 229888 67514 229900
rect 230474 229888 230480 229900
rect 67508 229860 230480 229888
rect 67508 229848 67514 229860
rect 230474 229848 230480 229860
rect 230532 229848 230538 229900
rect 127434 229780 127440 229832
rect 127492 229820 127498 229832
rect 173158 229820 173164 229832
rect 127492 229792 173164 229820
rect 127492 229780 127498 229792
rect 173158 229780 173164 229792
rect 173216 229780 173222 229832
rect 180058 229780 180064 229832
rect 180116 229820 180122 229832
rect 382274 229820 382280 229832
rect 180116 229792 382280 229820
rect 180116 229780 180122 229792
rect 382274 229780 382280 229792
rect 382332 229780 382338 229832
rect 48222 229712 48228 229764
rect 48280 229752 48286 229764
rect 276842 229752 276848 229764
rect 48280 229724 276848 229752
rect 48280 229712 48286 229724
rect 276842 229712 276848 229724
rect 276900 229712 276906 229764
rect 111886 228420 111892 228472
rect 111944 228460 111950 228472
rect 378134 228460 378140 228472
rect 111944 228432 378140 228460
rect 111944 228420 111950 228432
rect 378134 228420 378140 228432
rect 378192 228420 378198 228472
rect 98638 228352 98644 228404
rect 98696 228392 98702 228404
rect 418890 228392 418896 228404
rect 98696 228364 418896 228392
rect 98696 228352 98702 228364
rect 418890 228352 418896 228364
rect 418948 228352 418954 228404
rect 94038 226992 94044 227044
rect 94096 227032 94102 227044
rect 235994 227032 236000 227044
rect 94096 227004 236000 227032
rect 94096 226992 94102 227004
rect 235994 226992 236000 227004
rect 236052 226992 236058 227044
rect 60550 225700 60556 225752
rect 60608 225740 60614 225752
rect 164878 225740 164884 225752
rect 60608 225712 164884 225740
rect 60608 225700 60614 225712
rect 164878 225700 164884 225712
rect 164936 225700 164942 225752
rect 56318 225632 56324 225684
rect 56376 225672 56382 225684
rect 252554 225672 252560 225684
rect 56376 225644 252560 225672
rect 56376 225632 56382 225644
rect 252554 225632 252560 225644
rect 252612 225632 252618 225684
rect 74718 225564 74724 225616
rect 74776 225604 74782 225616
rect 303706 225604 303712 225616
rect 74776 225576 303712 225604
rect 74776 225564 74782 225576
rect 303706 225564 303712 225576
rect 303764 225564 303770 225616
rect 91738 224884 91744 224936
rect 91796 224924 91802 224936
rect 438946 224924 438952 224936
rect 91796 224896 438952 224924
rect 91796 224884 91802 224896
rect 438946 224884 438952 224896
rect 439004 224884 439010 224936
rect 438946 224476 438952 224528
rect 439004 224516 439010 224528
rect 439498 224516 439504 224528
rect 439004 224488 439504 224516
rect 439004 224476 439010 224488
rect 439498 224476 439504 224488
rect 439556 224476 439562 224528
rect 59170 224272 59176 224324
rect 59228 224312 59234 224324
rect 187050 224312 187056 224324
rect 59228 224284 187056 224312
rect 59228 224272 59234 224284
rect 187050 224272 187056 224284
rect 187108 224272 187114 224324
rect 65978 224204 65984 224256
rect 66036 224244 66042 224256
rect 230566 224244 230572 224256
rect 66036 224216 230572 224244
rect 66036 224204 66042 224216
rect 230566 224204 230572 224216
rect 230624 224204 230630 224256
rect 59078 222844 59084 222896
rect 59136 222884 59142 222896
rect 417418 222884 417424 222896
rect 59136 222856 417424 222884
rect 59136 222844 59142 222856
rect 417418 222844 417424 222856
rect 417476 222844 417482 222896
rect 82906 222640 82912 222692
rect 82964 222680 82970 222692
rect 83458 222680 83464 222692
rect 82964 222652 83464 222680
rect 82964 222640 82970 222652
rect 83458 222640 83464 222652
rect 83516 222640 83522 222692
rect 4798 222164 4804 222216
rect 4856 222204 4862 222216
rect 82906 222204 82912 222216
rect 4856 222176 82912 222204
rect 4856 222164 4862 222176
rect 82906 222164 82912 222176
rect 82964 222164 82970 222216
rect 118234 222096 118240 222148
rect 118292 222136 118298 222148
rect 146294 222136 146300 222148
rect 118292 222108 146300 222136
rect 118292 222096 118298 222108
rect 146294 222096 146300 222108
rect 146352 222136 146358 222148
rect 146754 222136 146760 222148
rect 146352 222108 146760 222136
rect 146352 222096 146358 222108
rect 146754 222096 146760 222108
rect 146812 222096 146818 222148
rect 282270 221552 282276 221604
rect 282328 221592 282334 221604
rect 299474 221592 299480 221604
rect 282328 221564 299480 221592
rect 282328 221552 282334 221564
rect 299474 221552 299480 221564
rect 299532 221552 299538 221604
rect 146754 221484 146760 221536
rect 146812 221524 146818 221536
rect 301498 221524 301504 221536
rect 146812 221496 301504 221524
rect 146812 221484 146818 221496
rect 301498 221484 301504 221496
rect 301556 221484 301562 221536
rect 86310 221416 86316 221468
rect 86368 221456 86374 221468
rect 440234 221456 440240 221468
rect 86368 221428 440240 221456
rect 86368 221416 86374 221428
rect 440234 221416 440240 221428
rect 440292 221416 440298 221468
rect 233878 220124 233884 220176
rect 233936 220164 233942 220176
rect 309134 220164 309140 220176
rect 233936 220136 309140 220164
rect 233936 220124 233942 220136
rect 309134 220124 309140 220136
rect 309192 220124 309198 220176
rect 48038 220056 48044 220108
rect 48096 220096 48102 220108
rect 260190 220096 260196 220108
rect 48096 220068 260196 220096
rect 48096 220056 48102 220068
rect 260190 220056 260196 220068
rect 260248 220056 260254 220108
rect 89806 218764 89812 218816
rect 89864 218804 89870 218816
rect 233418 218804 233424 218816
rect 89864 218776 233424 218804
rect 89864 218764 89870 218776
rect 233418 218764 233424 218776
rect 233476 218764 233482 218816
rect 61378 218696 61384 218748
rect 61436 218736 61442 218748
rect 363598 218736 363604 218748
rect 61436 218708 363604 218736
rect 61436 218696 61442 218708
rect 363598 218696 363604 218708
rect 363656 218696 363662 218748
rect 446398 218696 446404 218748
rect 446456 218736 446462 218748
rect 580166 218736 580172 218748
rect 446456 218708 580172 218736
rect 446456 218696 446462 218708
rect 580166 218696 580172 218708
rect 580224 218696 580230 218748
rect 74626 217404 74632 217456
rect 74684 217444 74690 217456
rect 147674 217444 147680 217456
rect 74684 217416 147680 217444
rect 74684 217404 74690 217416
rect 147674 217404 147680 217416
rect 147732 217404 147738 217456
rect 41230 217336 41236 217388
rect 41288 217376 41294 217388
rect 275278 217376 275284 217388
rect 41288 217348 275284 217376
rect 41288 217336 41294 217348
rect 275278 217336 275284 217348
rect 275336 217336 275342 217388
rect 104158 217268 104164 217320
rect 104216 217308 104222 217320
rect 400214 217308 400220 217320
rect 104216 217280 400220 217308
rect 104216 217268 104222 217280
rect 400214 217268 400220 217280
rect 400272 217268 400278 217320
rect 54846 215908 54852 215960
rect 54904 215948 54910 215960
rect 414014 215948 414020 215960
rect 54904 215920 414020 215948
rect 54904 215908 54910 215920
rect 414014 215908 414020 215920
rect 414072 215908 414078 215960
rect 81526 215228 81532 215280
rect 81584 215268 81590 215280
rect 151814 215268 151820 215280
rect 81584 215240 151820 215268
rect 81584 215228 81590 215240
rect 151814 215228 151820 215240
rect 151872 215268 151878 215280
rect 153102 215268 153108 215280
rect 151872 215240 153108 215268
rect 151872 215228 151878 215240
rect 153102 215228 153108 215240
rect 153160 215228 153166 215280
rect 3326 214616 3332 214668
rect 3384 214656 3390 214668
rect 7558 214656 7564 214668
rect 3384 214628 7564 214656
rect 3384 214616 3390 214628
rect 7558 214616 7564 214628
rect 7616 214656 7622 214668
rect 209038 214656 209044 214668
rect 7616 214628 209044 214656
rect 7616 214616 7622 214628
rect 209038 214616 209044 214628
rect 209096 214616 209102 214668
rect 153102 214548 153108 214600
rect 153160 214588 153166 214600
rect 407114 214588 407120 214600
rect 153160 214560 407120 214588
rect 153160 214548 153166 214560
rect 407114 214548 407120 214560
rect 407172 214548 407178 214600
rect 69014 213188 69020 213240
rect 69072 213228 69078 213240
rect 391934 213228 391940 213240
rect 69072 213200 391940 213228
rect 69072 213188 69078 213200
rect 391934 213188 391940 213200
rect 391992 213188 391998 213240
rect 58618 211760 58624 211812
rect 58676 211800 58682 211812
rect 401594 211800 401600 211812
rect 58676 211772 401600 211800
rect 58676 211760 58682 211772
rect 401594 211760 401600 211772
rect 401652 211760 401658 211812
rect 45370 210400 45376 210452
rect 45428 210440 45434 210452
rect 307754 210440 307760 210452
rect 45428 210412 307760 210440
rect 45428 210400 45434 210412
rect 307754 210400 307760 210412
rect 307812 210400 307818 210452
rect 109678 209788 109684 209840
rect 109736 209828 109742 209840
rect 389174 209828 389180 209840
rect 109736 209800 389180 209828
rect 109736 209788 109742 209800
rect 389174 209788 389180 209800
rect 389232 209788 389238 209840
rect 113174 209108 113180 209160
rect 113232 209148 113238 209160
rect 302234 209148 302240 209160
rect 113232 209120 302240 209148
rect 113232 209108 113238 209120
rect 302234 209108 302240 209120
rect 302292 209108 302298 209160
rect 50890 209040 50896 209092
rect 50948 209080 50954 209092
rect 247034 209080 247040 209092
rect 50948 209052 247040 209080
rect 50948 209040 50954 209052
rect 247034 209040 247040 209052
rect 247092 209040 247098 209092
rect 111794 207680 111800 207732
rect 111852 207720 111858 207732
rect 249886 207720 249892 207732
rect 111852 207692 249892 207720
rect 111852 207680 111858 207692
rect 249886 207680 249892 207692
rect 249944 207680 249950 207732
rect 56410 207612 56416 207664
rect 56468 207652 56474 207664
rect 387794 207652 387800 207664
rect 56468 207624 387800 207652
rect 56468 207612 56474 207624
rect 387794 207612 387800 207624
rect 387852 207612 387858 207664
rect 100754 206320 100760 206372
rect 100812 206360 100818 206372
rect 225690 206360 225696 206372
rect 100812 206332 225696 206360
rect 100812 206320 100818 206332
rect 225690 206320 225696 206332
rect 225748 206320 225754 206372
rect 78766 206252 78772 206304
rect 78824 206292 78830 206304
rect 285674 206292 285680 206304
rect 78824 206264 285680 206292
rect 78824 206252 78830 206264
rect 285674 206252 285680 206264
rect 285732 206252 285738 206304
rect 450538 206252 450544 206304
rect 450596 206292 450602 206304
rect 580166 206292 580172 206304
rect 450596 206264 580172 206292
rect 450596 206252 450602 206264
rect 580166 206252 580172 206264
rect 580224 206252 580230 206304
rect 82814 205572 82820 205624
rect 82872 205612 82878 205624
rect 133874 205612 133880 205624
rect 82872 205584 133880 205612
rect 82872 205572 82878 205584
rect 133874 205572 133880 205584
rect 133932 205612 133938 205624
rect 135162 205612 135168 205624
rect 133932 205584 135168 205612
rect 133932 205572 133938 205584
rect 135162 205572 135168 205584
rect 135220 205572 135226 205624
rect 122098 205096 122104 205148
rect 122156 205136 122162 205148
rect 310606 205136 310612 205148
rect 122156 205108 310612 205136
rect 122156 205096 122162 205108
rect 310606 205096 310612 205108
rect 310664 205096 310670 205148
rect 55030 205028 55036 205080
rect 55088 205068 55094 205080
rect 248506 205068 248512 205080
rect 55088 205040 248512 205068
rect 55088 205028 55094 205040
rect 248506 205028 248512 205040
rect 248564 205028 248570 205080
rect 92566 204960 92572 205012
rect 92624 205000 92630 205012
rect 288434 205000 288440 205012
rect 92624 204972 288440 205000
rect 92624 204960 92630 204972
rect 288434 204960 288440 204972
rect 288492 204960 288498 205012
rect 135162 204892 135168 204944
rect 135220 204932 135226 204944
rect 429470 204932 429476 204944
rect 135220 204904 429476 204932
rect 135220 204892 135226 204904
rect 429470 204892 429476 204904
rect 429528 204892 429534 204944
rect 114462 203804 114468 203856
rect 114520 203844 114526 203856
rect 166350 203844 166356 203856
rect 114520 203816 166356 203844
rect 114520 203804 114526 203816
rect 166350 203804 166356 203816
rect 166408 203804 166414 203856
rect 86954 203736 86960 203788
rect 87012 203776 87018 203788
rect 251266 203776 251272 203788
rect 87012 203748 251272 203776
rect 87012 203736 87018 203748
rect 251266 203736 251272 203748
rect 251324 203736 251330 203788
rect 114554 203668 114560 203720
rect 114612 203708 114618 203720
rect 283190 203708 283196 203720
rect 114612 203680 283196 203708
rect 114612 203668 114618 203680
rect 283190 203668 283196 203680
rect 283248 203668 283254 203720
rect 63126 203600 63132 203652
rect 63184 203640 63190 203652
rect 299566 203640 299572 203652
rect 63184 203612 299572 203640
rect 63184 203600 63190 203612
rect 299566 203600 299572 203612
rect 299624 203600 299630 203652
rect 3326 203532 3332 203584
rect 3384 203572 3390 203584
rect 120074 203572 120080 203584
rect 3384 203544 120080 203572
rect 3384 203532 3390 203544
rect 120074 203532 120080 203544
rect 120132 203532 120138 203584
rect 164878 203532 164884 203584
rect 164936 203572 164942 203584
rect 439130 203572 439136 203584
rect 164936 203544 439136 203572
rect 164936 203532 164942 203544
rect 439130 203532 439136 203544
rect 439188 203532 439194 203584
rect 157978 202240 157984 202292
rect 158036 202280 158042 202292
rect 296714 202280 296720 202292
rect 158036 202252 296720 202280
rect 158036 202240 158042 202252
rect 296714 202240 296720 202252
rect 296772 202240 296778 202292
rect 86218 202172 86224 202224
rect 86276 202212 86282 202224
rect 242986 202212 242992 202224
rect 86276 202184 242992 202212
rect 86276 202172 86282 202184
rect 242986 202172 242992 202184
rect 243044 202172 243050 202224
rect 80146 202104 80152 202156
rect 80204 202144 80210 202156
rect 278222 202144 278228 202156
rect 80204 202116 278228 202144
rect 80204 202104 80210 202116
rect 278222 202104 278228 202116
rect 278280 202104 278286 202156
rect 228450 201084 228456 201136
rect 228508 201124 228514 201136
rect 298186 201124 298192 201136
rect 228508 201096 298192 201124
rect 228508 201084 228514 201096
rect 298186 201084 298192 201096
rect 298244 201084 298250 201136
rect 96706 201016 96712 201068
rect 96764 201056 96770 201068
rect 241606 201056 241612 201068
rect 96764 201028 241612 201056
rect 96764 201016 96770 201028
rect 241606 201016 241612 201028
rect 241664 201016 241670 201068
rect 104894 200948 104900 201000
rect 104952 200988 104958 201000
rect 272610 200988 272616 201000
rect 104952 200960 272616 200988
rect 104952 200948 104958 200960
rect 272610 200948 272616 200960
rect 272668 200948 272674 201000
rect 49510 200880 49516 200932
rect 49568 200920 49574 200932
rect 237374 200920 237380 200932
rect 49568 200892 237380 200920
rect 49568 200880 49574 200892
rect 237374 200880 237380 200892
rect 237432 200880 237438 200932
rect 67358 200812 67364 200864
rect 67416 200852 67422 200864
rect 307938 200852 307944 200864
rect 67416 200824 307944 200852
rect 67416 200812 67422 200824
rect 307938 200812 307944 200824
rect 307996 200812 308002 200864
rect 99190 200744 99196 200796
rect 99248 200784 99254 200796
rect 443086 200784 443092 200796
rect 99248 200756 443092 200784
rect 99248 200744 99254 200756
rect 443086 200744 443092 200756
rect 443144 200744 443150 200796
rect 144178 199520 144184 199572
rect 144236 199560 144242 199572
rect 223022 199560 223028 199572
rect 144236 199532 223028 199560
rect 144236 199520 144242 199532
rect 223022 199520 223028 199532
rect 223080 199520 223086 199572
rect 116026 199452 116032 199504
rect 116084 199492 116090 199504
rect 428090 199492 428096 199504
rect 116084 199464 428096 199492
rect 116084 199452 116090 199464
rect 428090 199452 428096 199464
rect 428148 199452 428154 199504
rect 82078 199384 82084 199436
rect 82136 199424 82142 199436
rect 432230 199424 432236 199436
rect 82136 199396 432236 199424
rect 82136 199384 82142 199396
rect 432230 199384 432236 199396
rect 432288 199384 432294 199436
rect 50798 198092 50804 198144
rect 50856 198132 50862 198144
rect 217318 198132 217324 198144
rect 50856 198104 217324 198132
rect 50856 198092 50862 198104
rect 217318 198092 217324 198104
rect 217376 198092 217382 198144
rect 280890 198092 280896 198144
rect 280948 198132 280954 198144
rect 301038 198132 301044 198144
rect 280948 198104 301044 198132
rect 280948 198092 280954 198104
rect 301038 198092 301044 198104
rect 301096 198092 301102 198144
rect 93946 198024 93952 198076
rect 94004 198064 94010 198076
rect 305086 198064 305092 198076
rect 94004 198036 305092 198064
rect 94004 198024 94010 198036
rect 305086 198024 305092 198036
rect 305144 198024 305150 198076
rect 61838 197956 61844 198008
rect 61896 197996 61902 198008
rect 302326 197996 302332 198008
rect 61896 197968 302332 197996
rect 61896 197956 61902 197968
rect 302326 197956 302332 197968
rect 302384 197956 302390 198008
rect 110414 196800 110420 196852
rect 110472 196840 110478 196852
rect 233326 196840 233332 196852
rect 110472 196812 233332 196840
rect 110472 196800 110478 196812
rect 233326 196800 233332 196812
rect 233384 196800 233390 196852
rect 105538 196732 105544 196784
rect 105596 196772 105602 196784
rect 240226 196772 240232 196784
rect 105596 196744 240232 196772
rect 105596 196732 105602 196744
rect 240226 196732 240232 196744
rect 240284 196732 240290 196784
rect 65886 196664 65892 196716
rect 65944 196704 65950 196716
rect 295426 196704 295432 196716
rect 65944 196676 295432 196704
rect 65944 196664 65950 196676
rect 295426 196664 295432 196676
rect 295484 196664 295490 196716
rect 83458 196596 83464 196648
rect 83516 196636 83522 196648
rect 369854 196636 369860 196648
rect 83516 196608 369860 196636
rect 83516 196596 83522 196608
rect 369854 196596 369860 196608
rect 369912 196596 369918 196648
rect 92474 195440 92480 195492
rect 92532 195480 92538 195492
rect 211890 195480 211896 195492
rect 92532 195452 211896 195480
rect 92532 195440 92538 195452
rect 211890 195440 211896 195452
rect 211948 195440 211954 195492
rect 222838 195440 222844 195492
rect 222896 195480 222902 195492
rect 294046 195480 294052 195492
rect 222896 195452 294052 195480
rect 222896 195440 222902 195452
rect 294046 195440 294052 195452
rect 294104 195440 294110 195492
rect 209130 195372 209136 195424
rect 209188 195412 209194 195424
rect 437566 195412 437572 195424
rect 209188 195384 437572 195412
rect 209188 195372 209194 195384
rect 437566 195372 437572 195384
rect 437624 195372 437630 195424
rect 49418 195304 49424 195356
rect 49476 195344 49482 195356
rect 306466 195344 306472 195356
rect 49476 195316 306472 195344
rect 49476 195304 49482 195316
rect 306466 195304 306472 195316
rect 306524 195304 306530 195356
rect 59262 195236 59268 195288
rect 59320 195276 59326 195288
rect 436094 195276 436100 195288
rect 59320 195248 436100 195276
rect 59320 195236 59326 195248
rect 436094 195236 436100 195248
rect 436152 195236 436158 195288
rect 89714 194148 89720 194200
rect 89772 194188 89778 194200
rect 252646 194188 252652 194200
rect 89772 194160 252652 194188
rect 89772 194148 89778 194160
rect 252646 194148 252652 194160
rect 252704 194148 252710 194200
rect 64598 194080 64604 194132
rect 64656 194120 64662 194132
rect 230658 194120 230664 194132
rect 64656 194092 230664 194120
rect 64656 194080 64662 194092
rect 230658 194080 230664 194092
rect 230716 194080 230722 194132
rect 93854 194012 93860 194064
rect 93912 194052 93918 194064
rect 309226 194052 309232 194064
rect 93912 194024 309232 194052
rect 93912 194012 93918 194024
rect 309226 194012 309232 194024
rect 309284 194012 309290 194064
rect 60642 193944 60648 193996
rect 60700 193984 60706 193996
rect 278314 193984 278320 193996
rect 60700 193956 278320 193984
rect 60700 193944 60706 193956
rect 278314 193944 278320 193956
rect 278372 193944 278378 193996
rect 99282 193876 99288 193928
rect 99340 193916 99346 193928
rect 329098 193916 329104 193928
rect 99340 193888 329104 193916
rect 99340 193876 99346 193888
rect 329098 193876 329104 193888
rect 329156 193876 329162 193928
rect 155218 193808 155224 193860
rect 155276 193848 155282 193860
rect 447134 193848 447140 193860
rect 155276 193820 447140 193848
rect 155276 193808 155282 193820
rect 447134 193808 447140 193820
rect 447192 193808 447198 193860
rect 53558 192584 53564 192636
rect 53616 192624 53622 192636
rect 221642 192624 221648 192636
rect 53616 192596 221648 192624
rect 53616 192584 53622 192596
rect 221642 192584 221648 192596
rect 221700 192584 221706 192636
rect 160738 192516 160744 192568
rect 160796 192556 160802 192568
rect 434806 192556 434812 192568
rect 160796 192528 434812 192556
rect 160796 192516 160802 192528
rect 434806 192516 434812 192528
rect 434864 192516 434870 192568
rect 60458 192448 60464 192500
rect 60516 192488 60522 192500
rect 451274 192488 451280 192500
rect 60516 192460 451280 192488
rect 60516 192448 60522 192460
rect 451274 192448 451280 192460
rect 451332 192448 451338 192500
rect 475378 192448 475384 192500
rect 475436 192488 475442 192500
rect 579614 192488 579620 192500
rect 475436 192460 579620 192488
rect 475436 192448 475442 192460
rect 579614 192448 579620 192460
rect 579672 192448 579678 192500
rect 203518 191360 203524 191412
rect 203576 191400 203582 191412
rect 244274 191400 244280 191412
rect 203576 191372 244280 191400
rect 203576 191360 203582 191372
rect 244274 191360 244280 191372
rect 244332 191360 244338 191412
rect 244918 191360 244924 191412
rect 244976 191400 244982 191412
rect 337470 191400 337476 191412
rect 244976 191372 337476 191400
rect 244976 191360 244982 191372
rect 337470 191360 337476 191372
rect 337528 191360 337534 191412
rect 102134 191292 102140 191344
rect 102192 191332 102198 191344
rect 292666 191332 292672 191344
rect 102192 191304 292672 191332
rect 102192 191292 102198 191304
rect 292666 191292 292672 191304
rect 292724 191292 292730 191344
rect 66070 191224 66076 191276
rect 66128 191264 66134 191276
rect 256786 191264 256792 191276
rect 66128 191236 256792 191264
rect 66128 191224 66134 191236
rect 256786 191224 256792 191236
rect 256844 191224 256850 191276
rect 50982 191156 50988 191208
rect 51040 191196 51046 191208
rect 245746 191196 245752 191208
rect 51040 191168 245752 191196
rect 51040 191156 51046 191168
rect 245746 191156 245752 191168
rect 245804 191156 245810 191208
rect 88334 191088 88340 191140
rect 88392 191128 88398 191140
rect 285950 191128 285956 191140
rect 88392 191100 285956 191128
rect 88392 191088 88398 191100
rect 285950 191088 285956 191100
rect 286008 191088 286014 191140
rect 108942 190476 108948 190528
rect 109000 190516 109006 190528
rect 214742 190516 214748 190528
rect 109000 190488 214748 190516
rect 109000 190476 109006 190488
rect 214742 190476 214748 190488
rect 214800 190476 214806 190528
rect 77294 189864 77300 189916
rect 77352 189904 77358 189916
rect 229186 189904 229192 189916
rect 77352 189876 229192 189904
rect 77352 189864 77358 189876
rect 229186 189864 229192 189876
rect 229244 189864 229250 189916
rect 73246 189796 73252 189848
rect 73304 189836 73310 189848
rect 285858 189836 285864 189848
rect 73304 189808 285864 189836
rect 73304 189796 73310 189808
rect 285858 189796 285864 189808
rect 285916 189796 285922 189848
rect 169018 189728 169024 189780
rect 169076 189768 169082 189780
rect 436370 189768 436376 189780
rect 169076 189740 436376 189768
rect 169076 189728 169082 189740
rect 436370 189728 436376 189740
rect 436428 189728 436434 189780
rect 106182 189184 106188 189236
rect 106240 189224 106246 189236
rect 169110 189224 169116 189236
rect 106240 189196 169116 189224
rect 106240 189184 106246 189196
rect 169110 189184 169116 189196
rect 169168 189184 169174 189236
rect 104802 189116 104808 189168
rect 104860 189156 104866 189168
rect 173250 189156 173256 189168
rect 104860 189128 173256 189156
rect 104860 189116 104866 189128
rect 173250 189116 173256 189128
rect 173308 189116 173314 189168
rect 3510 189048 3516 189100
rect 3568 189088 3574 189100
rect 4062 189088 4068 189100
rect 3568 189060 4068 189088
rect 3568 189048 3574 189060
rect 4062 189048 4068 189060
rect 4120 189088 4126 189100
rect 441706 189088 441712 189100
rect 4120 189060 441712 189088
rect 4120 189048 4126 189060
rect 441706 189048 441712 189060
rect 441764 189048 441770 189100
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 11698 189020 11704 189032
rect 3476 188992 11704 189020
rect 3476 188980 3482 188992
rect 11698 188980 11704 188992
rect 11756 188980 11762 189032
rect 279510 188640 279516 188692
rect 279568 188680 279574 188692
rect 292758 188680 292764 188692
rect 279568 188652 292764 188680
rect 279568 188640 279574 188652
rect 292758 188640 292764 188652
rect 292816 188640 292822 188692
rect 278130 188572 278136 188624
rect 278188 188612 278194 188624
rect 306558 188612 306564 188624
rect 278188 188584 306564 188612
rect 278188 188572 278194 188584
rect 306558 188572 306564 188584
rect 306616 188572 306622 188624
rect 99374 188504 99380 188556
rect 99432 188544 99438 188556
rect 280338 188544 280344 188556
rect 99432 188516 280344 188544
rect 99432 188504 99438 188516
rect 280338 188504 280344 188516
rect 280396 188504 280402 188556
rect 118694 188436 118700 188488
rect 118752 188476 118758 188488
rect 309318 188476 309324 188488
rect 118752 188448 309324 188476
rect 118752 188436 118758 188448
rect 309318 188436 309324 188448
rect 309376 188436 309382 188488
rect 71774 188368 71780 188420
rect 71832 188408 71838 188420
rect 280154 188408 280160 188420
rect 71832 188380 280160 188408
rect 71832 188368 71838 188380
rect 280154 188368 280160 188380
rect 280212 188368 280218 188420
rect 54938 188300 54944 188352
rect 54996 188340 55002 188352
rect 305178 188340 305184 188352
rect 54996 188312 305184 188340
rect 54996 188300 55002 188312
rect 305178 188300 305184 188312
rect 305236 188300 305242 188352
rect 103422 187756 103428 187808
rect 103480 187796 103486 187808
rect 171778 187796 171784 187808
rect 103480 187768 171784 187796
rect 103480 187756 103486 187768
rect 171778 187756 171784 187768
rect 171836 187756 171842 187808
rect 131022 187688 131028 187740
rect 131080 187728 131086 187740
rect 209130 187728 209136 187740
rect 131080 187700 209136 187728
rect 131080 187688 131086 187700
rect 209130 187688 209136 187700
rect 209188 187688 209194 187740
rect 146938 187076 146944 187128
rect 146996 187116 147002 187128
rect 175918 187116 175924 187128
rect 146996 187088 175924 187116
rect 146996 187076 147002 187088
rect 175918 187076 175924 187088
rect 175976 187076 175982 187128
rect 95234 187008 95240 187060
rect 95292 187048 95298 187060
rect 274082 187048 274088 187060
rect 95292 187020 274088 187048
rect 95292 187008 95298 187020
rect 274082 187008 274088 187020
rect 274140 187008 274146 187060
rect 73154 186940 73160 186992
rect 73212 186980 73218 186992
rect 291286 186980 291292 186992
rect 73212 186952 291292 186980
rect 73212 186940 73218 186952
rect 291286 186940 291292 186952
rect 291344 186940 291350 186992
rect 348970 186940 348976 186992
rect 349028 186980 349034 186992
rect 580902 186980 580908 186992
rect 349028 186952 580908 186980
rect 349028 186940 349034 186952
rect 580902 186940 580908 186952
rect 580960 186940 580966 186992
rect 153838 185852 153844 185904
rect 153896 185892 153902 185904
rect 289906 185892 289912 185904
rect 153896 185864 289912 185892
rect 153896 185852 153902 185864
rect 289906 185852 289912 185864
rect 289964 185852 289970 185904
rect 84194 185784 84200 185836
rect 84252 185824 84258 185836
rect 280246 185824 280252 185836
rect 84252 185796 280252 185824
rect 84252 185784 84258 185796
rect 280246 185784 280252 185796
rect 280304 185784 280310 185836
rect 52270 185716 52276 185768
rect 52328 185756 52334 185768
rect 251358 185756 251364 185768
rect 52328 185728 251364 185756
rect 52328 185716 52334 185728
rect 251358 185716 251364 185728
rect 251416 185716 251422 185768
rect 264238 185716 264244 185768
rect 264296 185756 264302 185768
rect 448606 185756 448612 185768
rect 264296 185728 448612 185756
rect 264296 185716 264302 185728
rect 448606 185716 448612 185728
rect 448664 185716 448670 185768
rect 80054 185648 80060 185700
rect 80112 185688 80118 185700
rect 310698 185688 310704 185700
rect 80112 185660 310704 185688
rect 80112 185648 80118 185660
rect 310698 185648 310704 185660
rect 310756 185648 310762 185700
rect 39942 185580 39948 185632
rect 40000 185620 40006 185632
rect 295518 185620 295524 185632
rect 40000 185592 295524 185620
rect 40000 185580 40006 185592
rect 295518 185580 295524 185592
rect 295576 185580 295582 185632
rect 350810 185580 350816 185632
rect 350868 185620 350874 185632
rect 381538 185620 381544 185632
rect 350868 185592 381544 185620
rect 350868 185580 350874 185592
rect 381538 185580 381544 185592
rect 381596 185580 381602 185632
rect 395338 185580 395344 185632
rect 395396 185620 395402 185632
rect 425790 185620 425796 185632
rect 395396 185592 425796 185620
rect 395396 185580 395402 185592
rect 425790 185580 425796 185592
rect 425848 185580 425854 185632
rect 100662 184900 100668 184952
rect 100720 184940 100726 184952
rect 169202 184940 169208 184952
rect 100720 184912 169208 184940
rect 100720 184900 100726 184912
rect 169202 184900 169208 184912
rect 169260 184900 169266 184952
rect 151078 184424 151084 184476
rect 151136 184464 151142 184476
rect 174538 184464 174544 184476
rect 151136 184436 174544 184464
rect 151136 184424 151142 184436
rect 174538 184424 174544 184436
rect 174596 184424 174602 184476
rect 210418 184424 210424 184476
rect 210476 184464 210482 184476
rect 243078 184464 243084 184476
rect 210476 184436 243084 184464
rect 210476 184424 210482 184436
rect 243078 184424 243084 184436
rect 243136 184424 243142 184476
rect 103698 184356 103704 184408
rect 103756 184396 103762 184408
rect 284478 184396 284484 184408
rect 103756 184368 284484 184396
rect 103756 184356 103762 184368
rect 284478 184356 284484 184368
rect 284536 184356 284542 184408
rect 63218 184288 63224 184340
rect 63276 184328 63282 184340
rect 247126 184328 247132 184340
rect 63276 184300 247132 184328
rect 63276 184288 63282 184300
rect 247126 184288 247132 184300
rect 247184 184288 247190 184340
rect 271138 184288 271144 184340
rect 271196 184328 271202 184340
rect 445846 184328 445852 184340
rect 271196 184300 445852 184328
rect 271196 184288 271202 184300
rect 445846 184288 445852 184300
rect 445904 184288 445910 184340
rect 75914 184220 75920 184272
rect 75972 184260 75978 184272
rect 285766 184260 285772 184272
rect 75972 184232 285772 184260
rect 75972 184220 75978 184232
rect 285766 184220 285772 184232
rect 285824 184220 285830 184272
rect 44082 184152 44088 184204
rect 44140 184192 44146 184204
rect 291194 184192 291200 184204
rect 44140 184164 291200 184192
rect 44140 184152 44146 184164
rect 291194 184152 291200 184164
rect 291252 184152 291258 184204
rect 358078 184152 358084 184204
rect 358136 184192 358142 184204
rect 374638 184192 374644 184204
rect 358136 184164 374644 184192
rect 358136 184152 358142 184164
rect 374638 184152 374644 184164
rect 374696 184152 374702 184204
rect 129642 183540 129648 183592
rect 129700 183580 129706 183592
rect 209314 183580 209320 183592
rect 129700 183552 209320 183580
rect 129700 183540 129706 183552
rect 209314 183540 209320 183552
rect 209372 183540 209378 183592
rect 187050 183064 187056 183116
rect 187108 183104 187114 183116
rect 244366 183104 244372 183116
rect 187108 183076 244372 183104
rect 187108 183064 187114 183076
rect 244366 183064 244372 183076
rect 244424 183064 244430 183116
rect 255958 183064 255964 183116
rect 256016 183104 256022 183116
rect 296898 183104 296904 183116
rect 256016 183076 296904 183104
rect 256016 183064 256022 183076
rect 296898 183064 296904 183076
rect 296956 183064 296962 183116
rect 142798 182996 142804 183048
rect 142856 183036 142862 183048
rect 238754 183036 238760 183048
rect 142856 183008 238760 183036
rect 142856 182996 142862 183008
rect 238754 182996 238760 183008
rect 238812 182996 238818 183048
rect 265618 182996 265624 183048
rect 265676 183036 265682 183048
rect 316862 183036 316868 183048
rect 265676 183008 316868 183036
rect 265676 182996 265682 183008
rect 316862 182996 316868 183008
rect 316920 182996 316926 183048
rect 411898 182996 411904 183048
rect 411956 183036 411962 183048
rect 443178 183036 443184 183048
rect 411956 183008 443184 183036
rect 411956 182996 411962 183008
rect 443178 182996 443184 183008
rect 443236 182996 443242 183048
rect 115934 182928 115940 182980
rect 115992 182968 115998 182980
rect 241698 182968 241704 182980
rect 115992 182940 241704 182968
rect 115992 182928 115998 182940
rect 241698 182928 241704 182940
rect 241756 182928 241762 182980
rect 262950 182928 262956 182980
rect 263008 182968 263014 182980
rect 319438 182968 319444 182980
rect 263008 182940 319444 182968
rect 263008 182928 263014 182940
rect 319438 182928 319444 182940
rect 319496 182928 319502 182980
rect 400858 182928 400864 182980
rect 400916 182968 400922 182980
rect 449894 182968 449900 182980
rect 400916 182940 449900 182968
rect 400916 182928 400922 182940
rect 449894 182928 449900 182940
rect 449952 182928 449958 182980
rect 64690 182860 64696 182912
rect 64748 182900 64754 182912
rect 230750 182900 230756 182912
rect 64748 182872 230756 182900
rect 64748 182860 64754 182872
rect 230750 182860 230756 182872
rect 230808 182860 230814 182912
rect 269758 182860 269764 182912
rect 269816 182900 269822 182912
rect 434898 182900 434904 182912
rect 269816 182872 434904 182900
rect 269816 182860 269822 182872
rect 434898 182860 434904 182872
rect 434956 182860 434962 182912
rect 107654 182792 107660 182844
rect 107712 182832 107718 182844
rect 307846 182832 307852 182844
rect 107712 182804 307852 182832
rect 107712 182792 107718 182804
rect 307846 182792 307852 182804
rect 307904 182792 307910 182844
rect 360838 182792 360844 182844
rect 360896 182832 360902 182844
rect 444466 182832 444472 182844
rect 360896 182804 444472 182832
rect 360896 182792 360902 182804
rect 444466 182792 444472 182804
rect 444524 182792 444530 182844
rect 119522 182180 119528 182232
rect 119580 182220 119586 182232
rect 211798 182220 211804 182232
rect 119580 182192 211804 182220
rect 119580 182180 119586 182192
rect 211798 182180 211804 182192
rect 211856 182180 211862 182232
rect 220262 181772 220268 181824
rect 220320 181812 220326 181824
rect 237466 181812 237472 181824
rect 220320 181784 237472 181812
rect 220320 181772 220326 181784
rect 237466 181772 237472 181784
rect 237524 181772 237530 181824
rect 269850 181772 269856 181824
rect 269908 181812 269914 181824
rect 314102 181812 314108 181824
rect 269908 181784 314108 181812
rect 269908 181772 269914 181784
rect 314102 181772 314108 181784
rect 314160 181772 314166 181824
rect 162118 181704 162124 181756
rect 162176 181744 162182 181756
rect 200758 181744 200764 181756
rect 162176 181716 200764 181744
rect 162176 181704 162182 181716
rect 200758 181704 200764 181716
rect 200816 181704 200822 181756
rect 200850 181704 200856 181756
rect 200908 181744 200914 181756
rect 240318 181744 240324 181756
rect 200908 181716 240324 181744
rect 200908 181704 200914 181716
rect 240318 181704 240324 181716
rect 240376 181704 240382 181756
rect 251818 181704 251824 181756
rect 251876 181744 251882 181756
rect 296806 181744 296812 181756
rect 251876 181716 296812 181744
rect 251876 181704 251882 181716
rect 296806 181704 296812 181716
rect 296864 181704 296870 181756
rect 199378 181636 199384 181688
rect 199436 181676 199442 181688
rect 248598 181676 248604 181688
rect 199436 181648 248604 181676
rect 199436 181636 199442 181648
rect 248598 181636 248604 181648
rect 248656 181636 248662 181688
rect 249058 181636 249064 181688
rect 249116 181676 249122 181688
rect 300210 181676 300216 181688
rect 249116 181648 300216 181676
rect 249116 181636 249122 181648
rect 300210 181636 300216 181648
rect 300268 181636 300274 181688
rect 167638 181568 167644 181620
rect 167696 181608 167702 181620
rect 244458 181608 244464 181620
rect 167696 181580 244464 181608
rect 167696 181568 167702 181580
rect 244458 181568 244464 181580
rect 244516 181568 244522 181620
rect 264330 181568 264336 181620
rect 264388 181608 264394 181620
rect 323670 181608 323676 181620
rect 264388 181580 323676 181608
rect 264388 181568 264394 181580
rect 323670 181568 323676 181580
rect 323728 181568 323734 181620
rect 96614 181500 96620 181552
rect 96672 181540 96678 181552
rect 202230 181540 202236 181552
rect 96672 181512 202236 181540
rect 96672 181500 96678 181512
rect 202230 181500 202236 181512
rect 202288 181500 202294 181552
rect 214650 181500 214656 181552
rect 214708 181540 214714 181552
rect 237558 181540 237564 181552
rect 214708 181512 237564 181540
rect 214708 181500 214714 181512
rect 237558 181500 237564 181512
rect 237616 181500 237622 181552
rect 245010 181500 245016 181552
rect 245068 181540 245074 181552
rect 424410 181540 424416 181552
rect 245068 181512 424416 181540
rect 245068 181500 245074 181512
rect 424410 181500 424416 181512
rect 424468 181500 424474 181552
rect 53742 181432 53748 181484
rect 53800 181472 53806 181484
rect 298278 181472 298284 181484
rect 53800 181444 298284 181472
rect 53800 181432 53806 181444
rect 298278 181432 298284 181444
rect 298336 181432 298342 181484
rect 361298 181432 361304 181484
rect 361356 181472 361362 181484
rect 405734 181472 405740 181484
rect 361356 181444 405740 181472
rect 361356 181432 361362 181444
rect 405734 181432 405740 181444
rect 405792 181432 405798 181484
rect 132402 180956 132408 181008
rect 132460 180996 132466 181008
rect 164878 180996 164884 181008
rect 132460 180968 164884 180996
rect 132460 180956 132466 180968
rect 164878 180956 164884 180968
rect 164936 180956 164942 181008
rect 122006 180888 122012 180940
rect 122064 180928 122070 180940
rect 167822 180928 167828 180940
rect 122064 180900 167828 180928
rect 122064 180888 122070 180900
rect 167822 180888 167828 180900
rect 167880 180888 167886 180940
rect 116946 180820 116952 180872
rect 117004 180860 117010 180872
rect 167730 180860 167736 180872
rect 117004 180832 167736 180860
rect 117004 180820 117010 180832
rect 167730 180820 167736 180832
rect 167788 180820 167794 180872
rect 223022 180412 223028 180464
rect 223080 180452 223086 180464
rect 236178 180452 236184 180464
rect 223080 180424 236184 180452
rect 223080 180412 223086 180424
rect 236178 180412 236184 180424
rect 236236 180412 236242 180464
rect 272518 180412 272524 180464
rect 272576 180452 272582 180464
rect 288618 180452 288624 180464
rect 272576 180424 288624 180452
rect 272576 180412 272582 180424
rect 288618 180412 288624 180424
rect 288676 180412 288682 180464
rect 222930 180344 222936 180396
rect 222988 180384 222994 180396
rect 236086 180384 236092 180396
rect 222988 180356 236092 180384
rect 222988 180344 222994 180356
rect 236086 180344 236092 180356
rect 236144 180344 236150 180396
rect 273898 180344 273904 180396
rect 273956 180384 273962 180396
rect 302418 180384 302424 180396
rect 273956 180356 302424 180384
rect 273956 180344 273962 180356
rect 302418 180344 302424 180356
rect 302476 180344 302482 180396
rect 225598 180276 225604 180328
rect 225656 180316 225662 180328
rect 245838 180316 245844 180328
rect 225656 180288 245844 180316
rect 225656 180276 225662 180288
rect 245838 180276 245844 180288
rect 245896 180276 245902 180328
rect 273990 180276 273996 180328
rect 274048 180316 274054 180328
rect 303798 180316 303804 180328
rect 274048 180288 303804 180316
rect 274048 180276 274054 180288
rect 303798 180276 303804 180288
rect 303856 180276 303862 180328
rect 414658 180276 414664 180328
rect 414716 180316 414722 180328
rect 444374 180316 444380 180328
rect 414716 180288 444380 180316
rect 414716 180276 414722 180288
rect 444374 180276 444380 180288
rect 444432 180276 444438 180328
rect 220170 180208 220176 180260
rect 220228 180248 220234 180260
rect 247218 180248 247224 180260
rect 220228 180220 247224 180248
rect 220228 180208 220234 180220
rect 247218 180208 247224 180220
rect 247276 180208 247282 180260
rect 258718 180208 258724 180260
rect 258776 180248 258782 180260
rect 294138 180248 294144 180260
rect 258776 180220 294144 180248
rect 258776 180208 258782 180220
rect 294138 180208 294144 180220
rect 294196 180208 294202 180260
rect 363782 180208 363788 180260
rect 363840 180248 363846 180260
rect 376754 180248 376760 180260
rect 363840 180220 376760 180248
rect 363840 180208 363846 180220
rect 376754 180208 376760 180220
rect 376812 180208 376818 180260
rect 407758 180208 407764 180260
rect 407816 180248 407822 180260
rect 439038 180248 439044 180260
rect 407816 180220 439044 180248
rect 407816 180208 407822 180220
rect 439038 180208 439044 180220
rect 439096 180208 439102 180260
rect 159358 180140 159364 180192
rect 159416 180180 159422 180192
rect 192478 180180 192484 180192
rect 159416 180152 192484 180180
rect 159416 180140 159422 180152
rect 192478 180140 192484 180152
rect 192536 180140 192542 180192
rect 198090 180140 198096 180192
rect 198148 180180 198154 180192
rect 347314 180180 347320 180192
rect 198148 180152 347320 180180
rect 198148 180140 198154 180152
rect 347314 180140 347320 180152
rect 347372 180140 347378 180192
rect 359458 180140 359464 180192
rect 359516 180180 359522 180192
rect 437474 180180 437480 180192
rect 359516 180152 437480 180180
rect 359516 180140 359522 180152
rect 437474 180140 437480 180152
rect 437532 180140 437538 180192
rect 173158 180072 173164 180124
rect 173216 180112 173222 180124
rect 438854 180112 438860 180124
rect 173216 180084 438860 180112
rect 173216 180072 173222 180084
rect 438854 180072 438860 180084
rect 438912 180072 438918 180124
rect 133138 179664 133144 179716
rect 133196 179704 133202 179716
rect 164418 179704 164424 179716
rect 133196 179676 164424 179704
rect 133196 179664 133202 179676
rect 164418 179664 164424 179676
rect 164476 179664 164482 179716
rect 120994 179596 121000 179648
rect 121052 179636 121058 179648
rect 166534 179636 166540 179648
rect 121052 179608 166540 179636
rect 121052 179596 121058 179608
rect 166534 179596 166540 179608
rect 166592 179596 166598 179648
rect 115842 179528 115848 179580
rect 115900 179568 115906 179580
rect 166442 179568 166448 179580
rect 115900 179540 166448 179568
rect 115900 179528 115906 179540
rect 166442 179528 166448 179540
rect 166500 179528 166506 179580
rect 97350 179460 97356 179512
rect 97408 179500 97414 179512
rect 173342 179500 173348 179512
rect 97408 179472 173348 179500
rect 97408 179460 97414 179472
rect 173342 179460 173348 179472
rect 173400 179460 173406 179512
rect 112254 179392 112260 179444
rect 112312 179432 112318 179444
rect 198182 179432 198188 179444
rect 112312 179404 198188 179432
rect 112312 179392 112318 179404
rect 198182 179392 198188 179404
rect 198240 179392 198246 179444
rect 276750 178984 276756 179036
rect 276808 179024 276814 179036
rect 289998 179024 290004 179036
rect 276808 178996 290004 179024
rect 276808 178984 276814 178996
rect 289998 178984 290004 178996
rect 290056 178984 290062 179036
rect 217318 178916 217324 178968
rect 217376 178956 217382 178968
rect 238938 178956 238944 178968
rect 217376 178928 238944 178956
rect 217376 178916 217382 178928
rect 238938 178916 238944 178928
rect 238996 178916 239002 178968
rect 272610 178916 272616 178968
rect 272668 178956 272674 178968
rect 287238 178956 287244 178968
rect 272668 178928 287244 178956
rect 272668 178916 272674 178928
rect 287238 178916 287244 178928
rect 287296 178916 287302 178968
rect 178770 178848 178776 178900
rect 178828 178888 178834 178900
rect 224954 178888 224960 178900
rect 178828 178860 224960 178888
rect 178828 178848 178834 178860
rect 224954 178848 224960 178860
rect 225012 178848 225018 178900
rect 257338 178848 257344 178900
rect 257396 178888 257402 178900
rect 295334 178888 295340 178900
rect 257396 178860 295340 178888
rect 257396 178848 257402 178860
rect 295334 178848 295340 178860
rect 295392 178848 295398 178900
rect 418798 178848 418804 178900
rect 418856 178888 418862 178900
rect 436186 178888 436192 178900
rect 418856 178860 436192 178888
rect 418856 178848 418862 178860
rect 436186 178848 436192 178860
rect 436244 178848 436250 178900
rect 214558 178780 214564 178832
rect 214616 178820 214622 178832
rect 312538 178820 312544 178832
rect 214616 178792 312544 178820
rect 214616 178780 214622 178792
rect 312538 178780 312544 178792
rect 312596 178780 312602 178832
rect 399478 178780 399484 178832
rect 399536 178820 399542 178832
rect 429378 178820 429384 178832
rect 399536 178792 429384 178820
rect 399536 178780 399542 178792
rect 429378 178780 429384 178792
rect 429436 178780 429442 178832
rect 64506 178712 64512 178764
rect 64564 178752 64570 178764
rect 254026 178752 254032 178764
rect 64564 178724 254032 178752
rect 64564 178712 64570 178724
rect 254026 178712 254032 178724
rect 254084 178712 254090 178764
rect 271230 178712 271236 178764
rect 271288 178752 271294 178764
rect 333330 178752 333336 178764
rect 271288 178724 333336 178752
rect 271288 178712 271294 178724
rect 333330 178712 333336 178724
rect 333388 178712 333394 178764
rect 358170 178712 358176 178764
rect 358228 178752 358234 178764
rect 433426 178752 433432 178764
rect 358228 178724 433432 178752
rect 358228 178712 358234 178724
rect 433426 178712 433432 178724
rect 433484 178712 433490 178764
rect 220078 178644 220084 178696
rect 220136 178684 220142 178696
rect 430574 178684 430580 178696
rect 220136 178656 430580 178684
rect 220136 178644 220142 178656
rect 430574 178644 430580 178656
rect 430632 178644 430638 178696
rect 148226 178304 148232 178356
rect 148284 178344 148290 178356
rect 169018 178344 169024 178356
rect 148284 178316 169024 178344
rect 148284 178304 148290 178316
rect 169018 178304 169024 178316
rect 169076 178304 169082 178356
rect 114370 178236 114376 178288
rect 114428 178276 114434 178288
rect 167914 178276 167920 178288
rect 114428 178248 167920 178276
rect 114428 178236 114434 178248
rect 167914 178236 167920 178248
rect 167972 178236 167978 178288
rect 109770 178168 109776 178220
rect 109828 178208 109834 178220
rect 170490 178208 170496 178220
rect 109828 178180 170496 178208
rect 109828 178168 109834 178180
rect 170490 178168 170496 178180
rect 170548 178168 170554 178220
rect 127066 178100 127072 178152
rect 127124 178140 127130 178152
rect 211982 178140 211988 178152
rect 127124 178112 211988 178140
rect 127124 178100 127130 178112
rect 211982 178100 211988 178112
rect 212040 178100 212046 178152
rect 214650 178072 214656 178084
rect 122806 178044 214656 178072
rect 118418 177964 118424 178016
rect 118476 178004 118482 178016
rect 122806 178004 122834 178044
rect 214650 178032 214656 178044
rect 214708 178032 214714 178084
rect 468478 178032 468484 178084
rect 468536 178072 468542 178084
rect 580166 178072 580172 178084
rect 468536 178044 580172 178072
rect 468536 178032 468542 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 118476 177976 122834 178004
rect 118476 177964 118482 177976
rect 278038 177624 278044 177676
rect 278096 177664 278102 177676
rect 288710 177664 288716 177676
rect 278096 177636 288716 177664
rect 278096 177624 278102 177636
rect 288710 177624 288716 177636
rect 288768 177624 288774 177676
rect 221642 177556 221648 177608
rect 221700 177596 221706 177608
rect 229554 177596 229560 177608
rect 221700 177568 229560 177596
rect 221700 177556 221706 177568
rect 229554 177556 229560 177568
rect 229612 177556 229618 177608
rect 275278 177556 275284 177608
rect 275336 177596 275342 177608
rect 294230 177596 294236 177608
rect 275336 177568 294236 177596
rect 275336 177556 275342 177568
rect 294230 177556 294236 177568
rect 294288 177556 294294 177608
rect 417418 177556 417424 177608
rect 417476 177596 417482 177608
rect 426894 177596 426900 177608
rect 417476 177568 426900 177596
rect 417476 177556 417482 177568
rect 426894 177556 426900 177568
rect 426952 177556 426958 177608
rect 227162 177488 227168 177540
rect 227220 177528 227226 177540
rect 234890 177528 234896 177540
rect 227220 177500 234896 177528
rect 227220 177488 227226 177500
rect 234890 177488 234896 177500
rect 234948 177488 234954 177540
rect 250438 177488 250444 177540
rect 250496 177528 250502 177540
rect 292574 177528 292580 177540
rect 250496 177500 292580 177528
rect 250496 177488 250502 177500
rect 292574 177488 292580 177500
rect 292632 177488 292638 177540
rect 413278 177488 413284 177540
rect 413336 177528 413342 177540
rect 434990 177528 434996 177540
rect 413336 177500 434996 177528
rect 413336 177488 413342 177500
rect 434990 177488 434996 177500
rect 435048 177488 435054 177540
rect 211890 177420 211896 177472
rect 211948 177460 211954 177472
rect 237650 177460 237656 177472
rect 211948 177432 237656 177460
rect 211948 177420 211954 177432
rect 237650 177420 237656 177432
rect 237708 177420 237714 177472
rect 268378 177420 268384 177472
rect 268436 177460 268442 177472
rect 325142 177460 325148 177472
rect 268436 177432 325148 177460
rect 268436 177420 268442 177432
rect 325142 177420 325148 177432
rect 325200 177420 325206 177472
rect 352558 177420 352564 177472
rect 352616 177460 352622 177472
rect 397454 177460 397460 177472
rect 352616 177432 397460 177460
rect 352616 177420 352622 177432
rect 397454 177420 397460 177432
rect 397512 177420 397518 177472
rect 418890 177420 418896 177472
rect 418948 177460 418954 177472
rect 441614 177460 441620 177472
rect 418948 177432 441620 177460
rect 418948 177420 418954 177432
rect 441614 177420 441620 177432
rect 441672 177420 441678 177472
rect 206370 177352 206376 177404
rect 206428 177392 206434 177404
rect 279418 177392 279424 177404
rect 206428 177364 279424 177392
rect 206428 177352 206434 177364
rect 279418 177352 279424 177364
rect 279476 177352 279482 177404
rect 363598 177352 363604 177404
rect 363656 177392 363662 177404
rect 422294 177392 422300 177404
rect 363656 177364 422300 177392
rect 363656 177352 363662 177364
rect 422294 177352 422300 177364
rect 422352 177352 422358 177404
rect 166350 177284 166356 177336
rect 166408 177324 166414 177336
rect 353294 177324 353300 177336
rect 166408 177296 353300 177324
rect 166408 177284 166414 177296
rect 353294 177284 353300 177296
rect 353352 177284 353358 177336
rect 370498 177284 370504 177336
rect 370556 177324 370562 177336
rect 437658 177324 437664 177336
rect 370556 177296 437664 177324
rect 370556 177284 370562 177296
rect 437658 177284 437664 177296
rect 437716 177284 437722 177336
rect 134426 176944 134432 176996
rect 134484 176984 134490 176996
rect 165246 176984 165252 176996
rect 134484 176956 165252 176984
rect 134484 176944 134490 176956
rect 165246 176944 165252 176956
rect 165304 176944 165310 176996
rect 125778 176876 125784 176928
rect 125836 176916 125842 176928
rect 166626 176916 166632 176928
rect 125836 176888 166632 176916
rect 125836 176876 125842 176888
rect 166626 176876 166632 176888
rect 166684 176876 166690 176928
rect 111058 176848 111064 176860
rect 109420 176820 111064 176848
rect 109420 176792 109448 176820
rect 111058 176808 111064 176820
rect 111116 176808 111122 176860
rect 124490 176808 124496 176860
rect 124548 176848 124554 176860
rect 170582 176848 170588 176860
rect 124548 176820 170588 176848
rect 124548 176808 124554 176820
rect 170582 176808 170588 176820
rect 170640 176808 170646 176860
rect 14458 176740 14464 176792
rect 14516 176780 14522 176792
rect 109402 176780 109408 176792
rect 14516 176752 109408 176780
rect 14516 176740 14522 176752
rect 109402 176740 109408 176752
rect 109460 176740 109466 176792
rect 110690 176740 110696 176792
rect 110748 176780 110754 176792
rect 214558 176780 214564 176792
rect 110748 176752 214564 176780
rect 110748 176740 110754 176752
rect 214558 176740 214564 176752
rect 214616 176740 214622 176792
rect 102042 176672 102048 176724
rect 102100 176712 102106 176724
rect 213362 176712 213368 176724
rect 102100 176684 213368 176712
rect 102100 176672 102106 176684
rect 213362 176672 213368 176684
rect 213420 176672 213426 176724
rect 240778 176672 240784 176724
rect 240836 176712 240842 176724
rect 241514 176712 241520 176724
rect 240836 176684 241520 176712
rect 240836 176672 240842 176684
rect 241514 176672 241520 176684
rect 241572 176672 241578 176724
rect 403618 176672 403624 176724
rect 403676 176712 403682 176724
rect 404814 176712 404820 176724
rect 403676 176684 404820 176712
rect 403676 176672 403682 176684
rect 404814 176672 404820 176684
rect 404872 176672 404878 176724
rect 135714 176604 135720 176656
rect 135772 176644 135778 176656
rect 213914 176644 213920 176656
rect 135772 176616 213920 176644
rect 135772 176604 135778 176616
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 228358 176604 228364 176656
rect 228416 176644 228422 176656
rect 229462 176644 229468 176656
rect 228416 176616 229468 176644
rect 228416 176604 228422 176616
rect 229462 176604 229468 176616
rect 229520 176604 229526 176656
rect 260190 176604 260196 176656
rect 260248 176644 260254 176656
rect 279510 176644 279516 176656
rect 260248 176616 279516 176644
rect 260248 176604 260254 176616
rect 279510 176604 279516 176616
rect 279568 176604 279574 176656
rect 158898 176196 158904 176248
rect 158956 176236 158962 176248
rect 167638 176236 167644 176248
rect 158956 176208 167644 176236
rect 158956 176196 158962 176208
rect 167638 176196 167644 176208
rect 167696 176196 167702 176248
rect 123110 176128 123116 176180
rect 123168 176168 123174 176180
rect 166258 176168 166264 176180
rect 123168 176140 166264 176168
rect 123168 176128 123174 176140
rect 166258 176128 166264 176140
rect 166316 176128 166322 176180
rect 274082 176128 274088 176180
rect 274140 176168 274146 176180
rect 281534 176168 281540 176180
rect 274140 176140 281540 176168
rect 274140 176128 274146 176140
rect 281534 176128 281540 176140
rect 281592 176128 281598 176180
rect 128170 176060 128176 176112
rect 128228 176100 128234 176112
rect 214098 176100 214104 176112
rect 128228 176072 214104 176100
rect 128228 176060 128234 176072
rect 214098 176060 214104 176072
rect 214156 176060 214162 176112
rect 225690 176060 225696 176112
rect 225748 176100 225754 176112
rect 232038 176100 232044 176112
rect 225748 176072 232044 176100
rect 225748 176060 225754 176072
rect 232038 176060 232044 176072
rect 232096 176060 232102 176112
rect 278222 176060 278228 176112
rect 278280 176100 278286 176112
rect 287054 176100 287060 176112
rect 278280 176072 287060 176100
rect 278280 176060 278286 176072
rect 287054 176060 287060 176072
rect 287112 176060 287118 176112
rect 421558 176060 421564 176112
rect 421616 176100 421622 176112
rect 430666 176100 430672 176112
rect 421616 176072 430672 176100
rect 421616 176060 421622 176072
rect 430666 176060 430672 176072
rect 430724 176060 430730 176112
rect 25498 175992 25504 176044
rect 25556 176032 25562 176044
rect 109678 176032 109684 176044
rect 25556 176004 109684 176032
rect 25556 175992 25562 176004
rect 109678 175992 109684 176004
rect 109736 175992 109742 176044
rect 113174 175992 113180 176044
rect 113232 176032 113238 176044
rect 209222 176032 209228 176044
rect 113232 176004 209228 176032
rect 113232 175992 113238 176004
rect 209222 175992 209228 176004
rect 209280 175992 209286 176044
rect 221458 175992 221464 176044
rect 221516 176032 221522 176044
rect 229370 176032 229376 176044
rect 221516 176004 229376 176032
rect 221516 175992 221522 176004
rect 229370 175992 229376 176004
rect 229428 175992 229434 176044
rect 279602 175992 279608 176044
rect 279660 176032 279666 176044
rect 289814 176032 289820 176044
rect 279660 176004 289820 176032
rect 279660 175992 279666 176004
rect 289814 175992 289820 176004
rect 289872 175992 289878 176044
rect 371878 175992 371884 176044
rect 371936 176032 371942 176044
rect 440326 176032 440332 176044
rect 371936 176004 440332 176032
rect 371936 175992 371942 176004
rect 440326 175992 440332 176004
rect 440384 175992 440390 176044
rect 98362 175924 98368 175976
rect 98420 175964 98426 175976
rect 206370 175964 206376 175976
rect 98420 175936 206376 175964
rect 98420 175924 98426 175936
rect 206370 175924 206376 175936
rect 206428 175924 206434 175976
rect 224218 175924 224224 175976
rect 224276 175964 224282 175976
rect 240410 175964 240416 175976
rect 224276 175936 240416 175964
rect 224276 175924 224282 175936
rect 240410 175924 240416 175936
rect 240468 175924 240474 175976
rect 276842 175924 276848 175976
rect 276900 175964 276906 175976
rect 291378 175964 291384 175976
rect 276900 175936 291384 175964
rect 276900 175924 276906 175936
rect 291378 175924 291384 175936
rect 291436 175924 291442 175976
rect 353938 175924 353944 175976
rect 353996 175964 354002 175976
rect 436278 175964 436284 175976
rect 353996 175936 436284 175964
rect 353996 175924 354002 175936
rect 436278 175924 436284 175936
rect 436336 175924 436342 175976
rect 425790 175856 425796 175908
rect 425848 175896 425854 175908
rect 429286 175896 429292 175908
rect 425848 175868 429292 175896
rect 425848 175856 425854 175868
rect 429286 175856 429292 175868
rect 429344 175856 429350 175908
rect 224954 175788 224960 175840
rect 225012 175828 225018 175840
rect 227714 175828 227720 175840
rect 225012 175800 227720 175828
rect 225012 175788 225018 175800
rect 227714 175788 227720 175800
rect 227772 175788 227778 175840
rect 333238 175244 333244 175296
rect 333296 175284 333302 175296
rect 333296 175256 425100 175284
rect 333296 175244 333302 175256
rect 165246 175176 165252 175228
rect 165304 175216 165310 175228
rect 213914 175216 213920 175228
rect 165304 175188 213920 175216
rect 165304 175176 165310 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 425072 175216 425100 175256
rect 427814 175216 427820 175228
rect 425072 175188 427820 175216
rect 427814 175176 427820 175188
rect 427872 175176 427878 175228
rect 164418 175108 164424 175160
rect 164476 175148 164482 175160
rect 214006 175148 214012 175160
rect 164476 175120 214012 175148
rect 164476 175108 164482 175120
rect 214006 175108 214012 175120
rect 214064 175108 214070 175160
rect 256050 174020 256056 174072
rect 256108 174060 256114 174072
rect 265342 174060 265348 174072
rect 256108 174032 265348 174060
rect 256108 174020 256114 174032
rect 265342 174020 265348 174032
rect 265400 174020 265406 174072
rect 250438 173952 250444 174004
rect 250496 173992 250502 174004
rect 265894 173992 265900 174004
rect 250496 173964 265900 173992
rect 250496 173952 250502 173964
rect 265894 173952 265900 173964
rect 265952 173952 265958 174004
rect 244918 173884 244924 173936
rect 244976 173924 244982 173936
rect 265802 173924 265808 173936
rect 244976 173896 265808 173924
rect 244976 173884 244982 173896
rect 265802 173884 265808 173896
rect 265860 173884 265866 173936
rect 322290 173884 322296 173936
rect 322348 173924 322354 173936
rect 347498 173924 347504 173936
rect 322348 173896 347504 173924
rect 322348 173884 322354 173896
rect 347498 173884 347504 173896
rect 347556 173884 347562 173936
rect 164878 173816 164884 173868
rect 164936 173856 164942 173868
rect 213914 173856 213920 173868
rect 164936 173828 213920 173856
rect 164936 173816 164942 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 231394 173816 231400 173868
rect 231452 173856 231458 173868
rect 238754 173856 238760 173868
rect 231452 173828 238760 173856
rect 231452 173816 231458 173828
rect 238754 173816 238760 173828
rect 238812 173816 238818 173868
rect 209130 173748 209136 173800
rect 209188 173788 209194 173800
rect 214006 173788 214012 173800
rect 209188 173760 214012 173788
rect 209188 173748 209194 173760
rect 214006 173748 214012 173760
rect 214064 173748 214070 173800
rect 260098 172660 260104 172712
rect 260156 172700 260162 172712
rect 265342 172700 265348 172712
rect 260156 172672 265348 172700
rect 260156 172660 260162 172672
rect 265342 172660 265348 172672
rect 265400 172660 265406 172712
rect 243814 172592 243820 172644
rect 243872 172632 243878 172644
rect 265802 172632 265808 172644
rect 243872 172604 265808 172632
rect 243872 172592 243878 172604
rect 265802 172592 265808 172604
rect 265860 172592 265866 172644
rect 239398 172524 239404 172576
rect 239456 172564 239462 172576
rect 265250 172564 265256 172576
rect 239456 172536 265256 172564
rect 239456 172524 239462 172536
rect 265250 172524 265256 172536
rect 265308 172524 265314 172576
rect 320910 172524 320916 172576
rect 320968 172564 320974 172576
rect 347498 172564 347504 172576
rect 320968 172536 347504 172564
rect 320968 172524 320974 172536
rect 347498 172524 347504 172536
rect 347556 172524 347562 172576
rect 430574 172524 430580 172576
rect 430632 172564 430638 172576
rect 433610 172564 433616 172576
rect 430632 172536 433616 172564
rect 430632 172524 430638 172536
rect 433610 172524 433616 172536
rect 433668 172524 433674 172576
rect 209314 172456 209320 172508
rect 209372 172496 209378 172508
rect 213914 172496 213920 172508
rect 209372 172468 213920 172496
rect 209372 172456 209378 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 240134 172456 240140 172508
rect 240192 172496 240198 172508
rect 241514 172496 241520 172508
rect 240192 172468 241520 172496
rect 240192 172456 240198 172468
rect 241514 172456 241520 172468
rect 241572 172456 241578 172508
rect 231670 172388 231676 172440
rect 231728 172428 231734 172440
rect 240042 172428 240048 172440
rect 231728 172400 240048 172428
rect 231728 172388 231734 172400
rect 240042 172388 240048 172400
rect 240100 172388 240106 172440
rect 231762 172320 231768 172372
rect 231820 172360 231826 172372
rect 240318 172360 240324 172372
rect 231820 172332 240324 172360
rect 231820 172320 231826 172332
rect 240318 172320 240324 172332
rect 240376 172320 240382 172372
rect 246390 171776 246396 171828
rect 246448 171816 246454 171828
rect 265986 171816 265992 171828
rect 246448 171788 265992 171816
rect 246448 171776 246454 171788
rect 265986 171776 265992 171788
rect 266044 171776 266050 171828
rect 167086 171300 167092 171352
rect 167144 171340 167150 171352
rect 169294 171340 169300 171352
rect 167144 171312 169300 171340
rect 167144 171300 167150 171312
rect 169294 171300 169300 171312
rect 169352 171300 169358 171352
rect 258718 171300 258724 171352
rect 258776 171340 258782 171352
rect 265158 171340 265164 171352
rect 258776 171312 265164 171340
rect 258776 171300 258782 171312
rect 265158 171300 265164 171312
rect 265216 171300 265222 171352
rect 242250 171096 242256 171148
rect 242308 171136 242314 171148
rect 265066 171136 265072 171148
rect 242308 171108 265072 171136
rect 242308 171096 242314 171108
rect 265066 171096 265072 171108
rect 265124 171096 265130 171148
rect 325050 171096 325056 171148
rect 325108 171136 325114 171148
rect 347498 171136 347504 171148
rect 325108 171108 347504 171136
rect 325108 171096 325114 171108
rect 347498 171096 347504 171108
rect 347556 171096 347562 171148
rect 166626 171028 166632 171080
rect 166684 171068 166690 171080
rect 213914 171068 213920 171080
rect 166684 171040 213920 171068
rect 166684 171028 166690 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 231762 171028 231768 171080
rect 231820 171068 231826 171080
rect 245654 171068 245660 171080
rect 231820 171040 245660 171068
rect 231820 171028 231826 171040
rect 245654 171028 245660 171040
rect 245712 171028 245718 171080
rect 282730 171028 282736 171080
rect 282788 171068 282794 171080
rect 291286 171068 291292 171080
rect 282788 171040 291292 171068
rect 282788 171028 282794 171040
rect 291286 171028 291292 171040
rect 291344 171028 291350 171080
rect 211982 170960 211988 171012
rect 212040 171000 212046 171012
rect 214006 171000 214012 171012
rect 212040 170972 214012 171000
rect 212040 170960 212046 170972
rect 214006 170960 214012 170972
rect 214064 170960 214070 171012
rect 282822 170960 282828 171012
rect 282880 171000 282886 171012
rect 289814 171000 289820 171012
rect 282880 170972 289820 171000
rect 282880 170960 282886 170972
rect 289814 170960 289820 170972
rect 289872 170960 289878 171012
rect 231670 170892 231676 170944
rect 231728 170932 231734 170944
rect 237558 170932 237564 170944
rect 231728 170904 237564 170932
rect 231728 170892 231734 170904
rect 237558 170892 237564 170904
rect 237616 170892 237622 170944
rect 231762 170144 231768 170196
rect 231820 170184 231826 170196
rect 237374 170184 237380 170196
rect 231820 170156 237380 170184
rect 231820 170144 231826 170156
rect 237374 170144 237380 170156
rect 237432 170144 237438 170196
rect 251910 169872 251916 169924
rect 251968 169912 251974 169924
rect 265250 169912 265256 169924
rect 251968 169884 265256 169912
rect 251968 169872 251974 169884
rect 265250 169872 265256 169884
rect 265308 169872 265314 169924
rect 250530 169804 250536 169856
rect 250588 169844 250594 169856
rect 265434 169844 265440 169856
rect 250588 169816 265440 169844
rect 250588 169804 250594 169816
rect 265434 169804 265440 169816
rect 265492 169804 265498 169856
rect 249702 169736 249708 169788
rect 249760 169776 249766 169788
rect 265618 169776 265624 169788
rect 249760 169748 265624 169776
rect 249760 169736 249766 169748
rect 265618 169736 265624 169748
rect 265676 169736 265682 169788
rect 166258 169668 166264 169720
rect 166316 169708 166322 169720
rect 214006 169708 214012 169720
rect 166316 169680 214012 169708
rect 166316 169668 166322 169680
rect 214006 169668 214012 169680
rect 214064 169668 214070 169720
rect 231670 169668 231676 169720
rect 231728 169708 231734 169720
rect 241606 169708 241612 169720
rect 231728 169680 241612 169708
rect 231728 169668 231734 169680
rect 241606 169668 241612 169680
rect 241664 169668 241670 169720
rect 170582 169600 170588 169652
rect 170640 169640 170646 169652
rect 213914 169640 213920 169652
rect 170640 169612 213920 169640
rect 170640 169600 170646 169612
rect 213914 169600 213920 169612
rect 213972 169600 213978 169652
rect 231394 169600 231400 169652
rect 231452 169640 231458 169652
rect 240134 169640 240140 169652
rect 231452 169612 240140 169640
rect 231452 169600 231458 169612
rect 240134 169600 240140 169612
rect 240192 169600 240198 169652
rect 231762 169532 231768 169584
rect 231820 169572 231826 169584
rect 240226 169572 240232 169584
rect 231820 169544 240232 169572
rect 231820 169532 231826 169544
rect 240226 169532 240232 169544
rect 240284 169532 240290 169584
rect 258994 169464 259000 169516
rect 259052 169504 259058 169516
rect 265342 169504 265348 169516
rect 259052 169476 265348 169504
rect 259052 169464 259058 169476
rect 265342 169464 265348 169476
rect 265400 169464 265406 169516
rect 281902 168852 281908 168904
rect 281960 168892 281966 168904
rect 287054 168892 287060 168904
rect 281960 168864 287060 168892
rect 281960 168852 281966 168864
rect 287054 168852 287060 168864
rect 287112 168852 287118 168904
rect 240962 168444 240968 168496
rect 241020 168484 241026 168496
rect 241020 168456 243216 168484
rect 241020 168444 241026 168456
rect 240870 168376 240876 168428
rect 240928 168416 240934 168428
rect 243078 168416 243084 168428
rect 240928 168388 243084 168416
rect 240928 168376 240934 168388
rect 243078 168376 243084 168388
rect 243136 168376 243142 168428
rect 243188 168416 243216 168456
rect 246666 168444 246672 168496
rect 246724 168484 246730 168496
rect 265342 168484 265348 168496
rect 246724 168456 265348 168484
rect 246724 168444 246730 168456
rect 265342 168444 265348 168456
rect 265400 168444 265406 168496
rect 265894 168416 265900 168428
rect 243188 168388 265900 168416
rect 265894 168376 265900 168388
rect 265952 168376 265958 168428
rect 307018 168376 307024 168428
rect 307076 168416 307082 168428
rect 347038 168416 347044 168428
rect 307076 168388 347044 168416
rect 307076 168376 307082 168388
rect 347038 168376 347044 168388
rect 347096 168376 347102 168428
rect 166534 168308 166540 168360
rect 166592 168348 166598 168360
rect 214006 168348 214012 168360
rect 166592 168320 214012 168348
rect 166592 168308 166598 168320
rect 214006 168308 214012 168320
rect 214064 168308 214070 168360
rect 231762 168308 231768 168360
rect 231820 168348 231826 168360
rect 238846 168348 238852 168360
rect 231820 168320 238852 168348
rect 231820 168308 231826 168320
rect 238846 168308 238852 168320
rect 238904 168308 238910 168360
rect 281902 168308 281908 168360
rect 281960 168348 281966 168360
rect 295426 168348 295432 168360
rect 281960 168320 295432 168348
rect 281960 168308 281966 168320
rect 295426 168308 295432 168320
rect 295484 168308 295490 168360
rect 167822 168240 167828 168292
rect 167880 168280 167886 168292
rect 213914 168280 213920 168292
rect 167880 168252 213920 168280
rect 167880 168240 167886 168252
rect 213914 168240 213920 168252
rect 213972 168240 213978 168292
rect 282362 168240 282368 168292
rect 282420 168280 282426 168292
rect 289998 168280 290004 168292
rect 282420 168252 290004 168280
rect 282420 168240 282426 168252
rect 289998 168240 290004 168252
rect 290056 168240 290062 168292
rect 231210 167968 231216 168020
rect 231268 168008 231274 168020
rect 237466 168008 237472 168020
rect 231268 167980 237472 168008
rect 231268 167968 231274 167980
rect 237466 167968 237472 167980
rect 237524 167968 237530 168020
rect 243722 167628 243728 167680
rect 243780 167668 243786 167680
rect 265802 167668 265808 167680
rect 243780 167640 265808 167668
rect 243780 167628 243786 167640
rect 265802 167628 265808 167640
rect 265860 167628 265866 167680
rect 249058 167152 249064 167204
rect 249116 167192 249122 167204
rect 265250 167192 265256 167204
rect 249116 167164 265256 167192
rect 249116 167152 249122 167164
rect 265250 167152 265256 167164
rect 265308 167152 265314 167204
rect 242158 167084 242164 167136
rect 242216 167124 242222 167136
rect 249702 167124 249708 167136
rect 242216 167096 249708 167124
rect 242216 167084 242222 167096
rect 249702 167084 249708 167096
rect 249760 167084 249766 167136
rect 238018 167016 238024 167068
rect 238076 167056 238082 167068
rect 265526 167056 265532 167068
rect 238076 167028 265532 167056
rect 238076 167016 238082 167028
rect 265526 167016 265532 167028
rect 265584 167016 265590 167068
rect 327810 167016 327816 167068
rect 327868 167056 327874 167068
rect 347498 167056 347504 167068
rect 327868 167028 347504 167056
rect 327868 167016 327874 167028
rect 347498 167016 347504 167028
rect 347556 167016 347562 167068
rect 167730 166948 167736 167000
rect 167788 166988 167794 167000
rect 213914 166988 213920 167000
rect 167788 166960 213920 166988
rect 167788 166948 167794 166960
rect 213914 166948 213920 166960
rect 213972 166948 213978 167000
rect 231762 166948 231768 167000
rect 231820 166988 231826 167000
rect 241790 166988 241796 167000
rect 231820 166960 241796 166988
rect 231820 166948 231826 166960
rect 241790 166948 241796 166960
rect 241848 166948 241854 167000
rect 282086 166948 282092 167000
rect 282144 166988 282150 167000
rect 295518 166988 295524 167000
rect 282144 166960 295524 166988
rect 282144 166948 282150 166960
rect 295518 166948 295524 166960
rect 295576 166948 295582 167000
rect 211798 166880 211804 166932
rect 211856 166920 211862 166932
rect 214098 166920 214104 166932
rect 211856 166892 214104 166920
rect 211856 166880 211862 166892
rect 214098 166880 214104 166892
rect 214156 166880 214162 166932
rect 231486 166880 231492 166932
rect 231544 166920 231550 166932
rect 238938 166920 238944 166932
rect 231544 166892 238944 166920
rect 231544 166880 231550 166892
rect 238938 166880 238944 166892
rect 238996 166880 239002 166932
rect 429102 166812 429108 166864
rect 429160 166852 429166 166864
rect 433426 166852 433432 166864
rect 429160 166824 433432 166852
rect 429160 166812 429166 166824
rect 433426 166812 433432 166824
rect 433484 166812 433490 166864
rect 230566 166268 230572 166320
rect 230624 166308 230630 166320
rect 230934 166308 230940 166320
rect 230624 166280 230940 166308
rect 230624 166268 230630 166280
rect 230934 166268 230940 166280
rect 230992 166268 230998 166320
rect 231578 166268 231584 166320
rect 231636 166308 231642 166320
rect 237650 166308 237656 166320
rect 231636 166280 237656 166308
rect 231636 166268 231642 166280
rect 237650 166268 237656 166280
rect 237708 166268 237714 166320
rect 280798 166268 280804 166320
rect 280856 166308 280862 166320
rect 281626 166308 281632 166320
rect 280856 166280 281632 166308
rect 280856 166268 280862 166280
rect 281626 166268 281632 166280
rect 281684 166268 281690 166320
rect 314010 166268 314016 166320
rect 314068 166308 314074 166320
rect 346670 166308 346676 166320
rect 314068 166280 346676 166308
rect 314068 166268 314074 166280
rect 346670 166268 346676 166280
rect 346728 166308 346734 166320
rect 346854 166308 346860 166320
rect 346728 166280 346860 166308
rect 346728 166268 346734 166280
rect 346854 166268 346860 166280
rect 346912 166268 346918 166320
rect 263134 165724 263140 165776
rect 263192 165764 263198 165776
rect 265802 165764 265808 165776
rect 263192 165736 265808 165764
rect 263192 165724 263198 165736
rect 265802 165724 265808 165736
rect 265860 165724 265866 165776
rect 253198 165656 253204 165708
rect 253256 165696 253262 165708
rect 265618 165696 265624 165708
rect 253256 165668 265624 165696
rect 253256 165656 253262 165668
rect 265618 165656 265624 165668
rect 265676 165656 265682 165708
rect 238386 165588 238392 165640
rect 238444 165628 238450 165640
rect 265894 165628 265900 165640
rect 238444 165600 265900 165628
rect 238444 165588 238450 165600
rect 265894 165588 265900 165600
rect 265952 165588 265958 165640
rect 166442 165520 166448 165572
rect 166500 165560 166506 165572
rect 213914 165560 213920 165572
rect 166500 165532 213920 165560
rect 166500 165520 166506 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 231026 165520 231032 165572
rect 231084 165560 231090 165572
rect 249794 165560 249800 165572
rect 231084 165532 249800 165560
rect 231084 165520 231090 165532
rect 249794 165520 249800 165532
rect 249852 165520 249858 165572
rect 282086 165520 282092 165572
rect 282144 165560 282150 165572
rect 292666 165560 292672 165572
rect 282144 165532 292672 165560
rect 282144 165520 282150 165532
rect 292666 165520 292672 165532
rect 292724 165520 292730 165572
rect 167914 165452 167920 165504
rect 167972 165492 167978 165504
rect 214006 165492 214012 165504
rect 167972 165464 214012 165492
rect 167972 165452 167978 165464
rect 214006 165452 214012 165464
rect 214064 165452 214070 165504
rect 231118 165452 231124 165504
rect 231176 165492 231182 165504
rect 233418 165492 233424 165504
rect 231176 165464 233424 165492
rect 231176 165452 231182 165464
rect 233418 165452 233424 165464
rect 233476 165452 233482 165504
rect 247862 164840 247868 164892
rect 247920 164880 247926 164892
rect 265434 164880 265440 164892
rect 247920 164852 265440 164880
rect 247920 164840 247926 164852
rect 265434 164840 265440 164852
rect 265492 164840 265498 164892
rect 327718 164840 327724 164892
rect 327776 164880 327782 164892
rect 339494 164880 339500 164892
rect 327776 164852 339500 164880
rect 327776 164840 327782 164852
rect 339494 164840 339500 164852
rect 339552 164840 339558 164892
rect 467098 164840 467104 164892
rect 467156 164880 467162 164892
rect 580166 164880 580172 164892
rect 467156 164852 580172 164880
rect 467156 164840 467162 164852
rect 580166 164840 580172 164852
rect 580224 164840 580230 164892
rect 282362 164228 282368 164280
rect 282420 164268 282426 164280
rect 288526 164268 288532 164280
rect 282420 164240 288532 164268
rect 282420 164228 282426 164240
rect 288526 164228 288532 164240
rect 288584 164228 288590 164280
rect 339494 164228 339500 164280
rect 339552 164268 339558 164280
rect 347498 164268 347504 164280
rect 339552 164240 347504 164268
rect 339552 164228 339558 164240
rect 347498 164228 347504 164240
rect 347556 164228 347562 164280
rect 198182 164160 198188 164212
rect 198240 164200 198246 164212
rect 214006 164200 214012 164212
rect 198240 164172 214012 164200
rect 198240 164160 198246 164172
rect 214006 164160 214012 164172
rect 214064 164160 214070 164212
rect 231762 164160 231768 164212
rect 231820 164200 231826 164212
rect 244458 164200 244464 164212
rect 231820 164172 244464 164200
rect 231820 164160 231826 164172
rect 244458 164160 244464 164172
rect 244516 164160 244522 164212
rect 282178 164160 282184 164212
rect 282236 164200 282242 164212
rect 299566 164200 299572 164212
rect 282236 164172 299572 164200
rect 282236 164160 282242 164172
rect 299566 164160 299572 164172
rect 299624 164160 299630 164212
rect 430574 164160 430580 164212
rect 430632 164200 430638 164212
rect 436370 164200 436376 164212
rect 430632 164172 436376 164200
rect 430632 164160 430638 164172
rect 436370 164160 436376 164172
rect 436428 164200 436434 164212
rect 436646 164200 436652 164212
rect 436428 164172 436652 164200
rect 436428 164160 436434 164172
rect 436646 164160 436652 164172
rect 436704 164160 436710 164212
rect 209222 164092 209228 164144
rect 209280 164132 209286 164144
rect 213914 164132 213920 164144
rect 209280 164104 213920 164132
rect 209280 164092 209286 164104
rect 213914 164092 213920 164104
rect 213972 164092 213978 164144
rect 231670 164092 231676 164144
rect 231728 164132 231734 164144
rect 244274 164132 244280 164144
rect 231728 164104 244280 164132
rect 231728 164092 231734 164104
rect 244274 164092 244280 164104
rect 244332 164092 244338 164144
rect 282822 164092 282828 164144
rect 282880 164132 282886 164144
rect 291378 164132 291384 164144
rect 282880 164104 291384 164132
rect 282880 164092 282886 164104
rect 291378 164092 291384 164104
rect 291436 164092 291442 164144
rect 231486 164024 231492 164076
rect 231544 164064 231550 164076
rect 239030 164064 239036 164076
rect 231544 164036 239036 164064
rect 231544 164024 231550 164036
rect 239030 164024 239036 164036
rect 239088 164024 239094 164076
rect 229922 163684 229928 163736
rect 229980 163724 229986 163736
rect 234890 163724 234896 163736
rect 229980 163696 234896 163724
rect 229980 163684 229986 163696
rect 234890 163684 234896 163696
rect 234948 163684 234954 163736
rect 229738 163480 229744 163532
rect 229796 163520 229802 163532
rect 242894 163520 242900 163532
rect 229796 163492 242900 163520
rect 229796 163480 229802 163492
rect 242894 163480 242900 163492
rect 242952 163480 242958 163532
rect 245010 163480 245016 163532
rect 245068 163520 245074 163532
rect 265158 163520 265164 163532
rect 245068 163492 265164 163520
rect 245068 163480 245074 163492
rect 265158 163480 265164 163492
rect 265216 163480 265222 163532
rect 336182 163480 336188 163532
rect 336240 163520 336246 163532
rect 345014 163520 345020 163532
rect 336240 163492 345020 163520
rect 336240 163480 336246 163492
rect 345014 163480 345020 163492
rect 345072 163520 345078 163532
rect 346670 163520 346676 163532
rect 345072 163492 346676 163520
rect 345072 163480 345078 163492
rect 346670 163480 346676 163492
rect 346728 163480 346734 163532
rect 436646 163480 436652 163532
rect 436704 163520 436710 163532
rect 471238 163520 471244 163532
rect 436704 163492 471244 163520
rect 436704 163480 436710 163492
rect 471238 163480 471244 163492
rect 471296 163480 471302 163532
rect 240134 163140 240140 163192
rect 240192 163180 240198 163192
rect 245746 163180 245752 163192
rect 240192 163152 245752 163180
rect 240192 163140 240198 163152
rect 245746 163140 245752 163152
rect 245804 163140 245810 163192
rect 260190 162936 260196 162988
rect 260248 162976 260254 162988
rect 265618 162976 265624 162988
rect 260248 162948 265624 162976
rect 260248 162936 260254 162948
rect 265618 162936 265624 162948
rect 265676 162936 265682 162988
rect 234154 162868 234160 162920
rect 234212 162908 234218 162920
rect 265526 162908 265532 162920
rect 234212 162880 265532 162908
rect 234212 162868 234218 162880
rect 265526 162868 265532 162880
rect 265584 162868 265590 162920
rect 170490 162800 170496 162852
rect 170548 162840 170554 162852
rect 213914 162840 213920 162852
rect 170548 162812 213920 162840
rect 170548 162800 170554 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 282086 162800 282092 162852
rect 282144 162840 282150 162852
rect 298094 162840 298100 162852
rect 282144 162812 298100 162840
rect 282144 162800 282150 162812
rect 298094 162800 298100 162812
rect 298152 162800 298158 162852
rect 430574 162800 430580 162852
rect 430632 162840 430638 162852
rect 434990 162840 434996 162852
rect 430632 162812 434996 162840
rect 430632 162800 430638 162812
rect 434990 162800 434996 162812
rect 435048 162840 435054 162852
rect 436002 162840 436008 162852
rect 435048 162812 436008 162840
rect 435048 162800 435054 162812
rect 436002 162800 436008 162812
rect 436060 162800 436066 162852
rect 231762 162732 231768 162784
rect 231820 162772 231826 162784
rect 244366 162772 244372 162784
rect 231820 162744 244372 162772
rect 231820 162732 231826 162744
rect 244366 162732 244372 162744
rect 244424 162732 244430 162784
rect 282822 162732 282828 162784
rect 282880 162772 282886 162784
rect 292758 162772 292764 162784
rect 282880 162744 292764 162772
rect 282880 162732 282886 162744
rect 292758 162732 292764 162744
rect 292816 162732 292822 162784
rect 430574 162188 430580 162240
rect 430632 162228 430638 162240
rect 439130 162228 439136 162240
rect 430632 162200 439136 162228
rect 430632 162188 430638 162200
rect 439130 162188 439136 162200
rect 439188 162188 439194 162240
rect 436002 162120 436008 162172
rect 436060 162160 436066 162172
rect 464338 162160 464344 162172
rect 436060 162132 464344 162160
rect 436060 162120 436066 162132
rect 464338 162120 464344 162132
rect 464396 162120 464402 162172
rect 234062 161780 234068 161832
rect 234120 161820 234126 161832
rect 240410 161820 240416 161832
rect 234120 161792 240416 161820
rect 234120 161780 234126 161792
rect 240410 161780 240416 161792
rect 240468 161780 240474 161832
rect 253290 161576 253296 161628
rect 253348 161616 253354 161628
rect 264514 161616 264520 161628
rect 253348 161588 264520 161616
rect 253348 161576 253354 161588
rect 264514 161576 264520 161588
rect 264572 161576 264578 161628
rect 246298 161508 246304 161560
rect 246356 161548 246362 161560
rect 265710 161548 265716 161560
rect 246356 161520 265716 161548
rect 246356 161508 246362 161520
rect 265710 161508 265716 161520
rect 265768 161508 265774 161560
rect 238110 161440 238116 161492
rect 238168 161480 238174 161492
rect 265802 161480 265808 161492
rect 238168 161452 265808 161480
rect 238168 161440 238174 161452
rect 265802 161440 265808 161452
rect 265860 161440 265866 161492
rect 231762 161372 231768 161424
rect 231820 161412 231826 161424
rect 241698 161412 241704 161424
rect 231820 161384 241704 161412
rect 231820 161372 231826 161384
rect 241698 161372 241704 161384
rect 241756 161372 241762 161424
rect 282730 161372 282736 161424
rect 282788 161412 282794 161424
rect 293954 161412 293960 161424
rect 282788 161384 293960 161412
rect 282788 161372 282794 161384
rect 293954 161372 293960 161384
rect 294012 161372 294018 161424
rect 343634 161372 343640 161424
rect 343692 161412 343698 161424
rect 347498 161412 347504 161424
rect 343692 161384 347504 161412
rect 343692 161372 343698 161384
rect 347498 161372 347504 161384
rect 347556 161372 347562 161424
rect 430574 161372 430580 161424
rect 430632 161412 430638 161424
rect 444466 161412 444472 161424
rect 430632 161384 444472 161412
rect 430632 161372 430638 161384
rect 444466 161372 444472 161384
rect 444524 161372 444530 161424
rect 231302 161304 231308 161356
rect 231360 161344 231366 161356
rect 238846 161344 238852 161356
rect 231360 161316 238852 161344
rect 231360 161304 231366 161316
rect 238846 161304 238852 161316
rect 238904 161304 238910 161356
rect 169294 160692 169300 160744
rect 169352 160732 169358 160744
rect 214558 160732 214564 160744
rect 169352 160704 214564 160732
rect 169352 160692 169358 160704
rect 214558 160692 214564 160704
rect 214616 160692 214622 160744
rect 318150 160692 318156 160744
rect 318208 160732 318214 160744
rect 343634 160732 343640 160744
rect 318208 160704 343640 160732
rect 318208 160692 318214 160704
rect 343634 160692 343640 160704
rect 343692 160692 343698 160744
rect 282822 160420 282828 160472
rect 282880 160460 282886 160472
rect 288710 160460 288716 160472
rect 282880 160432 288716 160460
rect 282880 160420 282886 160432
rect 288710 160420 288716 160432
rect 288768 160420 288774 160472
rect 257338 160216 257344 160268
rect 257396 160256 257402 160268
rect 265618 160256 265624 160268
rect 257396 160228 265624 160256
rect 257396 160216 257402 160228
rect 265618 160216 265624 160228
rect 265676 160216 265682 160268
rect 240778 160148 240784 160200
rect 240836 160188 240842 160200
rect 265342 160188 265348 160200
rect 240836 160160 265348 160188
rect 240836 160148 240842 160160
rect 265342 160148 265348 160160
rect 265400 160148 265406 160200
rect 239490 160080 239496 160132
rect 239548 160120 239554 160132
rect 265802 160120 265808 160132
rect 239548 160092 265808 160120
rect 239548 160080 239554 160092
rect 265802 160080 265808 160092
rect 265860 160080 265866 160132
rect 444466 160080 444472 160132
rect 444524 160120 444530 160132
rect 447778 160120 447784 160132
rect 444524 160092 447784 160120
rect 444524 160080 444530 160092
rect 447778 160080 447784 160092
rect 447836 160080 447842 160132
rect 169110 160012 169116 160064
rect 169168 160052 169174 160064
rect 213914 160052 213920 160064
rect 169168 160024 213920 160052
rect 169168 160012 169174 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 231762 160012 231768 160064
rect 231820 160052 231826 160064
rect 245838 160052 245844 160064
rect 231820 160024 245844 160052
rect 231820 160012 231826 160024
rect 245838 160012 245844 160024
rect 245896 160012 245902 160064
rect 282086 160012 282092 160064
rect 282144 160052 282150 160064
rect 313274 160052 313280 160064
rect 282144 160024 313280 160052
rect 282144 160012 282150 160024
rect 313274 160012 313280 160024
rect 313332 160012 313338 160064
rect 430574 160012 430580 160064
rect 430632 160052 430638 160064
rect 454034 160052 454040 160064
rect 430632 160024 454040 160052
rect 430632 160012 430638 160024
rect 454034 160012 454040 160024
rect 454092 160052 454098 160064
rect 467098 160052 467104 160064
rect 454092 160024 467104 160052
rect 454092 160012 454098 160024
rect 467098 160012 467104 160024
rect 467156 160012 467162 160064
rect 173250 159944 173256 159996
rect 173308 159984 173314 159996
rect 214006 159984 214012 159996
rect 173308 159956 214012 159984
rect 173308 159944 173314 159956
rect 214006 159944 214012 159956
rect 214064 159944 214070 159996
rect 231026 159944 231032 159996
rect 231084 159984 231090 159996
rect 240134 159984 240140 159996
rect 231084 159956 240140 159984
rect 231084 159944 231090 159956
rect 240134 159944 240140 159956
rect 240192 159944 240198 159996
rect 231578 159876 231584 159928
rect 231636 159916 231642 159928
rect 234062 159916 234068 159928
rect 231636 159888 234068 159916
rect 231636 159876 231642 159888
rect 234062 159876 234068 159888
rect 234120 159876 234126 159928
rect 250622 159332 250628 159384
rect 250680 159372 250686 159384
rect 265986 159372 265992 159384
rect 250680 159344 265992 159372
rect 250680 159332 250686 159344
rect 265986 159332 265992 159344
rect 266044 159332 266050 159384
rect 316770 159332 316776 159384
rect 316828 159372 316834 159384
rect 340874 159372 340880 159384
rect 316828 159344 340880 159372
rect 316828 159332 316834 159344
rect 340874 159332 340880 159344
rect 340932 159372 340938 159384
rect 347498 159372 347504 159384
rect 340932 159344 347504 159372
rect 340932 159332 340938 159344
rect 347498 159332 347504 159344
rect 347556 159332 347562 159384
rect 245194 158788 245200 158840
rect 245252 158828 245258 158840
rect 265802 158828 265808 158840
rect 245252 158800 265808 158828
rect 245252 158788 245258 158800
rect 265802 158788 265808 158800
rect 265860 158788 265866 158840
rect 239674 158720 239680 158772
rect 239732 158760 239738 158772
rect 265710 158760 265716 158772
rect 239732 158732 265716 158760
rect 239732 158720 239738 158732
rect 265710 158720 265716 158732
rect 265768 158720 265774 158772
rect 171778 158652 171784 158704
rect 171836 158692 171842 158704
rect 213914 158692 213920 158704
rect 171836 158664 213920 158692
rect 171836 158652 171842 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 231762 158652 231768 158704
rect 231820 158692 231826 158704
rect 252554 158692 252560 158704
rect 231820 158664 252560 158692
rect 231820 158652 231826 158664
rect 252554 158652 252560 158664
rect 252612 158652 252618 158704
rect 282730 158652 282736 158704
rect 282788 158692 282794 158704
rect 302418 158692 302424 158704
rect 282788 158664 302424 158692
rect 282788 158652 282794 158664
rect 302418 158652 302424 158664
rect 302476 158652 302482 158704
rect 430574 158652 430580 158704
rect 430632 158692 430638 158704
rect 450538 158692 450544 158704
rect 430632 158664 450544 158692
rect 430632 158652 430638 158664
rect 450538 158652 450544 158664
rect 450596 158652 450602 158704
rect 231210 158584 231216 158636
rect 231268 158624 231274 158636
rect 240870 158624 240876 158636
rect 231268 158596 240876 158624
rect 231268 158584 231274 158596
rect 240870 158584 240876 158596
rect 240928 158584 240934 158636
rect 282822 158584 282828 158636
rect 282880 158624 282886 158636
rect 300854 158624 300860 158636
rect 282880 158596 300860 158624
rect 282880 158584 282886 158596
rect 300854 158584 300860 158596
rect 300912 158584 300918 158636
rect 324958 157972 324964 158024
rect 325016 158012 325022 158024
rect 342346 158012 342352 158024
rect 325016 157984 342352 158012
rect 325016 157972 325022 157984
rect 342346 157972 342352 157984
rect 342404 157972 342410 158024
rect 261570 157496 261576 157548
rect 261628 157536 261634 157548
rect 265894 157536 265900 157548
rect 261628 157508 265900 157536
rect 261628 157496 261634 157508
rect 265894 157496 265900 157508
rect 265952 157496 265958 157548
rect 245286 157428 245292 157480
rect 245344 157468 245350 157480
rect 265710 157468 265716 157480
rect 245344 157440 265716 157468
rect 245344 157428 245350 157440
rect 265710 157428 265716 157440
rect 265768 157428 265774 157480
rect 342346 157428 342352 157480
rect 342404 157468 342410 157480
rect 347498 157468 347504 157480
rect 342404 157440 347504 157468
rect 342404 157428 342410 157440
rect 347498 157428 347504 157440
rect 347556 157428 347562 157480
rect 237374 157360 237380 157412
rect 237432 157400 237438 157412
rect 265618 157400 265624 157412
rect 237432 157372 265624 157400
rect 237432 157360 237438 157372
rect 265618 157360 265624 157372
rect 265676 157360 265682 157412
rect 169202 157292 169208 157344
rect 169260 157332 169266 157344
rect 213914 157332 213920 157344
rect 169260 157304 213920 157332
rect 169260 157292 169266 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 231762 157292 231768 157344
rect 231820 157332 231826 157344
rect 256694 157332 256700 157344
rect 231820 157304 256700 157332
rect 231820 157292 231826 157304
rect 256694 157292 256700 157304
rect 256752 157292 256758 157344
rect 282086 157292 282092 157344
rect 282144 157332 282150 157344
rect 303798 157332 303804 157344
rect 282144 157304 303804 157332
rect 282144 157292 282150 157304
rect 303798 157292 303804 157304
rect 303856 157292 303862 157344
rect 430574 157292 430580 157344
rect 430632 157332 430638 157344
rect 475378 157332 475384 157344
rect 430632 157304 475384 157332
rect 430632 157292 430638 157304
rect 475378 157292 475384 157304
rect 475436 157292 475442 157344
rect 231118 157224 231124 157276
rect 231176 157264 231182 157276
rect 248414 157264 248420 157276
rect 231176 157236 248420 157264
rect 231176 157224 231182 157236
rect 248414 157224 248420 157236
rect 248472 157224 248478 157276
rect 231578 156748 231584 156800
rect 231636 156788 231642 156800
rect 234706 156788 234712 156800
rect 231636 156760 234712 156788
rect 231636 156748 231642 156760
rect 234706 156748 234712 156760
rect 234764 156748 234770 156800
rect 232682 156680 232688 156732
rect 232740 156720 232746 156732
rect 251358 156720 251364 156732
rect 232740 156692 251364 156720
rect 232740 156680 232746 156692
rect 251358 156680 251364 156692
rect 251416 156680 251422 156732
rect 242434 156612 242440 156664
rect 242492 156652 242498 156664
rect 265158 156652 265164 156664
rect 242492 156624 265164 156652
rect 242492 156612 242498 156624
rect 265158 156612 265164 156624
rect 265216 156612 265222 156664
rect 336090 156068 336096 156120
rect 336148 156108 336154 156120
rect 343634 156108 343640 156120
rect 336148 156080 343640 156108
rect 336148 156068 336154 156080
rect 343634 156068 343640 156080
rect 343692 156108 343698 156120
rect 347038 156108 347044 156120
rect 343692 156080 347044 156108
rect 343692 156068 343698 156080
rect 347038 156068 347044 156080
rect 347096 156068 347102 156120
rect 252094 156000 252100 156052
rect 252152 156040 252158 156052
rect 265526 156040 265532 156052
rect 252152 156012 265532 156040
rect 252152 156000 252158 156012
rect 265526 156000 265532 156012
rect 265584 156000 265590 156052
rect 240870 155932 240876 155984
rect 240928 155972 240934 155984
rect 265894 155972 265900 155984
rect 240928 155944 265900 155972
rect 240928 155932 240934 155944
rect 265894 155932 265900 155944
rect 265952 155932 265958 155984
rect 281534 155932 281540 155984
rect 281592 155972 281598 155984
rect 283098 155972 283104 155984
rect 281592 155944 283104 155972
rect 281592 155932 281598 155944
rect 283098 155932 283104 155944
rect 283156 155932 283162 155984
rect 173342 155864 173348 155916
rect 173400 155904 173406 155916
rect 214006 155904 214012 155916
rect 173400 155876 214012 155904
rect 173400 155864 173406 155876
rect 214006 155864 214012 155876
rect 214064 155864 214070 155916
rect 231486 155864 231492 155916
rect 231544 155904 231550 155916
rect 247218 155904 247224 155916
rect 231544 155876 247224 155904
rect 231544 155864 231550 155876
rect 247218 155864 247224 155876
rect 247276 155864 247282 155916
rect 282362 155864 282368 155916
rect 282420 155904 282426 155916
rect 307938 155904 307944 155916
rect 282420 155876 307944 155904
rect 282420 155864 282426 155876
rect 307938 155864 307944 155876
rect 307996 155864 308002 155916
rect 430850 155864 430856 155916
rect 430908 155904 430914 155916
rect 482278 155904 482284 155916
rect 430908 155876 482284 155904
rect 430908 155864 430914 155876
rect 482278 155864 482284 155876
rect 482336 155864 482342 155916
rect 206370 155796 206376 155848
rect 206428 155836 206434 155848
rect 213914 155836 213920 155848
rect 206428 155808 213920 155836
rect 206428 155796 206434 155808
rect 213914 155796 213920 155808
rect 213972 155796 213978 155848
rect 231762 155796 231768 155848
rect 231820 155836 231826 155848
rect 242986 155836 242992 155848
rect 231820 155808 242992 155836
rect 231820 155796 231826 155808
rect 242986 155796 242992 155808
rect 243044 155796 243050 155848
rect 282086 155796 282092 155848
rect 282144 155836 282150 155848
rect 306558 155836 306564 155848
rect 282144 155808 306564 155836
rect 282144 155796 282150 155808
rect 306558 155796 306564 155808
rect 306616 155796 306622 155848
rect 430574 155796 430580 155848
rect 430632 155836 430638 155848
rect 438946 155836 438952 155848
rect 430632 155808 438952 155836
rect 430632 155796 430638 155808
rect 438946 155796 438952 155808
rect 439004 155796 439010 155848
rect 256326 155252 256332 155304
rect 256384 155292 256390 155304
rect 265342 155292 265348 155304
rect 256384 155264 265348 155292
rect 256384 155252 256390 155264
rect 265342 155252 265348 155264
rect 265400 155252 265406 155304
rect 238202 155184 238208 155236
rect 238260 155224 238266 155236
rect 265986 155224 265992 155236
rect 238260 155196 265992 155224
rect 238260 155184 238266 155196
rect 265986 155184 265992 155196
rect 266044 155184 266050 155236
rect 241146 154572 241152 154624
rect 241204 154612 241210 154624
rect 265802 154612 265808 154624
rect 241204 154584 265808 154612
rect 241204 154572 241210 154584
rect 265802 154572 265808 154584
rect 265860 154572 265866 154624
rect 231762 154504 231768 154556
rect 231820 154544 231826 154556
rect 251266 154544 251272 154556
rect 231820 154516 251272 154544
rect 231820 154504 231826 154516
rect 251266 154504 251272 154516
rect 251324 154504 251330 154556
rect 282454 154504 282460 154556
rect 282512 154544 282518 154556
rect 310698 154544 310704 154556
rect 282512 154516 310704 154544
rect 282512 154504 282518 154516
rect 310698 154504 310704 154516
rect 310756 154504 310762 154556
rect 430574 154504 430580 154556
rect 430632 154544 430638 154556
rect 479518 154544 479524 154556
rect 430632 154516 479524 154544
rect 430632 154504 430638 154516
rect 479518 154504 479524 154516
rect 479576 154504 479582 154556
rect 231670 154436 231676 154488
rect 231728 154476 231734 154488
rect 248506 154476 248512 154488
rect 231728 154448 248512 154476
rect 231728 154436 231734 154448
rect 248506 154436 248512 154448
rect 248564 154436 248570 154488
rect 281902 154164 281908 154216
rect 281960 154204 281966 154216
rect 285950 154204 285956 154216
rect 281960 154176 285956 154204
rect 281960 154164 281966 154176
rect 285950 154164 285956 154176
rect 286008 154164 286014 154216
rect 252186 153824 252192 153876
rect 252244 153864 252250 153876
rect 265986 153864 265992 153876
rect 252244 153836 265992 153864
rect 252244 153824 252250 153836
rect 265986 153824 265992 153836
rect 266044 153824 266050 153876
rect 309778 153824 309784 153876
rect 309836 153864 309842 153876
rect 345014 153864 345020 153876
rect 309836 153836 345020 153864
rect 309836 153824 309842 153836
rect 345014 153824 345020 153836
rect 345072 153864 345078 153876
rect 346670 153864 346676 153876
rect 345072 153836 346676 153864
rect 345072 153824 345078 153836
rect 346670 153824 346676 153836
rect 346728 153824 346734 153876
rect 231118 153756 231124 153808
rect 231176 153796 231182 153808
rect 238386 153796 238392 153808
rect 231176 153768 238392 153796
rect 231176 153756 231182 153768
rect 238386 153756 238392 153768
rect 238444 153756 238450 153808
rect 198090 153280 198096 153332
rect 198148 153320 198154 153332
rect 214006 153320 214012 153332
rect 198148 153292 214012 153320
rect 198148 153280 198154 153292
rect 214006 153280 214012 153292
rect 214064 153280 214070 153332
rect 238294 153280 238300 153332
rect 238352 153320 238358 153332
rect 265802 153320 265808 153332
rect 238352 153292 265808 153320
rect 238352 153280 238358 153292
rect 265802 153280 265808 153292
rect 265860 153280 265866 153332
rect 187050 153212 187056 153264
rect 187108 153252 187114 153264
rect 213914 153252 213920 153264
rect 187108 153224 213920 153252
rect 187108 153212 187114 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 236730 153212 236736 153264
rect 236788 153252 236794 153264
rect 265894 153252 265900 153264
rect 236788 153224 265900 153252
rect 236788 153212 236794 153224
rect 265894 153212 265900 153224
rect 265952 153212 265958 153264
rect 231762 153144 231768 153196
rect 231820 153184 231826 153196
rect 260834 153184 260840 153196
rect 231820 153156 260840 153184
rect 231820 153144 231826 153156
rect 260834 153144 260840 153156
rect 260892 153144 260898 153196
rect 430574 153144 430580 153196
rect 430632 153184 430638 153196
rect 457438 153184 457444 153196
rect 430632 153156 457444 153184
rect 430632 153144 430638 153156
rect 457438 153144 457444 153156
rect 457496 153144 457502 153196
rect 230474 152532 230480 152584
rect 230532 152572 230538 152584
rect 233234 152572 233240 152584
rect 230532 152544 233240 152572
rect 230532 152532 230538 152544
rect 233234 152532 233240 152544
rect 233292 152532 233298 152584
rect 234154 152464 234160 152516
rect 234212 152504 234218 152516
rect 265710 152504 265716 152516
rect 234212 152476 265716 152504
rect 234212 152464 234218 152476
rect 265710 152464 265716 152476
rect 265768 152464 265774 152516
rect 211798 152396 211804 152448
rect 211856 152436 211862 152448
rect 213914 152436 213920 152448
rect 211856 152408 213920 152436
rect 211856 152396 211862 152408
rect 213914 152396 213920 152408
rect 213972 152396 213978 152448
rect 345106 152056 345112 152108
rect 345164 152096 345170 152108
rect 346578 152096 346584 152108
rect 345164 152068 346584 152096
rect 345164 152056 345170 152068
rect 346578 152056 346584 152068
rect 346636 152056 346642 152108
rect 189718 151852 189724 151904
rect 189776 151892 189782 151904
rect 214006 151892 214012 151904
rect 189776 151864 214012 151892
rect 189776 151852 189782 151864
rect 214006 151852 214012 151864
rect 214064 151852 214070 151904
rect 341610 151852 341616 151904
rect 341668 151892 341674 151904
rect 345106 151892 345112 151904
rect 341668 151864 345112 151892
rect 341668 151852 341674 151864
rect 345106 151852 345112 151864
rect 345164 151852 345170 151904
rect 180242 151784 180248 151836
rect 180300 151824 180306 151836
rect 213914 151824 213920 151836
rect 180300 151796 213920 151824
rect 180300 151784 180306 151796
rect 213914 151784 213920 151796
rect 213972 151784 213978 151836
rect 257522 151784 257528 151836
rect 257580 151824 257586 151836
rect 265802 151824 265808 151836
rect 257580 151796 265808 151824
rect 257580 151784 257586 151796
rect 265802 151784 265808 151796
rect 265860 151784 265866 151836
rect 231670 151716 231676 151768
rect 231728 151756 231734 151768
rect 252646 151756 252652 151768
rect 231728 151728 252652 151756
rect 231728 151716 231734 151728
rect 252646 151716 252652 151728
rect 252704 151716 252710 151768
rect 281902 151716 281908 151768
rect 281960 151756 281966 151768
rect 284386 151756 284392 151768
rect 281960 151728 284392 151756
rect 281960 151716 281966 151728
rect 284386 151716 284392 151728
rect 284444 151716 284450 151768
rect 342254 151716 342260 151768
rect 342312 151756 342318 151768
rect 346670 151756 346676 151768
rect 342312 151728 346676 151756
rect 342312 151716 342318 151728
rect 346670 151716 346676 151728
rect 346728 151716 346734 151768
rect 430574 151716 430580 151768
rect 430632 151756 430638 151768
rect 465718 151756 465724 151768
rect 430632 151728 465724 151756
rect 430632 151716 430638 151728
rect 465718 151716 465724 151728
rect 465776 151716 465782 151768
rect 231762 151648 231768 151700
rect 231820 151688 231826 151700
rect 249886 151688 249892 151700
rect 231820 151660 249892 151688
rect 231820 151648 231826 151660
rect 249886 151648 249892 151660
rect 249944 151648 249950 151700
rect 282270 151104 282276 151156
rect 282328 151144 282334 151156
rect 285858 151144 285864 151156
rect 282328 151116 285864 151144
rect 282328 151104 282334 151116
rect 285858 151104 285864 151116
rect 285916 151104 285922 151156
rect 332042 151036 332048 151088
rect 332100 151076 332106 151088
rect 342254 151076 342260 151088
rect 332100 151048 342260 151076
rect 332100 151036 332106 151048
rect 342254 151036 342260 151048
rect 342312 151036 342318 151088
rect 249150 150492 249156 150544
rect 249208 150532 249214 150544
rect 265802 150532 265808 150544
rect 249208 150504 265808 150532
rect 249208 150492 249214 150504
rect 265802 150492 265808 150504
rect 265860 150492 265866 150544
rect 235442 150424 235448 150476
rect 235500 150464 235506 150476
rect 265894 150464 265900 150476
rect 235500 150436 265900 150464
rect 235500 150424 235506 150436
rect 265894 150424 265900 150436
rect 265952 150424 265958 150476
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 22738 150396 22744 150408
rect 3476 150368 22744 150396
rect 3476 150356 3482 150368
rect 22738 150356 22744 150368
rect 22796 150356 22802 150408
rect 169018 150356 169024 150408
rect 169076 150396 169082 150408
rect 213914 150396 213920 150408
rect 169076 150368 213920 150396
rect 169076 150356 169082 150368
rect 213914 150356 213920 150368
rect 213972 150356 213978 150408
rect 231670 150356 231676 150408
rect 231728 150396 231734 150408
rect 259454 150396 259460 150408
rect 231728 150368 259460 150396
rect 231728 150356 231734 150368
rect 259454 150356 259460 150368
rect 259512 150356 259518 150408
rect 282730 150356 282736 150408
rect 282788 150396 282794 150408
rect 310514 150396 310520 150408
rect 282788 150368 310520 150396
rect 282788 150356 282794 150368
rect 310514 150356 310520 150368
rect 310572 150356 310578 150408
rect 430574 150356 430580 150408
rect 430632 150396 430638 150408
rect 437658 150396 437664 150408
rect 430632 150368 437664 150396
rect 430632 150356 430638 150368
rect 437658 150356 437664 150368
rect 437716 150356 437722 150408
rect 282822 150288 282828 150340
rect 282880 150328 282886 150340
rect 294230 150328 294236 150340
rect 282880 150300 294236 150328
rect 282880 150288 282886 150300
rect 294230 150288 294236 150300
rect 294288 150288 294294 150340
rect 430850 150288 430856 150340
rect 430908 150328 430914 150340
rect 436094 150328 436100 150340
rect 430908 150300 436100 150328
rect 430908 150288 430914 150300
rect 436094 150288 436100 150300
rect 436152 150288 436158 150340
rect 231762 149812 231768 149864
rect 231820 149852 231826 149864
rect 235994 149852 236000 149864
rect 231820 149824 236000 149852
rect 231820 149812 231826 149824
rect 235994 149812 236000 149824
rect 236052 149812 236058 149864
rect 235258 149676 235264 149728
rect 235316 149716 235322 149728
rect 265986 149716 265992 149728
rect 235316 149688 265992 149716
rect 235316 149676 235322 149688
rect 265986 149676 265992 149688
rect 266044 149676 266050 149728
rect 323578 149676 323584 149728
rect 323636 149716 323642 149728
rect 342254 149716 342260 149728
rect 323636 149688 342260 149716
rect 323636 149676 323642 149688
rect 342254 149676 342260 149688
rect 342312 149676 342318 149728
rect 249242 149132 249248 149184
rect 249300 149172 249306 149184
rect 265250 149172 265256 149184
rect 249300 149144 265256 149172
rect 249300 149132 249306 149144
rect 265250 149132 265256 149144
rect 265308 149132 265314 149184
rect 342254 149132 342260 149184
rect 342312 149172 342318 149184
rect 347498 149172 347504 149184
rect 342312 149144 347504 149172
rect 342312 149132 342318 149144
rect 347498 149132 347504 149144
rect 347556 149132 347562 149184
rect 239582 149064 239588 149116
rect 239640 149104 239646 149116
rect 265894 149104 265900 149116
rect 239640 149076 265900 149104
rect 239640 149064 239646 149076
rect 265894 149064 265900 149076
rect 265952 149064 265958 149116
rect 167638 148996 167644 149048
rect 167696 149036 167702 149048
rect 213914 149036 213920 149048
rect 167696 149008 213920 149036
rect 167696 148996 167702 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 282822 148996 282828 149048
rect 282880 149036 282886 149048
rect 296898 149036 296904 149048
rect 282880 149008 296904 149036
rect 282880 148996 282886 149008
rect 296898 148996 296904 149008
rect 296956 148996 296962 149048
rect 430574 148996 430580 149048
rect 430632 149036 430638 149048
rect 434898 149036 434904 149048
rect 430632 149008 434904 149036
rect 430632 148996 430638 149008
rect 434898 148996 434904 149008
rect 434956 148996 434962 149048
rect 231302 148928 231308 148980
rect 231360 148968 231366 148980
rect 234614 148968 234620 148980
rect 231360 148940 234620 148968
rect 231360 148928 231366 148940
rect 234614 148928 234620 148940
rect 234672 148928 234678 148980
rect 177482 148316 177488 148368
rect 177540 148356 177546 148368
rect 214006 148356 214012 148368
rect 177540 148328 214012 148356
rect 177540 148316 177546 148328
rect 214006 148316 214012 148328
rect 214064 148316 214070 148368
rect 256234 148316 256240 148368
rect 256292 148356 256298 148368
rect 265802 148356 265808 148368
rect 256292 148328 265808 148356
rect 256292 148316 256298 148328
rect 265802 148316 265808 148328
rect 265860 148316 265866 148368
rect 231210 147704 231216 147756
rect 231268 147744 231274 147756
rect 238018 147744 238024 147756
rect 231268 147716 238024 147744
rect 231268 147704 231274 147716
rect 238018 147704 238024 147716
rect 238076 147704 238082 147756
rect 246482 147704 246488 147756
rect 246540 147744 246546 147756
rect 265710 147744 265716 147756
rect 246540 147716 265716 147744
rect 246540 147704 246546 147716
rect 265710 147704 265716 147716
rect 265768 147704 265774 147756
rect 191190 147636 191196 147688
rect 191248 147676 191254 147688
rect 213914 147676 213920 147688
rect 191248 147648 213920 147676
rect 191248 147636 191254 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 236914 147636 236920 147688
rect 236972 147676 236978 147688
rect 265434 147676 265440 147688
rect 236972 147648 265440 147676
rect 236972 147636 236978 147648
rect 265434 147636 265440 147648
rect 265492 147636 265498 147688
rect 282822 147568 282828 147620
rect 282880 147608 282886 147620
rect 289906 147608 289912 147620
rect 282880 147580 289912 147608
rect 282880 147568 282886 147580
rect 289906 147568 289912 147580
rect 289964 147568 289970 147620
rect 335998 146956 336004 147008
rect 336056 146996 336062 147008
rect 338206 146996 338212 147008
rect 336056 146968 338212 146996
rect 336056 146956 336062 146968
rect 338206 146956 338212 146968
rect 338264 146996 338270 147008
rect 338264 146968 345014 146996
rect 338264 146956 338270 146968
rect 344986 146928 345014 146968
rect 346670 146928 346676 146940
rect 344986 146900 346676 146928
rect 346670 146888 346676 146900
rect 346728 146888 346734 146940
rect 167638 146276 167644 146328
rect 167696 146316 167702 146328
rect 213914 146316 213920 146328
rect 167696 146288 213920 146316
rect 167696 146276 167702 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 235534 146276 235540 146328
rect 235592 146316 235598 146328
rect 265710 146316 265716 146328
rect 235592 146288 265716 146316
rect 235592 146276 235598 146288
rect 265710 146276 265716 146288
rect 265768 146276 265774 146328
rect 282822 146208 282828 146260
rect 282880 146248 282886 146260
rect 311894 146248 311900 146260
rect 282880 146220 311900 146248
rect 282880 146208 282886 146220
rect 311894 146208 311900 146220
rect 311952 146208 311958 146260
rect 430574 146208 430580 146260
rect 430632 146248 430638 146260
rect 436278 146248 436284 146260
rect 430632 146220 436284 146248
rect 430632 146208 430638 146220
rect 436278 146208 436284 146220
rect 436336 146208 436342 146260
rect 231762 146140 231768 146192
rect 231820 146180 231826 146192
rect 247034 146180 247040 146192
rect 231820 146152 247040 146180
rect 231820 146140 231826 146152
rect 247034 146140 247040 146152
rect 247092 146140 247098 146192
rect 282730 146140 282736 146192
rect 282788 146180 282794 146192
rect 291194 146180 291200 146192
rect 282788 146152 291200 146180
rect 282788 146140 282794 146152
rect 291194 146140 291200 146152
rect 291252 146140 291258 146192
rect 231394 146072 231400 146124
rect 231452 146112 231458 146124
rect 256786 146112 256792 146124
rect 231452 146084 256792 146112
rect 231452 146072 231458 146084
rect 256786 146072 256792 146084
rect 256844 146072 256850 146124
rect 230842 146004 230848 146056
rect 230900 146044 230906 146056
rect 232682 146044 232688 146056
rect 230900 146016 232688 146044
rect 230900 146004 230906 146016
rect 232682 146004 232688 146016
rect 232740 146004 232746 146056
rect 232590 145528 232596 145580
rect 232648 145568 232654 145580
rect 265526 145568 265532 145580
rect 232648 145540 265532 145568
rect 232648 145528 232654 145540
rect 265526 145528 265532 145540
rect 265584 145528 265590 145580
rect 313918 145528 313924 145580
rect 313976 145568 313982 145580
rect 346670 145568 346676 145580
rect 313976 145540 346676 145568
rect 313976 145528 313982 145540
rect 346670 145528 346676 145540
rect 346728 145528 346734 145580
rect 232498 145052 232504 145104
rect 232556 145092 232562 145104
rect 265802 145092 265808 145104
rect 232556 145064 265808 145092
rect 232556 145052 232562 145064
rect 265802 145052 265808 145064
rect 265860 145052 265866 145104
rect 196802 144984 196808 145036
rect 196860 145024 196866 145036
rect 213914 145024 213920 145036
rect 196860 144996 213920 145024
rect 196860 144984 196866 144996
rect 213914 144984 213920 144996
rect 213972 144984 213978 145036
rect 242342 144984 242348 145036
rect 242400 145024 242406 145036
rect 265894 145024 265900 145036
rect 242400 144996 265900 145024
rect 242400 144984 242406 144996
rect 265894 144984 265900 144996
rect 265952 144984 265958 145036
rect 171778 144916 171784 144968
rect 171836 144956 171842 144968
rect 214006 144956 214012 144968
rect 171836 144928 214012 144956
rect 171836 144916 171842 144928
rect 214006 144916 214012 144928
rect 214064 144916 214070 144968
rect 282730 144848 282736 144900
rect 282788 144888 282794 144900
rect 311986 144888 311992 144900
rect 282788 144860 311992 144888
rect 282788 144848 282794 144860
rect 311986 144848 311992 144860
rect 312044 144848 312050 144900
rect 430574 144848 430580 144900
rect 430632 144888 430638 144900
rect 441706 144888 441712 144900
rect 430632 144860 441712 144888
rect 430632 144848 430638 144860
rect 441706 144848 441712 144860
rect 441764 144848 441770 144900
rect 282822 144780 282828 144832
rect 282880 144820 282886 144832
rect 298278 144820 298284 144832
rect 282880 144792 298284 144820
rect 282880 144780 282886 144792
rect 298278 144780 298284 144792
rect 298336 144780 298342 144832
rect 430850 144780 430856 144832
rect 430908 144820 430914 144832
rect 440418 144820 440424 144832
rect 430908 144792 440424 144820
rect 430908 144780 430914 144792
rect 440418 144780 440424 144792
rect 440476 144780 440482 144832
rect 300854 144168 300860 144220
rect 300912 144208 300918 144220
rect 346302 144208 346308 144220
rect 300912 144180 346308 144208
rect 300912 144168 300918 144180
rect 346302 144168 346308 144180
rect 346360 144168 346366 144220
rect 231762 143964 231768 144016
rect 231820 144004 231826 144016
rect 234798 144004 234804 144016
rect 231820 143976 234804 144004
rect 231820 143964 231826 143976
rect 234798 143964 234804 143976
rect 234856 143964 234862 144016
rect 264514 143692 264520 143744
rect 264572 143732 264578 143744
rect 266078 143732 266084 143744
rect 264572 143704 266084 143732
rect 264572 143692 264578 143704
rect 266078 143692 266084 143704
rect 266136 143692 266142 143744
rect 210418 143624 210424 143676
rect 210476 143664 210482 143676
rect 214006 143664 214012 143676
rect 210476 143636 214012 143664
rect 210476 143624 210482 143636
rect 214006 143624 214012 143636
rect 214064 143624 214070 143676
rect 253106 143624 253112 143676
rect 253164 143664 253170 143676
rect 265526 143664 265532 143676
rect 253164 143636 265532 143664
rect 253164 143624 253170 143636
rect 265526 143624 265532 143636
rect 265584 143624 265590 143676
rect 176010 143556 176016 143608
rect 176068 143596 176074 143608
rect 213914 143596 213920 143608
rect 176068 143568 213920 143596
rect 176068 143556 176074 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 235350 143556 235356 143608
rect 235408 143596 235414 143608
rect 265802 143596 265808 143608
rect 235408 143568 265808 143596
rect 235408 143556 235414 143568
rect 265802 143556 265808 143568
rect 265860 143556 265866 143608
rect 344922 143556 344928 143608
rect 344980 143596 344986 143608
rect 346670 143596 346676 143608
rect 344980 143568 346676 143596
rect 344980 143556 344986 143568
rect 346670 143556 346676 143568
rect 346728 143556 346734 143608
rect 231762 143488 231768 143540
rect 231820 143528 231826 143540
rect 253934 143528 253940 143540
rect 231820 143500 253940 143528
rect 231820 143488 231826 143500
rect 253934 143488 253940 143500
rect 253992 143488 253998 143540
rect 282086 143488 282092 143540
rect 282144 143528 282150 143540
rect 307754 143528 307760 143540
rect 282144 143500 307760 143528
rect 282144 143488 282150 143500
rect 307754 143488 307760 143500
rect 307812 143488 307818 143540
rect 233970 142876 233976 142928
rect 234028 142916 234034 142928
rect 265710 142916 265716 142928
rect 234028 142888 265716 142916
rect 234028 142876 234034 142888
rect 265710 142876 265716 142888
rect 265768 142876 265774 142928
rect 169018 142808 169024 142860
rect 169076 142848 169082 142860
rect 214098 142848 214104 142860
rect 169076 142820 214104 142848
rect 169076 142808 169082 142820
rect 214098 142808 214104 142820
rect 214156 142808 214162 142860
rect 230014 142808 230020 142860
rect 230072 142848 230078 142860
rect 264422 142848 264428 142860
rect 230072 142820 264428 142848
rect 230072 142808 230078 142820
rect 264422 142808 264428 142820
rect 264480 142808 264486 142860
rect 322198 142808 322204 142860
rect 322256 142848 322262 142860
rect 346578 142848 346584 142860
rect 322256 142820 346584 142848
rect 322256 142808 322262 142820
rect 346578 142808 346584 142820
rect 346636 142808 346642 142860
rect 282822 142468 282828 142520
rect 282880 142508 282886 142520
rect 287330 142508 287336 142520
rect 282880 142480 287336 142508
rect 282880 142468 282886 142480
rect 287330 142468 287336 142480
rect 287388 142468 287394 142520
rect 254670 142196 254676 142248
rect 254728 142236 254734 142248
rect 265526 142236 265532 142248
rect 254728 142208 265532 142236
rect 254728 142196 254734 142208
rect 265526 142196 265532 142208
rect 265584 142196 265590 142248
rect 195422 142128 195428 142180
rect 195480 142168 195486 142180
rect 213914 142168 213920 142180
rect 195480 142140 213920 142168
rect 195480 142128 195486 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 253474 142128 253480 142180
rect 253532 142168 253538 142180
rect 265618 142168 265624 142180
rect 253532 142140 265624 142168
rect 253532 142128 253538 142140
rect 265618 142128 265624 142140
rect 265676 142128 265682 142180
rect 430574 142128 430580 142180
rect 430632 142168 430638 142180
rect 436094 142168 436100 142180
rect 430632 142140 436100 142168
rect 430632 142128 430638 142140
rect 436094 142128 436100 142140
rect 436152 142128 436158 142180
rect 231486 142060 231492 142112
rect 231544 142100 231550 142112
rect 251174 142100 251180 142112
rect 231544 142072 251180 142100
rect 231544 142060 231550 142072
rect 251174 142060 251180 142072
rect 251232 142060 251238 142112
rect 282730 142060 282736 142112
rect 282788 142100 282794 142112
rect 296806 142100 296812 142112
rect 282788 142072 296812 142100
rect 282788 142060 282794 142072
rect 296806 142060 296812 142072
rect 296864 142060 296870 142112
rect 231762 141992 231768 142044
rect 231820 142032 231826 142044
rect 248598 142032 248604 142044
rect 231820 142004 248604 142032
rect 231820 141992 231826 142004
rect 248598 141992 248604 142004
rect 248656 141992 248662 142044
rect 300118 141380 300124 141432
rect 300176 141420 300182 141432
rect 343818 141420 343824 141432
rect 300176 141392 343824 141420
rect 300176 141380 300182 141392
rect 343818 141380 343824 141392
rect 343876 141420 343882 141432
rect 346486 141420 346492 141432
rect 343876 141392 346492 141420
rect 343876 141380 343882 141392
rect 346486 141380 346492 141392
rect 346544 141380 346550 141432
rect 282822 141312 282828 141364
rect 282880 141352 282886 141364
rect 287146 141352 287152 141364
rect 282880 141324 287152 141352
rect 282880 141312 282886 141324
rect 287146 141312 287152 141324
rect 287204 141312 287210 141364
rect 259178 140904 259184 140956
rect 259236 140944 259242 140956
rect 264606 140944 264612 140956
rect 259236 140916 264612 140944
rect 259236 140904 259242 140916
rect 264606 140904 264612 140916
rect 264664 140904 264670 140956
rect 206370 140836 206376 140888
rect 206428 140876 206434 140888
rect 213914 140876 213920 140888
rect 206428 140848 213920 140876
rect 206428 140836 206434 140848
rect 213914 140836 213920 140848
rect 213972 140836 213978 140888
rect 232682 140836 232688 140888
rect 232740 140876 232746 140888
rect 264422 140876 264428 140888
rect 232740 140848 264428 140876
rect 232740 140836 232746 140848
rect 264422 140836 264428 140848
rect 264480 140836 264486 140888
rect 171870 140768 171876 140820
rect 171928 140808 171934 140820
rect 214006 140808 214012 140820
rect 171928 140780 214012 140808
rect 171928 140768 171934 140780
rect 214006 140768 214012 140780
rect 214064 140768 214070 140820
rect 232774 140768 232780 140820
rect 232832 140808 232838 140820
rect 265802 140808 265808 140820
rect 232832 140780 265808 140808
rect 232832 140768 232838 140780
rect 265802 140768 265808 140780
rect 265860 140768 265866 140820
rect 282822 140700 282828 140752
rect 282880 140740 282886 140752
rect 309134 140740 309140 140752
rect 282880 140712 309140 140740
rect 282880 140700 282886 140712
rect 309134 140700 309140 140712
rect 309192 140700 309198 140752
rect 430574 140700 430580 140752
rect 430632 140740 430638 140752
rect 445754 140740 445760 140752
rect 430632 140712 445760 140740
rect 430632 140700 430638 140712
rect 445754 140700 445760 140712
rect 445812 140700 445818 140752
rect 178862 140020 178868 140072
rect 178920 140060 178926 140072
rect 214650 140060 214656 140072
rect 178920 140032 214656 140060
rect 178920 140020 178926 140032
rect 214650 140020 214656 140032
rect 214708 140020 214714 140072
rect 231394 140020 231400 140072
rect 231452 140060 231458 140072
rect 240962 140060 240968 140072
rect 231452 140032 240968 140060
rect 231452 140020 231458 140032
rect 240962 140020 240968 140032
rect 241020 140020 241026 140072
rect 241054 140020 241060 140072
rect 241112 140060 241118 140072
rect 265710 140060 265716 140072
rect 241112 140032 265716 140060
rect 241112 140020 241118 140032
rect 265710 140020 265716 140032
rect 265768 140020 265774 140072
rect 445754 140020 445760 140072
rect 445812 140060 445818 140072
rect 493318 140060 493324 140072
rect 445812 140032 493324 140060
rect 445812 140020 445818 140032
rect 493318 140020 493324 140032
rect 493376 140020 493382 140072
rect 265710 139884 265716 139936
rect 265768 139924 265774 139936
rect 266170 139924 266176 139936
rect 265768 139896 266176 139924
rect 265768 139884 265774 139896
rect 266170 139884 266176 139896
rect 266228 139884 266234 139936
rect 231302 139748 231308 139800
rect 231360 139788 231366 139800
rect 236178 139788 236184 139800
rect 231360 139760 236184 139788
rect 231360 139748 231366 139760
rect 236178 139748 236184 139760
rect 236236 139748 236242 139800
rect 257430 139476 257436 139528
rect 257488 139516 257494 139528
rect 265250 139516 265256 139528
rect 257488 139488 265256 139516
rect 257488 139476 257494 139488
rect 265250 139476 265256 139488
rect 265308 139476 265314 139528
rect 209130 139408 209136 139460
rect 209188 139448 209194 139460
rect 213914 139448 213920 139460
rect 209188 139420 213920 139448
rect 209188 139408 209194 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 229922 139408 229928 139460
rect 229980 139448 229986 139460
rect 265894 139448 265900 139460
rect 229980 139420 265900 139448
rect 229980 139408 229986 139420
rect 265894 139408 265900 139420
rect 265952 139408 265958 139460
rect 282730 139340 282736 139392
rect 282788 139380 282794 139392
rect 305178 139380 305184 139392
rect 282788 139352 305184 139380
rect 282788 139340 282794 139352
rect 305178 139340 305184 139352
rect 305236 139340 305242 139392
rect 461670 139340 461676 139392
rect 461728 139380 461734 139392
rect 580166 139380 580172 139392
rect 461728 139352 580172 139380
rect 461728 139340 461734 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 231302 139272 231308 139324
rect 231360 139312 231366 139324
rect 233326 139312 233332 139324
rect 231360 139284 233332 139312
rect 231360 139272 231366 139284
rect 233326 139272 233332 139284
rect 233384 139272 233390 139324
rect 282822 139272 282828 139324
rect 282880 139312 282886 139324
rect 299474 139312 299480 139324
rect 282880 139284 299480 139312
rect 282880 139272 282886 139284
rect 299474 139272 299480 139284
rect 299532 139272 299538 139324
rect 231762 139204 231768 139256
rect 231820 139244 231826 139256
rect 247126 139244 247132 139256
rect 231820 139216 247132 139244
rect 231820 139204 231826 139216
rect 247126 139204 247132 139216
rect 247184 139204 247190 139256
rect 231578 138660 231584 138712
rect 231636 138700 231642 138712
rect 242250 138700 242256 138712
rect 231636 138672 242256 138700
rect 231636 138660 231642 138672
rect 242250 138660 242256 138672
rect 242308 138660 242314 138712
rect 327718 138660 327724 138712
rect 327776 138700 327782 138712
rect 346394 138700 346400 138712
rect 327776 138672 346400 138700
rect 327776 138660 327782 138672
rect 346394 138660 346400 138672
rect 346452 138700 346458 138712
rect 347130 138700 347136 138712
rect 346452 138672 347136 138700
rect 346452 138660 346458 138672
rect 347130 138660 347136 138672
rect 347188 138660 347194 138712
rect 436738 138660 436744 138712
rect 436796 138700 436802 138712
rect 460934 138700 460940 138712
rect 436796 138672 460940 138700
rect 436796 138660 436802 138672
rect 460934 138660 460940 138672
rect 460992 138700 460998 138712
rect 461670 138700 461676 138712
rect 460992 138672 461676 138700
rect 460992 138660 460998 138672
rect 461670 138660 461676 138672
rect 461728 138660 461734 138712
rect 231486 138252 231492 138304
rect 231544 138292 231550 138304
rect 236086 138292 236092 138304
rect 231544 138264 236092 138292
rect 231544 138252 231550 138264
rect 236086 138252 236092 138264
rect 236144 138252 236150 138304
rect 247770 138116 247776 138168
rect 247828 138156 247834 138168
rect 264422 138156 264428 138168
rect 247828 138128 264428 138156
rect 247828 138116 247834 138128
rect 264422 138116 264428 138128
rect 264480 138116 264486 138168
rect 243630 138048 243636 138100
rect 243688 138088 243694 138100
rect 265158 138088 265164 138100
rect 243688 138060 265164 138088
rect 243688 138048 243694 138060
rect 265158 138048 265164 138060
rect 265216 138048 265222 138100
rect 238018 137980 238024 138032
rect 238076 138020 238082 138032
rect 265434 138020 265440 138032
rect 238076 137992 265440 138020
rect 238076 137980 238082 137992
rect 265434 137980 265440 137992
rect 265492 137980 265498 138032
rect 429746 137980 429752 138032
rect 429804 138020 429810 138032
rect 436646 138020 436652 138032
rect 429804 137992 436652 138020
rect 429804 137980 429810 137992
rect 436646 137980 436652 137992
rect 436704 137980 436710 138032
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 17218 137952 17224 137964
rect 3292 137924 17224 137952
rect 3292 137912 3298 137924
rect 17218 137912 17224 137924
rect 17276 137912 17282 137964
rect 231394 137912 231400 137964
rect 231452 137952 231458 137964
rect 258074 137952 258080 137964
rect 231452 137924 258080 137952
rect 231452 137912 231458 137924
rect 258074 137912 258080 137924
rect 258132 137912 258138 137964
rect 282822 137912 282828 137964
rect 282880 137952 282886 137964
rect 304994 137952 305000 137964
rect 282880 137924 305000 137952
rect 282880 137912 282886 137924
rect 304994 137912 305000 137924
rect 305052 137912 305058 137964
rect 430850 137912 430856 137964
rect 430908 137952 430914 137964
rect 436738 137952 436744 137964
rect 430908 137924 436744 137952
rect 430908 137912 430914 137924
rect 436738 137912 436744 137924
rect 436796 137912 436802 137964
rect 231762 137844 231768 137896
rect 231820 137884 231826 137896
rect 254026 137884 254032 137896
rect 231820 137856 254032 137884
rect 231820 137844 231826 137856
rect 254026 137844 254032 137856
rect 254084 137844 254090 137896
rect 282270 137776 282276 137828
rect 282328 137816 282334 137828
rect 285674 137816 285680 137828
rect 282328 137788 285680 137816
rect 282328 137776 282334 137788
rect 285674 137776 285680 137788
rect 285732 137776 285738 137828
rect 174630 137232 174636 137284
rect 174688 137272 174694 137284
rect 213914 137272 213920 137284
rect 174688 137244 213920 137272
rect 174688 137232 174694 137244
rect 213914 137232 213920 137244
rect 213972 137232 213978 137284
rect 234246 137232 234252 137284
rect 234304 137272 234310 137284
rect 265710 137272 265716 137284
rect 234304 137244 265716 137272
rect 234304 137232 234310 137244
rect 265710 137232 265716 137244
rect 265768 137232 265774 137284
rect 334710 137232 334716 137284
rect 334768 137272 334774 137284
rect 343726 137272 343732 137284
rect 334768 137244 343732 137272
rect 334768 137232 334774 137244
rect 343726 137232 343732 137244
rect 343784 137232 343790 137284
rect 430574 137232 430580 137284
rect 430632 137272 430638 137284
rect 430632 137244 431954 137272
rect 430632 137232 430638 137244
rect 431926 137204 431954 137244
rect 436646 137232 436652 137284
rect 436704 137272 436710 137284
rect 580258 137272 580264 137284
rect 436704 137244 580264 137272
rect 436704 137232 436710 137244
rect 580258 137232 580264 137244
rect 580316 137232 580322 137284
rect 436186 137204 436192 137216
rect 431926 137176 436192 137204
rect 436186 137164 436192 137176
rect 436244 137204 436250 137216
rect 436738 137204 436744 137216
rect 436244 137176 436744 137204
rect 436244 137164 436250 137176
rect 436738 137164 436744 137176
rect 436796 137164 436802 137216
rect 343726 136688 343732 136740
rect 343784 136728 343790 136740
rect 346670 136728 346676 136740
rect 343784 136700 346676 136728
rect 343784 136688 343790 136700
rect 346670 136688 346676 136700
rect 346728 136688 346734 136740
rect 229830 136620 229836 136672
rect 229888 136660 229894 136672
rect 264422 136660 264428 136672
rect 229888 136632 264428 136660
rect 229888 136620 229894 136632
rect 264422 136620 264428 136632
rect 264480 136620 264486 136672
rect 231394 136552 231400 136604
rect 231452 136592 231458 136604
rect 250438 136592 250444 136604
rect 231452 136564 250444 136592
rect 231452 136552 231458 136564
rect 250438 136552 250444 136564
rect 250496 136552 250502 136604
rect 282362 136552 282368 136604
rect 282420 136592 282426 136604
rect 306374 136592 306380 136604
rect 282420 136564 306380 136592
rect 282420 136552 282426 136564
rect 306374 136552 306380 136564
rect 306432 136552 306438 136604
rect 331858 136552 331864 136604
rect 331916 136592 331922 136604
rect 337378 136592 337384 136604
rect 331916 136564 337384 136592
rect 331916 136552 331922 136564
rect 337378 136552 337384 136564
rect 337436 136552 337442 136604
rect 430574 136552 430580 136604
rect 430632 136592 430638 136604
rect 431126 136592 431132 136604
rect 430632 136564 431132 136592
rect 430632 136552 430638 136564
rect 431126 136552 431132 136564
rect 431184 136592 431190 136604
rect 468478 136592 468484 136604
rect 431184 136564 468484 136592
rect 431184 136552 431190 136564
rect 468478 136552 468484 136564
rect 468536 136552 468542 136604
rect 230750 136484 230756 136536
rect 230808 136524 230814 136536
rect 246390 136524 246396 136536
rect 230808 136496 246396 136524
rect 230808 136484 230814 136496
rect 246390 136484 246396 136496
rect 246448 136484 246454 136536
rect 295978 135872 295984 135924
rect 296036 135912 296042 135924
rect 340966 135912 340972 135924
rect 296036 135884 340972 135912
rect 296036 135872 296042 135884
rect 340966 135872 340972 135884
rect 341024 135872 341030 135924
rect 261662 135464 261668 135516
rect 261720 135504 261726 135516
rect 265802 135504 265808 135516
rect 261720 135476 265808 135504
rect 261720 135464 261726 135476
rect 265802 135464 265808 135476
rect 265860 135464 265866 135516
rect 254762 135396 254768 135448
rect 254820 135436 254826 135448
rect 264422 135436 264428 135448
rect 254820 135408 264428 135436
rect 254820 135396 254826 135408
rect 264422 135396 264428 135408
rect 264480 135396 264486 135448
rect 184290 135328 184296 135380
rect 184348 135368 184354 135380
rect 213914 135368 213920 135380
rect 184348 135340 213920 135368
rect 184348 135328 184354 135340
rect 213914 135328 213920 135340
rect 213972 135328 213978 135380
rect 246574 135328 246580 135380
rect 246632 135368 246638 135380
rect 261110 135368 261116 135380
rect 246632 135340 261116 135368
rect 246632 135328 246638 135340
rect 261110 135328 261116 135340
rect 261168 135328 261174 135380
rect 173250 135260 173256 135312
rect 173308 135300 173314 135312
rect 214006 135300 214012 135312
rect 173308 135272 214012 135300
rect 173308 135260 173314 135272
rect 214006 135260 214012 135272
rect 214064 135260 214070 135312
rect 236638 135260 236644 135312
rect 236696 135300 236702 135312
rect 260926 135300 260932 135312
rect 236696 135272 260932 135300
rect 236696 135260 236702 135272
rect 260926 135260 260932 135272
rect 260984 135260 260990 135312
rect 340966 135260 340972 135312
rect 341024 135300 341030 135312
rect 347498 135300 347504 135312
rect 341024 135272 347504 135300
rect 341024 135260 341030 135272
rect 347498 135260 347504 135272
rect 347556 135260 347562 135312
rect 231762 135192 231768 135244
rect 231820 135232 231826 135244
rect 256050 135232 256056 135244
rect 231820 135204 256056 135232
rect 231820 135192 231826 135204
rect 256050 135192 256056 135204
rect 256108 135192 256114 135244
rect 282730 135192 282736 135244
rect 282788 135232 282794 135244
rect 300946 135232 300952 135244
rect 282788 135204 300952 135232
rect 282788 135192 282794 135204
rect 300946 135192 300952 135204
rect 301004 135192 301010 135244
rect 430574 135192 430580 135244
rect 430632 135232 430638 135244
rect 446398 135232 446404 135244
rect 430632 135204 446404 135232
rect 430632 135192 430638 135204
rect 446398 135192 446404 135204
rect 446456 135192 446462 135244
rect 231670 135124 231676 135176
rect 231728 135164 231734 135176
rect 244918 135164 244924 135176
rect 231728 135136 244924 135164
rect 231728 135124 231734 135136
rect 244918 135124 244924 135136
rect 244976 135124 244982 135176
rect 282822 135124 282828 135176
rect 282880 135164 282886 135176
rect 298186 135164 298192 135176
rect 282880 135136 298192 135164
rect 282880 135124 282886 135136
rect 298186 135124 298192 135136
rect 298244 135124 298250 135176
rect 230566 135056 230572 135108
rect 230624 135096 230630 135108
rect 239398 135096 239404 135108
rect 230624 135068 239404 135096
rect 230624 135056 230630 135068
rect 239398 135056 239404 135068
rect 239456 135056 239462 135108
rect 255958 134036 255964 134088
rect 256016 134076 256022 134088
rect 265710 134076 265716 134088
rect 256016 134048 265716 134076
rect 256016 134036 256022 134048
rect 265710 134036 265716 134048
rect 265768 134036 265774 134088
rect 245102 133968 245108 134020
rect 245160 134008 245166 134020
rect 265526 134008 265532 134020
rect 245160 133980 265532 134008
rect 245160 133968 245166 133980
rect 265526 133968 265532 133980
rect 265584 133968 265590 134020
rect 181438 133900 181444 133952
rect 181496 133940 181502 133952
rect 213914 133940 213920 133952
rect 181496 133912 213920 133940
rect 181496 133900 181502 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 236822 133900 236828 133952
rect 236880 133940 236886 133952
rect 265802 133940 265808 133952
rect 236880 133912 265808 133940
rect 236880 133900 236886 133912
rect 265802 133900 265808 133912
rect 265860 133900 265866 133952
rect 231762 133832 231768 133884
rect 231820 133872 231826 133884
rect 260098 133872 260104 133884
rect 231820 133844 260104 133872
rect 231820 133832 231826 133844
rect 260098 133832 260104 133844
rect 260156 133832 260162 133884
rect 281994 133832 282000 133884
rect 282052 133872 282058 133884
rect 310606 133872 310612 133884
rect 282052 133844 310612 133872
rect 282052 133832 282058 133844
rect 310606 133832 310612 133844
rect 310664 133832 310670 133884
rect 430574 133832 430580 133884
rect 430632 133872 430638 133884
rect 485038 133872 485044 133884
rect 430632 133844 485044 133872
rect 430632 133832 430638 133844
rect 485038 133832 485044 133844
rect 485096 133832 485102 133884
rect 231670 133764 231676 133816
rect 231728 133804 231734 133816
rect 243814 133804 243820 133816
rect 231728 133776 243820 133804
rect 231728 133764 231734 133776
rect 243814 133764 243820 133776
rect 243872 133764 243878 133816
rect 282178 133424 282184 133476
rect 282236 133464 282242 133476
rect 284294 133464 284300 133476
rect 282236 133436 284300 133464
rect 282236 133424 282242 133436
rect 284294 133424 284300 133436
rect 284352 133424 284358 133476
rect 259086 133152 259092 133204
rect 259144 133192 259150 133204
rect 265986 133192 265992 133204
rect 259144 133164 265992 133192
rect 259144 133152 259150 133164
rect 265986 133152 265992 133164
rect 266044 133152 266050 133204
rect 309778 133152 309784 133204
rect 309836 133192 309842 133204
rect 346578 133192 346584 133204
rect 309836 133164 346584 133192
rect 309836 133152 309842 133164
rect 346578 133152 346584 133164
rect 346636 133152 346642 133204
rect 180150 132540 180156 132592
rect 180208 132580 180214 132592
rect 214006 132580 214012 132592
rect 180208 132552 214012 132580
rect 180208 132540 180214 132552
rect 214006 132540 214012 132552
rect 214064 132540 214070 132592
rect 250438 132540 250444 132592
rect 250496 132580 250502 132592
rect 265894 132580 265900 132592
rect 250496 132552 265900 132580
rect 250496 132540 250502 132552
rect 265894 132540 265900 132552
rect 265952 132540 265958 132592
rect 170582 132472 170588 132524
rect 170640 132512 170646 132524
rect 213914 132512 213920 132524
rect 170640 132484 213920 132512
rect 170640 132472 170646 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 243538 132472 243544 132524
rect 243596 132512 243602 132524
rect 265710 132512 265716 132524
rect 243596 132484 265716 132512
rect 243596 132472 243602 132484
rect 265710 132472 265716 132484
rect 265768 132472 265774 132524
rect 231670 132404 231676 132456
rect 231728 132444 231734 132456
rect 258994 132444 259000 132456
rect 231728 132416 259000 132444
rect 231728 132404 231734 132416
rect 258994 132404 259000 132416
rect 259052 132404 259058 132456
rect 282822 132404 282828 132456
rect 282880 132444 282886 132456
rect 314654 132444 314660 132456
rect 282880 132416 314660 132444
rect 282880 132404 282886 132416
rect 314654 132404 314660 132416
rect 314712 132404 314718 132456
rect 430574 132404 430580 132456
rect 430632 132444 430638 132456
rect 452654 132444 452660 132456
rect 430632 132416 452660 132444
rect 430632 132404 430638 132416
rect 452654 132404 452660 132416
rect 452712 132404 452718 132456
rect 230658 132336 230664 132388
rect 230716 132376 230722 132388
rect 258718 132376 258724 132388
rect 230716 132348 258724 132376
rect 230716 132336 230722 132348
rect 258718 132336 258724 132348
rect 258776 132336 258782 132388
rect 430850 132336 430856 132388
rect 430908 132376 430914 132388
rect 440234 132376 440240 132388
rect 430908 132348 440240 132376
rect 430908 132336 430914 132348
rect 440234 132336 440240 132348
rect 440292 132336 440298 132388
rect 231762 132268 231768 132320
rect 231820 132308 231826 132320
rect 250530 132308 250536 132320
rect 231820 132280 250536 132308
rect 231820 132268 231826 132280
rect 250530 132268 250536 132280
rect 250588 132268 250594 132320
rect 320818 131724 320824 131776
rect 320876 131764 320882 131776
rect 345198 131764 345204 131776
rect 320876 131736 345204 131764
rect 320876 131724 320882 131736
rect 345198 131724 345204 131736
rect 345256 131764 345262 131776
rect 347406 131764 347412 131776
rect 345256 131736 347412 131764
rect 345256 131724 345262 131736
rect 347406 131724 347412 131736
rect 347464 131724 347470 131776
rect 282270 131316 282276 131368
rect 282328 131356 282334 131368
rect 288618 131356 288624 131368
rect 282328 131328 288624 131356
rect 282328 131316 282334 131328
rect 288618 131316 288624 131328
rect 288676 131316 288682 131368
rect 258810 131248 258816 131300
rect 258868 131288 258874 131300
rect 265710 131288 265716 131300
rect 258868 131260 265716 131288
rect 258868 131248 258874 131260
rect 265710 131248 265716 131260
rect 265768 131248 265774 131300
rect 258902 131180 258908 131232
rect 258960 131220 258966 131232
rect 265434 131220 265440 131232
rect 258960 131192 265440 131220
rect 258960 131180 258966 131192
rect 265434 131180 265440 131192
rect 265492 131180 265498 131232
rect 193858 131112 193864 131164
rect 193916 131152 193922 131164
rect 213914 131152 213920 131164
rect 193916 131124 213920 131152
rect 193916 131112 193922 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 253382 131112 253388 131164
rect 253440 131152 253446 131164
rect 265894 131152 265900 131164
rect 253440 131124 265900 131152
rect 253440 131112 253446 131124
rect 265894 131112 265900 131124
rect 265952 131112 265958 131164
rect 231762 131044 231768 131096
rect 231820 131084 231826 131096
rect 251910 131084 251916 131096
rect 231820 131056 251916 131084
rect 231820 131044 231826 131056
rect 251910 131044 251916 131056
rect 251968 131044 251974 131096
rect 231394 130976 231400 131028
rect 231452 131016 231458 131028
rect 242158 131016 242164 131028
rect 231452 130988 242164 131016
rect 231452 130976 231458 130988
rect 242158 130976 242164 130988
rect 242216 130976 242222 131028
rect 231578 130364 231584 130416
rect 231636 130404 231642 130416
rect 263134 130404 263140 130416
rect 231636 130376 263140 130404
rect 231636 130364 231642 130376
rect 263134 130364 263140 130376
rect 263192 130364 263198 130416
rect 281626 129820 281632 129872
rect 281684 129860 281690 129872
rect 288434 129860 288440 129872
rect 281684 129832 288440 129860
rect 281684 129820 281690 129832
rect 288434 129820 288440 129832
rect 288492 129820 288498 129872
rect 251818 129752 251824 129804
rect 251876 129792 251882 129804
rect 265250 129792 265256 129804
rect 251876 129764 265256 129792
rect 251876 129752 251882 129764
rect 265250 129752 265256 129764
rect 265308 129752 265314 129804
rect 231762 129684 231768 129736
rect 231820 129724 231826 129736
rect 247862 129724 247868 129736
rect 231820 129696 247868 129724
rect 231820 129684 231826 129696
rect 247862 129684 247868 129696
rect 247920 129684 247926 129736
rect 282822 129684 282828 129736
rect 282880 129724 282886 129736
rect 309318 129724 309324 129736
rect 282880 129696 309324 129724
rect 282880 129684 282886 129696
rect 309318 129684 309324 129696
rect 309376 129684 309382 129736
rect 430574 129684 430580 129736
rect 430632 129724 430638 129736
rect 444374 129724 444380 129736
rect 430632 129696 444380 129724
rect 430632 129684 430638 129696
rect 444374 129684 444380 129696
rect 444432 129684 444438 129736
rect 231394 129616 231400 129668
rect 231452 129656 231458 129668
rect 246666 129656 246672 129668
rect 231452 129628 246672 129656
rect 231452 129616 231458 129628
rect 246666 129616 246672 129628
rect 246724 129616 246730 129668
rect 207658 128392 207664 128444
rect 207716 128432 207722 128444
rect 213914 128432 213920 128444
rect 207716 128404 213920 128432
rect 207716 128392 207722 128404
rect 213914 128392 213920 128404
rect 213972 128392 213978 128444
rect 247678 128392 247684 128444
rect 247736 128432 247742 128444
rect 264422 128432 264428 128444
rect 247736 128404 264428 128432
rect 247736 128392 247742 128404
rect 264422 128392 264428 128404
rect 264480 128392 264486 128444
rect 173158 128324 173164 128376
rect 173216 128364 173222 128376
rect 214006 128364 214012 128376
rect 173216 128336 214012 128364
rect 173216 128324 173222 128336
rect 214006 128324 214012 128336
rect 214064 128324 214070 128376
rect 246390 128324 246396 128376
rect 246448 128364 246454 128376
rect 265710 128364 265716 128376
rect 246448 128336 265716 128364
rect 246448 128324 246454 128336
rect 265710 128324 265716 128336
rect 265768 128324 265774 128376
rect 231670 128256 231676 128308
rect 231728 128296 231734 128308
rect 249058 128296 249064 128308
rect 231728 128268 249064 128296
rect 231728 128256 231734 128268
rect 249058 128256 249064 128268
rect 249116 128256 249122 128308
rect 281626 128256 281632 128308
rect 281684 128296 281690 128308
rect 307846 128296 307852 128308
rect 281684 128268 307852 128296
rect 281684 128256 281690 128268
rect 307846 128256 307852 128268
rect 307904 128256 307910 128308
rect 312538 128256 312544 128308
rect 312596 128296 312602 128308
rect 347958 128296 347964 128308
rect 312596 128268 347964 128296
rect 312596 128256 312602 128268
rect 347958 128256 347964 128268
rect 348016 128256 348022 128308
rect 231762 128188 231768 128240
rect 231820 128228 231826 128240
rect 243722 128228 243728 128240
rect 231820 128200 243728 128228
rect 231820 128188 231826 128200
rect 243722 128188 243728 128200
rect 243780 128188 243786 128240
rect 231486 127576 231492 127628
rect 231544 127616 231550 127628
rect 252094 127616 252100 127628
rect 231544 127588 252100 127616
rect 231544 127576 231550 127588
rect 252094 127576 252100 127588
rect 252152 127576 252158 127628
rect 287054 127576 287060 127628
rect 287112 127616 287118 127628
rect 345106 127616 345112 127628
rect 287112 127588 345112 127616
rect 287112 127576 287118 127588
rect 345106 127576 345112 127588
rect 345164 127576 345170 127628
rect 282270 127440 282276 127492
rect 282328 127480 282334 127492
rect 285766 127480 285772 127492
rect 282328 127452 285772 127480
rect 282328 127440 282334 127452
rect 285766 127440 285772 127452
rect 285824 127440 285830 127492
rect 252002 127032 252008 127084
rect 252060 127072 252066 127084
rect 265894 127072 265900 127084
rect 252060 127044 265900 127072
rect 252060 127032 252066 127044
rect 265894 127032 265900 127044
rect 265952 127032 265958 127084
rect 250530 126964 250536 127016
rect 250588 127004 250594 127016
rect 264422 127004 264428 127016
rect 250588 126976 264428 127004
rect 250588 126964 250594 126976
rect 264422 126964 264428 126976
rect 264480 126964 264486 127016
rect 231670 126896 231676 126948
rect 231728 126936 231734 126948
rect 253198 126936 253204 126948
rect 231728 126908 253204 126936
rect 231728 126896 231734 126908
rect 253198 126896 253204 126908
rect 253256 126896 253262 126948
rect 282822 126896 282828 126948
rect 282880 126936 282886 126948
rect 301038 126936 301044 126948
rect 282880 126908 301044 126936
rect 282880 126896 282886 126908
rect 301038 126896 301044 126908
rect 301096 126896 301102 126948
rect 323670 126896 323676 126948
rect 323728 126936 323734 126948
rect 347682 126936 347688 126948
rect 323728 126908 347688 126936
rect 323728 126896 323734 126908
rect 347682 126896 347688 126908
rect 347740 126896 347746 126948
rect 447778 126896 447784 126948
rect 447836 126936 447842 126948
rect 580166 126936 580172 126948
rect 447836 126908 580172 126936
rect 447836 126896 447842 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 231762 126828 231768 126880
rect 231820 126868 231826 126880
rect 245010 126868 245016 126880
rect 231820 126840 245016 126868
rect 231820 126828 231826 126840
rect 245010 126828 245016 126840
rect 245068 126828 245074 126880
rect 305638 126216 305644 126268
rect 305696 126256 305702 126268
rect 347682 126256 347688 126268
rect 305696 126228 347688 126256
rect 305696 126216 305702 126228
rect 347682 126216 347688 126228
rect 347740 126216 347746 126268
rect 180334 125672 180340 125724
rect 180392 125712 180398 125724
rect 214006 125712 214012 125724
rect 180392 125684 214012 125712
rect 180392 125672 180398 125684
rect 214006 125672 214012 125684
rect 214064 125672 214070 125724
rect 59262 125604 59268 125656
rect 59320 125644 59326 125656
rect 65150 125644 65156 125656
rect 59320 125616 65156 125644
rect 59320 125604 59326 125616
rect 65150 125604 65156 125616
rect 65208 125604 65214 125656
rect 176102 125604 176108 125656
rect 176160 125644 176166 125656
rect 213914 125644 213920 125656
rect 176160 125616 213920 125644
rect 176160 125604 176166 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 254854 125604 254860 125656
rect 254912 125644 254918 125656
rect 265894 125644 265900 125656
rect 254912 125616 265900 125644
rect 254912 125604 254918 125616
rect 265894 125604 265900 125616
rect 265952 125604 265958 125656
rect 231302 125536 231308 125588
rect 231360 125576 231366 125588
rect 264238 125576 264244 125588
rect 231360 125548 264244 125576
rect 231360 125536 231366 125548
rect 264238 125536 264244 125548
rect 264296 125536 264302 125588
rect 282822 125536 282828 125588
rect 282880 125576 282886 125588
rect 292574 125576 292580 125588
rect 282880 125548 292580 125576
rect 282880 125536 282886 125548
rect 292574 125536 292580 125548
rect 292632 125536 292638 125588
rect 430574 125536 430580 125588
rect 430632 125576 430638 125588
rect 439038 125576 439044 125588
rect 430632 125548 439044 125576
rect 430632 125536 430638 125548
rect 439038 125536 439044 125548
rect 439096 125536 439102 125588
rect 231670 125468 231676 125520
rect 231728 125508 231734 125520
rect 263042 125508 263048 125520
rect 231728 125480 263048 125508
rect 231728 125468 231734 125480
rect 263042 125468 263048 125480
rect 263100 125468 263106 125520
rect 311894 124856 311900 124908
rect 311952 124896 311958 124908
rect 343818 124896 343824 124908
rect 311952 124868 343824 124896
rect 311952 124856 311958 124868
rect 343818 124856 343824 124868
rect 343876 124856 343882 124908
rect 170674 124244 170680 124296
rect 170732 124284 170738 124296
rect 213914 124284 213920 124296
rect 170732 124256 213920 124284
rect 170732 124244 170738 124256
rect 213914 124244 213920 124256
rect 213972 124244 213978 124296
rect 264606 124244 264612 124296
rect 264664 124284 264670 124296
rect 265618 124284 265624 124296
rect 264664 124256 265624 124284
rect 264664 124244 264670 124256
rect 265618 124244 265624 124256
rect 265676 124244 265682 124296
rect 169110 124176 169116 124228
rect 169168 124216 169174 124228
rect 214006 124216 214012 124228
rect 169168 124188 214012 124216
rect 169168 124176 169174 124188
rect 214006 124176 214012 124188
rect 214064 124176 214070 124228
rect 242158 124176 242164 124228
rect 242216 124216 242222 124228
rect 265894 124216 265900 124228
rect 242216 124188 265900 124216
rect 242216 124176 242222 124188
rect 265894 124176 265900 124188
rect 265952 124176 265958 124228
rect 231486 124108 231492 124160
rect 231544 124148 231550 124160
rect 260190 124148 260196 124160
rect 231544 124120 260196 124148
rect 231544 124108 231550 124120
rect 260190 124108 260196 124120
rect 260248 124108 260254 124160
rect 338758 124108 338764 124160
rect 338816 124148 338822 124160
rect 348970 124148 348976 124160
rect 338816 124120 348976 124148
rect 338816 124108 338822 124120
rect 348970 124108 348976 124120
rect 349028 124108 349034 124160
rect 430574 124108 430580 124160
rect 430632 124148 430638 124160
rect 443178 124148 443184 124160
rect 430632 124120 443184 124148
rect 430632 124108 430638 124120
rect 443178 124108 443184 124120
rect 443236 124108 443242 124160
rect 231302 124040 231308 124092
rect 231360 124080 231366 124092
rect 250622 124080 250628 124092
rect 231360 124052 250628 124080
rect 231360 124040 231366 124052
rect 250622 124040 250628 124052
rect 250680 124040 250686 124092
rect 231302 123428 231308 123480
rect 231360 123468 231366 123480
rect 257338 123468 257344 123480
rect 231360 123440 257344 123468
rect 231360 123428 231366 123440
rect 257338 123428 257344 123440
rect 257396 123428 257402 123480
rect 325694 123428 325700 123480
rect 325752 123468 325758 123480
rect 338298 123468 338304 123480
rect 325752 123440 338304 123468
rect 325752 123428 325758 123440
rect 338298 123428 338304 123440
rect 338356 123428 338362 123480
rect 261478 123088 261484 123140
rect 261536 123128 261542 123140
rect 265894 123128 265900 123140
rect 261536 123100 265900 123128
rect 261536 123088 261542 123100
rect 265894 123088 265900 123100
rect 265952 123088 265958 123140
rect 177390 122884 177396 122936
rect 177448 122924 177454 122936
rect 214006 122924 214012 122936
rect 177448 122896 214012 122924
rect 177448 122884 177454 122896
rect 214006 122884 214012 122896
rect 214064 122884 214070 122936
rect 260098 122884 260104 122936
rect 260156 122924 260162 122936
rect 265894 122924 265900 122936
rect 260156 122896 265900 122924
rect 260156 122884 260162 122896
rect 265894 122884 265900 122896
rect 265952 122884 265958 122936
rect 167822 122816 167828 122868
rect 167880 122856 167886 122868
rect 213914 122856 213920 122868
rect 167880 122828 213920 122856
rect 167880 122816 167886 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 256142 122816 256148 122868
rect 256200 122856 256206 122868
rect 265986 122856 265992 122868
rect 256200 122828 265992 122856
rect 256200 122816 256206 122828
rect 265986 122816 265992 122828
rect 266044 122816 266050 122868
rect 231762 122748 231768 122800
rect 231820 122788 231826 122800
rect 256326 122788 256332 122800
rect 231820 122760 256332 122788
rect 231820 122748 231826 122760
rect 256326 122748 256332 122760
rect 256384 122748 256390 122800
rect 430574 122748 430580 122800
rect 430632 122788 430638 122800
rect 449894 122788 449900 122800
rect 430632 122760 449900 122788
rect 430632 122748 430638 122760
rect 449894 122748 449900 122760
rect 449952 122748 449958 122800
rect 231486 122680 231492 122732
rect 231544 122720 231550 122732
rect 246298 122720 246304 122732
rect 231544 122692 246304 122720
rect 231544 122680 231550 122692
rect 246298 122680 246304 122692
rect 246356 122680 246362 122732
rect 282822 122680 282828 122732
rect 282880 122720 282886 122732
rect 303706 122720 303712 122732
rect 282880 122692 303712 122720
rect 282880 122680 282886 122692
rect 303706 122680 303712 122692
rect 303764 122680 303770 122732
rect 231578 122612 231584 122664
rect 231636 122652 231642 122664
rect 234062 122652 234068 122664
rect 231636 122624 234068 122652
rect 231636 122612 231642 122624
rect 234062 122612 234068 122624
rect 234120 122612 234126 122664
rect 257338 121592 257344 121644
rect 257396 121632 257402 121644
rect 264238 121632 264244 121644
rect 257396 121604 264244 121632
rect 257396 121592 257402 121604
rect 264238 121592 264244 121604
rect 264296 121592 264302 121644
rect 172054 121524 172060 121576
rect 172112 121564 172118 121576
rect 213914 121564 213920 121576
rect 172112 121536 213920 121564
rect 172112 121524 172118 121536
rect 213914 121524 213920 121536
rect 213972 121524 213978 121576
rect 249058 121524 249064 121576
rect 249116 121564 249122 121576
rect 265986 121564 265992 121576
rect 249116 121536 265992 121564
rect 249116 121524 249122 121536
rect 265986 121524 265992 121536
rect 266044 121524 266050 121576
rect 170490 121456 170496 121508
rect 170548 121496 170554 121508
rect 214006 121496 214012 121508
rect 170548 121468 214012 121496
rect 170548 121456 170554 121468
rect 214006 121456 214012 121468
rect 214064 121456 214070 121508
rect 233878 121456 233884 121508
rect 233936 121496 233942 121508
rect 265894 121496 265900 121508
rect 233936 121468 265900 121496
rect 233936 121456 233942 121468
rect 265894 121456 265900 121468
rect 265952 121456 265958 121508
rect 231762 121388 231768 121440
rect 231820 121428 231826 121440
rect 253290 121428 253296 121440
rect 231820 121400 253296 121428
rect 231820 121388 231826 121400
rect 253290 121388 253296 121400
rect 253348 121388 253354 121440
rect 281902 121388 281908 121440
rect 281960 121428 281966 121440
rect 309226 121428 309232 121440
rect 281960 121400 309232 121428
rect 281960 121388 281966 121400
rect 309226 121388 309232 121400
rect 309284 121388 309290 121440
rect 430574 121388 430580 121440
rect 430632 121428 430638 121440
rect 437566 121428 437572 121440
rect 430632 121400 437572 121428
rect 430632 121388 430638 121400
rect 437566 121388 437572 121400
rect 437624 121388 437630 121440
rect 231486 121320 231492 121372
rect 231544 121360 231550 121372
rect 240778 121360 240784 121372
rect 231544 121332 240784 121360
rect 231544 121320 231550 121332
rect 240778 121320 240784 121332
rect 240836 121320 240842 121372
rect 281626 121320 281632 121372
rect 281684 121360 281690 121372
rect 303614 121360 303620 121372
rect 281684 121332 303620 121360
rect 281684 121320 281690 121332
rect 303614 121320 303620 121332
rect 303672 121320 303678 121372
rect 231118 120912 231124 120964
rect 231176 120952 231182 120964
rect 238110 120952 238116 120964
rect 231176 120924 238116 120952
rect 231176 120912 231182 120924
rect 238110 120912 238116 120924
rect 238168 120912 238174 120964
rect 430574 120844 430580 120896
rect 430632 120884 430638 120896
rect 433334 120884 433340 120896
rect 430632 120856 433340 120884
rect 430632 120844 430638 120856
rect 433334 120844 433340 120856
rect 433392 120844 433398 120896
rect 170398 120708 170404 120760
rect 170456 120748 170462 120760
rect 203518 120748 203524 120760
rect 170456 120720 203524 120748
rect 170456 120708 170462 120720
rect 203518 120708 203524 120720
rect 203576 120708 203582 120760
rect 260190 120232 260196 120284
rect 260248 120272 260254 120284
rect 265526 120272 265532 120284
rect 260248 120244 265532 120272
rect 260248 120232 260254 120244
rect 265526 120232 265532 120244
rect 265584 120232 265590 120284
rect 178770 120164 178776 120216
rect 178828 120204 178834 120216
rect 214006 120204 214012 120216
rect 178828 120176 214012 120204
rect 178828 120164 178834 120176
rect 214006 120164 214012 120176
rect 214064 120164 214070 120216
rect 253198 120164 253204 120216
rect 253256 120204 253262 120216
rect 265710 120204 265716 120216
rect 253256 120176 265716 120204
rect 253256 120164 253262 120176
rect 265710 120164 265716 120176
rect 265768 120164 265774 120216
rect 173434 120096 173440 120148
rect 173492 120136 173498 120148
rect 213914 120136 213920 120148
rect 173492 120108 213920 120136
rect 173492 120096 173498 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 239398 120096 239404 120148
rect 239456 120136 239462 120148
rect 265618 120136 265624 120148
rect 239456 120108 265624 120136
rect 239456 120096 239462 120108
rect 265618 120096 265624 120108
rect 265676 120096 265682 120148
rect 231762 120028 231768 120080
rect 231820 120068 231826 120080
rect 261570 120068 261576 120080
rect 231820 120040 261576 120068
rect 231820 120028 231826 120040
rect 261570 120028 261576 120040
rect 261628 120028 261634 120080
rect 282086 120028 282092 120080
rect 282144 120068 282150 120080
rect 294138 120068 294144 120080
rect 282144 120040 294144 120068
rect 282144 120028 282150 120040
rect 294138 120028 294144 120040
rect 294196 120028 294202 120080
rect 315298 120028 315304 120080
rect 315356 120068 315362 120080
rect 347038 120068 347044 120080
rect 315356 120040 347044 120068
rect 315356 120028 315362 120040
rect 347038 120028 347044 120040
rect 347096 120028 347102 120080
rect 231394 119960 231400 120012
rect 231452 120000 231458 120012
rect 239490 120000 239496 120012
rect 231452 119972 239496 120000
rect 231452 119960 231458 119972
rect 239490 119960 239496 119972
rect 239548 119960 239554 120012
rect 430574 119892 430580 119944
rect 430632 119932 430638 119944
rect 433518 119932 433524 119944
rect 430632 119904 433524 119932
rect 430632 119892 430638 119904
rect 433518 119892 433524 119904
rect 433576 119892 433582 119944
rect 231302 119348 231308 119400
rect 231360 119388 231366 119400
rect 259178 119388 259184 119400
rect 231360 119360 259184 119388
rect 231360 119348 231366 119360
rect 259178 119348 259184 119360
rect 259236 119348 259242 119400
rect 210510 118804 210516 118856
rect 210568 118844 210574 118856
rect 214098 118844 214104 118856
rect 210568 118816 214104 118844
rect 210568 118804 210574 118816
rect 214098 118804 214104 118816
rect 214156 118804 214162 118856
rect 185578 118736 185584 118788
rect 185636 118776 185642 118788
rect 213914 118776 213920 118788
rect 185636 118748 213920 118776
rect 185636 118736 185642 118748
rect 213914 118736 213920 118748
rect 213972 118736 213978 118788
rect 258718 118736 258724 118788
rect 258776 118776 258782 118788
rect 265710 118776 265716 118788
rect 258776 118748 265716 118776
rect 258776 118736 258782 118748
rect 265710 118736 265716 118748
rect 265768 118736 265774 118788
rect 178954 118668 178960 118720
rect 179012 118708 179018 118720
rect 214006 118708 214012 118720
rect 179012 118680 214012 118708
rect 179012 118668 179018 118680
rect 214006 118668 214012 118680
rect 214064 118668 214070 118720
rect 246298 118668 246304 118720
rect 246356 118708 246362 118720
rect 265618 118708 265624 118720
rect 246356 118680 265624 118708
rect 246356 118668 246362 118680
rect 265618 118668 265624 118680
rect 265676 118668 265682 118720
rect 231486 118600 231492 118652
rect 231544 118640 231550 118652
rect 245286 118640 245292 118652
rect 231544 118612 245292 118640
rect 231544 118600 231550 118612
rect 245286 118600 245292 118612
rect 245344 118600 245350 118652
rect 282454 118600 282460 118652
rect 282512 118640 282518 118652
rect 305086 118640 305092 118652
rect 282512 118612 305092 118640
rect 282512 118600 282518 118612
rect 305086 118600 305092 118612
rect 305144 118600 305150 118652
rect 231762 118532 231768 118584
rect 231820 118572 231826 118584
rect 245194 118572 245200 118584
rect 231820 118544 245200 118572
rect 231820 118532 231826 118544
rect 245194 118532 245200 118544
rect 245252 118532 245258 118584
rect 231118 118464 231124 118516
rect 231176 118504 231182 118516
rect 239674 118504 239680 118516
rect 231176 118476 239680 118504
rect 231176 118464 231182 118476
rect 239674 118464 239680 118476
rect 239732 118464 239738 118516
rect 430574 118396 430580 118448
rect 430632 118436 430638 118448
rect 432230 118436 432236 118448
rect 430632 118408 432236 118436
rect 430632 118396 430638 118408
rect 432230 118396 432236 118408
rect 432288 118396 432294 118448
rect 282822 117988 282828 118040
rect 282880 118028 282886 118040
rect 287238 118028 287244 118040
rect 282880 118000 287244 118028
rect 282880 117988 282886 118000
rect 287238 117988 287244 118000
rect 287296 117988 287302 118040
rect 318794 117920 318800 117972
rect 318852 117960 318858 117972
rect 343726 117960 343732 117972
rect 318852 117932 343732 117960
rect 318852 117920 318858 117932
rect 343726 117920 343732 117932
rect 343784 117920 343790 117972
rect 244918 117444 244924 117496
rect 244976 117484 244982 117496
rect 265986 117484 265992 117496
rect 244976 117456 265992 117484
rect 244976 117444 244982 117456
rect 265986 117444 265992 117456
rect 266044 117444 266050 117496
rect 177574 117376 177580 117428
rect 177632 117416 177638 117428
rect 213914 117416 213920 117428
rect 177632 117388 213920 117416
rect 177632 117376 177638 117388
rect 213914 117376 213920 117388
rect 213972 117376 213978 117428
rect 245010 117376 245016 117428
rect 245068 117416 245074 117428
rect 265710 117416 265716 117428
rect 245068 117388 265716 117416
rect 245068 117376 245074 117388
rect 265710 117376 265716 117388
rect 265768 117376 265774 117428
rect 166350 117308 166356 117360
rect 166408 117348 166414 117360
rect 214006 117348 214012 117360
rect 166408 117320 214012 117348
rect 166408 117308 166414 117320
rect 214006 117308 214012 117320
rect 214064 117308 214070 117360
rect 239490 117308 239496 117360
rect 239548 117348 239554 117360
rect 265342 117348 265348 117360
rect 239548 117320 265348 117348
rect 239548 117308 239554 117320
rect 265342 117308 265348 117320
rect 265400 117308 265406 117360
rect 231486 117240 231492 117292
rect 231544 117280 231550 117292
rect 242434 117280 242440 117292
rect 231544 117252 242440 117280
rect 231544 117240 231550 117252
rect 242434 117240 242440 117252
rect 242492 117240 242498 117292
rect 282546 117240 282552 117292
rect 282604 117280 282610 117292
rect 302234 117280 302240 117292
rect 282604 117252 302240 117280
rect 282604 117240 282610 117252
rect 302234 117240 302240 117252
rect 302292 117240 302298 117292
rect 430574 117240 430580 117292
rect 430632 117280 430638 117292
rect 448606 117280 448612 117292
rect 430632 117252 448612 117280
rect 430632 117240 430638 117252
rect 448606 117240 448612 117252
rect 448664 117240 448670 117292
rect 231210 116764 231216 116816
rect 231268 116804 231274 116816
rect 238294 116804 238300 116816
rect 231268 116776 238300 116804
rect 231268 116764 231274 116776
rect 238294 116764 238300 116776
rect 238352 116764 238358 116816
rect 231118 116560 231124 116612
rect 231176 116600 231182 116612
rect 241146 116600 241152 116612
rect 231176 116572 241152 116600
rect 231176 116560 231182 116572
rect 241146 116560 241152 116572
rect 241204 116560 241210 116612
rect 323026 116560 323032 116612
rect 323084 116600 323090 116612
rect 340966 116600 340972 116612
rect 323084 116572 340972 116600
rect 323084 116560 323090 116572
rect 340966 116560 340972 116572
rect 341024 116560 341030 116612
rect 256050 116084 256056 116136
rect 256108 116124 256114 116136
rect 266078 116124 266084 116136
rect 256108 116096 266084 116124
rect 256108 116084 256114 116096
rect 266078 116084 266084 116096
rect 266136 116084 266142 116136
rect 176194 116016 176200 116068
rect 176252 116056 176258 116068
rect 213914 116056 213920 116068
rect 176252 116028 213920 116056
rect 176252 116016 176258 116028
rect 213914 116016 213920 116028
rect 213972 116016 213978 116068
rect 242250 116016 242256 116068
rect 242308 116056 242314 116068
rect 265986 116056 265992 116068
rect 242308 116028 265992 116056
rect 242308 116016 242314 116028
rect 265986 116016 265992 116028
rect 266044 116016 266050 116068
rect 173342 115948 173348 116000
rect 173400 115988 173406 116000
rect 214006 115988 214012 116000
rect 173400 115960 214012 115988
rect 173400 115948 173406 115960
rect 214006 115948 214012 115960
rect 214064 115948 214070 116000
rect 240962 115948 240968 116000
rect 241020 115988 241026 116000
rect 265710 115988 265716 116000
rect 241020 115960 265716 115988
rect 241020 115948 241026 115960
rect 265710 115948 265716 115960
rect 265768 115948 265774 116000
rect 282546 115880 282552 115932
rect 282604 115920 282610 115932
rect 306466 115920 306472 115932
rect 282604 115892 306472 115920
rect 282604 115880 282610 115892
rect 306466 115880 306472 115892
rect 306524 115880 306530 115932
rect 330478 115880 330484 115932
rect 330536 115920 330542 115932
rect 347498 115920 347504 115932
rect 330536 115892 347504 115920
rect 330536 115880 330542 115892
rect 347498 115880 347504 115892
rect 347556 115880 347562 115932
rect 430574 115880 430580 115932
rect 430632 115920 430638 115932
rect 434806 115920 434812 115932
rect 430632 115892 434812 115920
rect 430632 115880 430638 115892
rect 434806 115880 434812 115892
rect 434864 115880 434870 115932
rect 282822 115812 282828 115864
rect 282880 115852 282886 115864
rect 302326 115852 302332 115864
rect 282880 115824 302332 115852
rect 282880 115812 282886 115824
rect 302326 115812 302332 115824
rect 302384 115812 302390 115864
rect 230658 115744 230664 115796
rect 230716 115784 230722 115796
rect 240870 115784 240876 115796
rect 230716 115756 240876 115784
rect 230716 115744 230722 115756
rect 240870 115744 240876 115756
rect 240928 115744 240934 115796
rect 231670 115472 231676 115524
rect 231728 115512 231734 115524
rect 238202 115512 238208 115524
rect 231728 115484 238208 115512
rect 231728 115472 231734 115484
rect 238202 115472 238208 115484
rect 238260 115472 238266 115524
rect 230566 114792 230572 114844
rect 230624 114832 230630 114844
rect 232590 114832 232596 114844
rect 230624 114804 232596 114832
rect 230624 114792 230630 114804
rect 232590 114792 232596 114804
rect 232648 114792 232654 114844
rect 247862 114656 247868 114708
rect 247920 114696 247926 114708
rect 265986 114696 265992 114708
rect 247920 114668 265992 114696
rect 247920 114656 247926 114668
rect 265986 114656 265992 114668
rect 266044 114656 266050 114708
rect 209222 114588 209228 114640
rect 209280 114628 209286 114640
rect 213914 114628 213920 114640
rect 209280 114600 213920 114628
rect 209280 114588 209286 114600
rect 213914 114588 213920 114600
rect 213972 114588 213978 114640
rect 240778 114588 240784 114640
rect 240836 114628 240842 114640
rect 265710 114628 265716 114640
rect 240836 114600 265716 114628
rect 240836 114588 240842 114600
rect 265710 114588 265716 114600
rect 265768 114588 265774 114640
rect 169202 114520 169208 114572
rect 169260 114560 169266 114572
rect 214006 114560 214012 114572
rect 169260 114532 214012 114560
rect 169260 114520 169266 114532
rect 214006 114520 214012 114532
rect 214064 114520 214070 114572
rect 238294 114520 238300 114572
rect 238352 114560 238358 114572
rect 265250 114560 265256 114572
rect 238352 114532 265256 114560
rect 238352 114520 238358 114532
rect 265250 114520 265256 114532
rect 265308 114520 265314 114572
rect 231762 114452 231768 114504
rect 231820 114492 231826 114504
rect 252186 114492 252192 114504
rect 231820 114464 252192 114492
rect 231820 114452 231826 114464
rect 252186 114452 252192 114464
rect 252244 114452 252250 114504
rect 430850 114452 430856 114504
rect 430908 114492 430914 114504
rect 447134 114492 447140 114504
rect 430908 114464 447140 114492
rect 430908 114452 430914 114464
rect 447134 114452 447140 114464
rect 447192 114452 447198 114504
rect 230566 114384 230572 114436
rect 230624 114424 230630 114436
rect 234154 114424 234160 114436
rect 230624 114396 234160 114424
rect 230624 114384 230630 114396
rect 234154 114384 234160 114396
rect 234212 114384 234218 114436
rect 430574 114384 430580 114436
rect 430632 114424 430638 114436
rect 445846 114424 445852 114436
rect 430632 114396 445852 114424
rect 430632 114384 430638 114396
rect 445846 114384 445852 114396
rect 445904 114384 445910 114436
rect 230658 113772 230664 113824
rect 230716 113812 230722 113824
rect 249150 113812 249156 113824
rect 230716 113784 249156 113812
rect 230716 113772 230722 113784
rect 249150 113772 249156 113784
rect 249208 113772 249214 113824
rect 252094 113296 252100 113348
rect 252152 113336 252158 113348
rect 265710 113336 265716 113348
rect 252152 113308 265716 113336
rect 252152 113296 252158 113308
rect 265710 113296 265716 113308
rect 265768 113296 265774 113348
rect 198182 113228 198188 113280
rect 198240 113268 198246 113280
rect 213914 113268 213920 113280
rect 198240 113240 213920 113268
rect 198240 113228 198246 113240
rect 213914 113228 213920 113240
rect 213972 113228 213978 113280
rect 251910 113228 251916 113280
rect 251968 113268 251974 113280
rect 265250 113268 265256 113280
rect 251968 113240 265256 113268
rect 251968 113228 251974 113240
rect 265250 113228 265256 113240
rect 265308 113228 265314 113280
rect 167730 113160 167736 113212
rect 167788 113200 167794 113212
rect 214006 113200 214012 113212
rect 167788 113172 214012 113200
rect 167788 113160 167794 113172
rect 214006 113160 214012 113172
rect 214064 113160 214070 113212
rect 229738 113160 229744 113212
rect 229796 113200 229802 113212
rect 265710 113200 265716 113212
rect 229796 113172 265716 113200
rect 229796 113160 229802 113172
rect 265710 113160 265716 113172
rect 265768 113160 265774 113212
rect 282086 113092 282092 113144
rect 282144 113132 282150 113144
rect 295334 113132 295340 113144
rect 282144 113104 295340 113132
rect 282144 113092 282150 113104
rect 295334 113092 295340 113104
rect 295392 113092 295398 113144
rect 231762 112820 231768 112872
rect 231820 112860 231826 112872
rect 236730 112860 236736 112872
rect 231820 112832 236736 112860
rect 231820 112820 231826 112832
rect 236730 112820 236736 112832
rect 236788 112820 236794 112872
rect 230566 112480 230572 112532
rect 230624 112520 230630 112532
rect 249242 112520 249248 112532
rect 230624 112492 249248 112520
rect 230624 112480 230630 112492
rect 249242 112480 249248 112492
rect 249300 112480 249306 112532
rect 231118 112412 231124 112464
rect 231176 112452 231182 112464
rect 264330 112452 264336 112464
rect 231176 112424 264336 112452
rect 231176 112412 231182 112424
rect 264330 112412 264336 112424
rect 264388 112412 264394 112464
rect 188522 111868 188528 111920
rect 188580 111908 188586 111920
rect 213914 111908 213920 111920
rect 188580 111880 213920 111908
rect 188580 111868 188586 111880
rect 213914 111868 213920 111880
rect 213972 111868 213978 111920
rect 181530 111800 181536 111852
rect 181588 111840 181594 111852
rect 214006 111840 214012 111852
rect 181588 111812 214012 111840
rect 181588 111800 181594 111812
rect 214006 111800 214012 111812
rect 214064 111800 214070 111852
rect 249150 111800 249156 111852
rect 249208 111840 249214 111852
rect 265710 111840 265716 111852
rect 249208 111812 265716 111840
rect 249208 111800 249214 111812
rect 265710 111800 265716 111812
rect 265768 111800 265774 111852
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 14458 111772 14464 111784
rect 3476 111744 14464 111772
rect 3476 111732 3482 111744
rect 14458 111732 14464 111744
rect 14516 111732 14522 111784
rect 167914 111732 167920 111784
rect 167972 111772 167978 111784
rect 177482 111772 177488 111784
rect 167972 111744 177488 111772
rect 167972 111732 167978 111744
rect 177482 111732 177488 111744
rect 177540 111732 177546 111784
rect 231762 111732 231768 111784
rect 231820 111772 231826 111784
rect 264514 111772 264520 111784
rect 231820 111744 264520 111772
rect 231820 111732 231826 111744
rect 264514 111732 264520 111744
rect 264572 111732 264578 111784
rect 282822 111732 282828 111784
rect 282880 111772 282886 111784
rect 296714 111772 296720 111784
rect 282880 111744 296720 111772
rect 282880 111732 282886 111744
rect 296714 111732 296720 111744
rect 296772 111732 296778 111784
rect 430574 111732 430580 111784
rect 430632 111772 430638 111784
rect 451274 111772 451280 111784
rect 430632 111744 451280 111772
rect 430632 111732 430638 111744
rect 451274 111732 451280 111744
rect 451332 111732 451338 111784
rect 231486 111664 231492 111716
rect 231544 111704 231550 111716
rect 235258 111704 235264 111716
rect 231544 111676 235264 111704
rect 231544 111664 231550 111676
rect 235258 111664 235264 111676
rect 235316 111664 235322 111716
rect 316034 111052 316040 111104
rect 316092 111092 316098 111104
rect 327718 111092 327724 111104
rect 316092 111064 327724 111092
rect 316092 111052 316098 111064
rect 327718 111052 327724 111064
rect 327776 111052 327782 111104
rect 329834 111052 329840 111104
rect 329892 111092 329898 111104
rect 345198 111092 345204 111104
rect 329892 111064 345204 111092
rect 329892 111052 329898 111064
rect 345198 111052 345204 111064
rect 345256 111052 345262 111104
rect 238202 110576 238208 110628
rect 238260 110616 238266 110628
rect 265986 110616 265992 110628
rect 238260 110588 265992 110616
rect 238260 110576 238266 110588
rect 265986 110576 265992 110588
rect 266044 110576 266050 110628
rect 207750 110508 207756 110560
rect 207808 110548 207814 110560
rect 214006 110548 214012 110560
rect 207808 110520 214012 110548
rect 207808 110508 207814 110520
rect 214006 110508 214012 110520
rect 214064 110508 214070 110560
rect 166258 110440 166264 110492
rect 166316 110480 166322 110492
rect 213914 110480 213920 110492
rect 166316 110452 213920 110480
rect 166316 110440 166322 110452
rect 213914 110440 213920 110452
rect 213972 110440 213978 110492
rect 260282 110440 260288 110492
rect 260340 110480 260346 110492
rect 265710 110480 265716 110492
rect 260340 110452 265716 110480
rect 260340 110440 260346 110452
rect 265710 110440 265716 110452
rect 265768 110440 265774 110492
rect 168098 110372 168104 110424
rect 168156 110412 168162 110424
rect 178862 110412 178868 110424
rect 168156 110384 178868 110412
rect 168156 110372 168162 110384
rect 178862 110372 178868 110384
rect 178920 110372 178926 110424
rect 231762 110372 231768 110424
rect 231820 110412 231826 110424
rect 257522 110412 257528 110424
rect 231820 110384 257528 110412
rect 231820 110372 231826 110384
rect 257522 110372 257528 110384
rect 257580 110372 257586 110424
rect 282270 110372 282276 110424
rect 282328 110412 282334 110424
rect 294046 110412 294052 110424
rect 282328 110384 294052 110412
rect 282328 110372 282334 110384
rect 294046 110372 294052 110384
rect 294104 110372 294110 110424
rect 344278 110372 344284 110424
rect 344336 110412 344342 110424
rect 347038 110412 347044 110424
rect 344336 110384 347044 110412
rect 344336 110372 344342 110384
rect 347038 110372 347044 110384
rect 347096 110372 347102 110424
rect 231762 109964 231768 110016
rect 231820 110004 231826 110016
rect 235442 110004 235448 110016
rect 231820 109976 235448 110004
rect 231820 109964 231826 109976
rect 235442 109964 235448 109976
rect 235500 109964 235506 110016
rect 257614 109148 257620 109200
rect 257672 109188 257678 109200
rect 265710 109188 265716 109200
rect 257672 109160 265716 109188
rect 257672 109148 257678 109160
rect 265710 109148 265716 109160
rect 265768 109148 265774 109200
rect 206462 109080 206468 109132
rect 206520 109120 206526 109132
rect 214006 109120 214012 109132
rect 206520 109092 214012 109120
rect 206520 109080 206526 109092
rect 214006 109080 214012 109092
rect 214064 109080 214070 109132
rect 235258 109080 235264 109132
rect 235316 109120 235322 109132
rect 265158 109120 265164 109132
rect 235316 109092 265164 109120
rect 235316 109080 235322 109092
rect 265158 109080 265164 109092
rect 265216 109080 265222 109132
rect 171962 109012 171968 109064
rect 172020 109052 172026 109064
rect 213914 109052 213920 109064
rect 172020 109024 213920 109052
rect 172020 109012 172026 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 234062 109012 234068 109064
rect 234120 109052 234126 109064
rect 265526 109052 265532 109064
rect 234120 109024 265532 109052
rect 234120 109012 234126 109024
rect 265526 109012 265532 109024
rect 265584 109012 265590 109064
rect 167914 108944 167920 108996
rect 167972 108984 167978 108996
rect 180242 108984 180248 108996
rect 167972 108956 180248 108984
rect 167972 108944 167978 108956
rect 180242 108944 180248 108956
rect 180300 108944 180306 108996
rect 231762 108944 231768 108996
rect 231820 108984 231826 108996
rect 260374 108984 260380 108996
rect 231820 108956 260380 108984
rect 231820 108944 231826 108956
rect 260374 108944 260380 108956
rect 260432 108944 260438 108996
rect 301498 108944 301504 108996
rect 301556 108984 301562 108996
rect 347498 108984 347504 108996
rect 301556 108956 347504 108984
rect 301556 108944 301562 108956
rect 347498 108944 347504 108956
rect 347556 108944 347562 108996
rect 430574 108944 430580 108996
rect 430632 108984 430638 108996
rect 434714 108984 434720 108996
rect 430632 108956 434720 108984
rect 430632 108944 430638 108956
rect 434714 108944 434720 108956
rect 434772 108944 434778 108996
rect 231670 108876 231676 108928
rect 231728 108916 231734 108928
rect 239582 108916 239588 108928
rect 231728 108888 239588 108916
rect 231728 108876 231734 108888
rect 239582 108876 239588 108888
rect 239640 108876 239646 108928
rect 231394 108264 231400 108316
rect 231452 108304 231458 108316
rect 253474 108304 253480 108316
rect 231452 108276 253480 108304
rect 231452 108264 231458 108276
rect 253474 108264 253480 108276
rect 253532 108264 253538 108316
rect 240870 107856 240876 107908
rect 240928 107896 240934 107908
rect 265710 107896 265716 107908
rect 240928 107868 265716 107896
rect 240928 107856 240934 107868
rect 265710 107856 265716 107868
rect 265768 107856 265774 107908
rect 281534 107856 281540 107908
rect 281592 107896 281598 107908
rect 283190 107896 283196 107908
rect 281592 107868 283196 107896
rect 281592 107856 281598 107868
rect 283190 107856 283196 107868
rect 283248 107856 283254 107908
rect 261570 107788 261576 107840
rect 261628 107828 261634 107840
rect 265986 107828 265992 107840
rect 261628 107800 265992 107828
rect 261628 107788 261634 107800
rect 265986 107788 265992 107800
rect 266044 107788 266050 107840
rect 178862 107720 178868 107772
rect 178920 107760 178926 107772
rect 214006 107760 214012 107772
rect 178920 107732 214012 107760
rect 178920 107720 178926 107732
rect 214006 107720 214012 107732
rect 214064 107720 214070 107772
rect 253290 107720 253296 107772
rect 253348 107760 253354 107772
rect 265710 107760 265716 107772
rect 253348 107732 265716 107760
rect 253348 107720 253354 107732
rect 265710 107720 265716 107732
rect 265768 107720 265774 107772
rect 174722 107652 174728 107704
rect 174780 107692 174786 107704
rect 213914 107692 213920 107704
rect 174780 107664 213920 107692
rect 174780 107652 174786 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 263042 107652 263048 107704
rect 263100 107692 263106 107704
rect 265158 107692 265164 107704
rect 263100 107664 265164 107692
rect 263100 107652 263106 107664
rect 265158 107652 265164 107664
rect 265216 107652 265222 107704
rect 231762 107584 231768 107636
rect 231820 107624 231826 107636
rect 256234 107624 256240 107636
rect 231820 107596 256240 107624
rect 231820 107584 231826 107596
rect 256234 107584 256240 107596
rect 256292 107584 256298 107636
rect 333330 107584 333336 107636
rect 333388 107624 333394 107636
rect 347498 107624 347504 107636
rect 333388 107596 347504 107624
rect 333388 107584 333394 107596
rect 347498 107584 347504 107596
rect 347556 107584 347562 107636
rect 430574 107584 430580 107636
rect 430632 107624 430638 107636
rect 442994 107624 443000 107636
rect 430632 107596 443000 107624
rect 430632 107584 430638 107596
rect 442994 107584 443000 107596
rect 443052 107584 443058 107636
rect 231670 107516 231676 107568
rect 231728 107556 231734 107568
rect 246482 107556 246488 107568
rect 231728 107528 246488 107556
rect 231728 107516 231734 107528
rect 246482 107516 246488 107528
rect 246540 107516 246546 107568
rect 231762 107040 231768 107092
rect 231820 107080 231826 107092
rect 236914 107080 236920 107092
rect 231820 107052 236920 107080
rect 231820 107040 231826 107052
rect 236914 107040 236920 107052
rect 236972 107040 236978 107092
rect 177482 106360 177488 106412
rect 177540 106400 177546 106412
rect 214006 106400 214012 106412
rect 177540 106372 214012 106400
rect 177540 106360 177546 106372
rect 214006 106360 214012 106372
rect 214064 106360 214070 106412
rect 249242 106360 249248 106412
rect 249300 106400 249306 106412
rect 265526 106400 265532 106412
rect 249300 106372 265532 106400
rect 249300 106360 249306 106372
rect 265526 106360 265532 106372
rect 265584 106360 265590 106412
rect 170398 106292 170404 106344
rect 170456 106332 170462 106344
rect 213914 106332 213920 106344
rect 170456 106304 213920 106332
rect 170456 106292 170462 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 245194 106292 245200 106344
rect 245252 106332 245258 106344
rect 265710 106332 265716 106344
rect 245252 106304 265716 106332
rect 245252 106292 245258 106304
rect 265710 106292 265716 106304
rect 265768 106292 265774 106344
rect 231762 106224 231768 106276
rect 231820 106264 231826 106276
rect 261846 106264 261852 106276
rect 231820 106236 261852 106264
rect 231820 106224 231826 106236
rect 261846 106224 261852 106236
rect 261904 106224 261910 106276
rect 262858 106224 262864 106276
rect 262916 106264 262922 106276
rect 267182 106264 267188 106276
rect 262916 106236 267188 106264
rect 262916 106224 262922 106236
rect 267182 106224 267188 106236
rect 267240 106224 267246 106276
rect 430574 106224 430580 106276
rect 430632 106264 430638 106276
rect 438854 106264 438860 106276
rect 430632 106236 438860 106264
rect 430632 106224 430638 106236
rect 438854 106224 438860 106236
rect 438912 106224 438918 106276
rect 231670 105340 231676 105392
rect 231728 105380 231734 105392
rect 235534 105380 235540 105392
rect 231728 105352 235540 105380
rect 231728 105340 231734 105352
rect 235534 105340 235540 105352
rect 235592 105340 235598 105392
rect 192570 105000 192576 105052
rect 192628 105040 192634 105052
rect 214006 105040 214012 105052
rect 192628 105012 214012 105040
rect 192628 105000 192634 105012
rect 214006 105000 214012 105012
rect 214064 105000 214070 105052
rect 261754 105000 261760 105052
rect 261812 105040 261818 105052
rect 265526 105040 265532 105052
rect 261812 105012 265532 105040
rect 261812 105000 261818 105012
rect 265526 105000 265532 105012
rect 265584 105000 265590 105052
rect 205082 104932 205088 104984
rect 205140 104972 205146 104984
rect 213914 104972 213920 104984
rect 205140 104944 213920 104972
rect 205140 104932 205146 104944
rect 213914 104932 213920 104944
rect 213972 104932 213978 104984
rect 256234 104932 256240 104984
rect 256292 104972 256298 104984
rect 265986 104972 265992 104984
rect 256292 104944 265992 104972
rect 256292 104932 256298 104944
rect 265986 104932 265992 104944
rect 266044 104932 266050 104984
rect 239582 104864 239588 104916
rect 239640 104904 239646 104916
rect 265710 104904 265716 104916
rect 239640 104876 265716 104904
rect 239640 104864 239646 104876
rect 265710 104864 265716 104876
rect 265768 104864 265774 104916
rect 231762 104796 231768 104848
rect 231820 104836 231826 104848
rect 264606 104836 264612 104848
rect 231820 104808 264612 104836
rect 231820 104796 231826 104808
rect 264606 104796 264612 104808
rect 264664 104796 264670 104848
rect 281994 104796 282000 104848
rect 282052 104836 282058 104848
rect 284478 104836 284484 104848
rect 282052 104808 284484 104836
rect 282052 104796 282058 104808
rect 284478 104796 284484 104808
rect 284536 104796 284542 104848
rect 311158 104796 311164 104848
rect 311216 104836 311222 104848
rect 347038 104836 347044 104848
rect 311216 104808 347044 104836
rect 311216 104796 311222 104808
rect 347038 104796 347044 104808
rect 347096 104796 347102 104848
rect 430574 104796 430580 104848
rect 430632 104836 430638 104848
rect 441614 104836 441620 104848
rect 430632 104808 441620 104836
rect 430632 104796 430638 104808
rect 441614 104796 441620 104808
rect 441672 104796 441678 104848
rect 231486 104728 231492 104780
rect 231544 104768 231550 104780
rect 242342 104768 242348 104780
rect 231544 104740 242348 104768
rect 231544 104728 231550 104740
rect 242342 104728 242348 104740
rect 242400 104728 242406 104780
rect 231670 104660 231676 104712
rect 231728 104700 231734 104712
rect 234246 104700 234252 104712
rect 231728 104672 234252 104700
rect 231728 104660 231734 104672
rect 234246 104660 234252 104672
rect 234304 104660 234310 104712
rect 262858 103708 262864 103760
rect 262916 103748 262922 103760
rect 265986 103748 265992 103760
rect 262916 103720 265992 103748
rect 262916 103708 262922 103720
rect 265986 103708 265992 103720
rect 266044 103708 266050 103760
rect 242434 103640 242440 103692
rect 242492 103680 242498 103692
rect 265710 103680 265716 103692
rect 242492 103652 265716 103680
rect 242492 103640 242498 103652
rect 265710 103640 265716 103652
rect 265768 103640 265774 103692
rect 202322 103572 202328 103624
rect 202380 103612 202386 103624
rect 214006 103612 214012 103624
rect 202380 103584 214012 103612
rect 202380 103572 202386 103584
rect 214006 103572 214012 103584
rect 214064 103572 214070 103624
rect 199378 103504 199384 103556
rect 199436 103544 199442 103556
rect 213914 103544 213920 103556
rect 199436 103516 213920 103544
rect 199436 103504 199442 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 430574 103436 430580 103488
rect 430632 103476 430638 103488
rect 440326 103476 440332 103488
rect 430632 103448 440332 103476
rect 430632 103436 430638 103448
rect 440326 103436 440332 103448
rect 440384 103436 440390 103488
rect 430758 103368 430764 103420
rect 430816 103408 430822 103420
rect 437474 103408 437480 103420
rect 430816 103380 437480 103408
rect 430816 103368 430822 103380
rect 437474 103368 437480 103380
rect 437532 103368 437538 103420
rect 230566 102960 230572 103012
rect 230624 103000 230630 103012
rect 232498 103000 232504 103012
rect 230624 102972 232504 103000
rect 230624 102960 230630 102972
rect 232498 102960 232504 102972
rect 232556 102960 232562 103012
rect 175918 102756 175924 102808
rect 175976 102796 175982 102808
rect 216214 102796 216220 102808
rect 175976 102768 216220 102796
rect 175976 102756 175982 102768
rect 216214 102756 216220 102768
rect 216272 102756 216278 102808
rect 293954 102756 293960 102808
rect 294012 102796 294018 102808
rect 342254 102796 342260 102808
rect 294012 102768 342260 102796
rect 294012 102756 294018 102768
rect 342254 102756 342260 102768
rect 342312 102756 342318 102808
rect 253474 102348 253480 102400
rect 253532 102388 253538 102400
rect 264606 102388 264612 102400
rect 253532 102360 264612 102388
rect 253532 102348 253538 102360
rect 264606 102348 264612 102360
rect 264664 102348 264670 102400
rect 233602 102280 233608 102332
rect 233660 102320 233666 102332
rect 266078 102320 266084 102332
rect 233660 102292 266084 102320
rect 233660 102280 233666 102292
rect 266078 102280 266084 102292
rect 266136 102280 266142 102332
rect 232590 102212 232596 102264
rect 232648 102252 232654 102264
rect 265710 102252 265716 102264
rect 232648 102224 265716 102252
rect 232648 102212 232654 102224
rect 265710 102212 265716 102224
rect 265768 102212 265774 102264
rect 200850 102144 200856 102196
rect 200908 102184 200914 102196
rect 213914 102184 213920 102196
rect 200908 102156 213920 102184
rect 200908 102144 200914 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 231118 102144 231124 102196
rect 231176 102184 231182 102196
rect 265158 102184 265164 102196
rect 231176 102156 265164 102184
rect 231176 102144 231182 102156
rect 265158 102144 265164 102156
rect 265216 102144 265222 102196
rect 231486 102076 231492 102128
rect 231544 102116 231550 102128
rect 233970 102116 233976 102128
rect 231544 102088 233976 102116
rect 231544 102076 231550 102088
rect 233970 102076 233976 102088
rect 234028 102076 234034 102128
rect 282822 102076 282828 102128
rect 282880 102116 282886 102128
rect 290090 102116 290096 102128
rect 282880 102088 290096 102116
rect 282880 102076 282886 102088
rect 290090 102076 290096 102088
rect 290148 102076 290154 102128
rect 336274 102076 336280 102128
rect 336332 102116 336338 102128
rect 347222 102116 347228 102128
rect 336332 102088 347228 102116
rect 336332 102076 336338 102088
rect 347222 102076 347228 102088
rect 347280 102076 347286 102128
rect 430574 102076 430580 102128
rect 430632 102116 430638 102128
rect 448514 102116 448520 102128
rect 430632 102088 448520 102116
rect 430632 102076 430638 102088
rect 448514 102076 448520 102088
rect 448572 102076 448578 102128
rect 231762 101940 231768 101992
rect 231820 101980 231826 101992
rect 259086 101980 259092 101992
rect 231820 101952 259092 101980
rect 231820 101940 231826 101952
rect 259086 101940 259092 101952
rect 259144 101940 259150 101992
rect 231578 101464 231584 101516
rect 231636 101504 231642 101516
rect 235350 101504 235356 101516
rect 231636 101476 235356 101504
rect 231636 101464 231642 101476
rect 235350 101464 235356 101476
rect 235408 101464 235414 101516
rect 231670 101396 231676 101448
rect 231728 101436 231734 101448
rect 254670 101436 254676 101448
rect 231728 101408 254676 101436
rect 231728 101396 231734 101408
rect 254670 101396 254676 101408
rect 254728 101396 254734 101448
rect 280430 101396 280436 101448
rect 280488 101436 280494 101448
rect 343634 101436 343640 101448
rect 280488 101408 343640 101436
rect 280488 101396 280494 101408
rect 343634 101396 343640 101408
rect 343692 101396 343698 101448
rect 258994 100852 259000 100904
rect 259052 100892 259058 100904
rect 265710 100892 265716 100904
rect 259052 100864 265716 100892
rect 259052 100852 259058 100864
rect 265710 100852 265716 100864
rect 265768 100852 265774 100904
rect 257522 100784 257528 100836
rect 257580 100824 257586 100836
rect 265342 100824 265348 100836
rect 257580 100796 265348 100824
rect 257580 100784 257586 100796
rect 265342 100784 265348 100796
rect 265400 100784 265406 100836
rect 203702 100716 203708 100768
rect 203760 100756 203766 100768
rect 213914 100756 213920 100768
rect 203760 100728 213920 100756
rect 203760 100716 203766 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 246482 100716 246488 100768
rect 246540 100756 246546 100768
rect 265526 100756 265532 100768
rect 246540 100728 265532 100756
rect 246540 100716 246546 100728
rect 265526 100716 265532 100728
rect 265584 100716 265590 100768
rect 231762 100648 231768 100700
rect 231820 100688 231826 100700
rect 241054 100688 241060 100700
rect 231820 100660 241060 100688
rect 231820 100648 231826 100660
rect 241054 100648 241060 100660
rect 241112 100648 241118 100700
rect 319438 100648 319444 100700
rect 319496 100688 319502 100700
rect 347498 100688 347504 100700
rect 319496 100660 347504 100688
rect 319496 100648 319502 100660
rect 347498 100648 347504 100660
rect 347556 100648 347562 100700
rect 436738 100648 436744 100700
rect 436796 100688 436802 100700
rect 580166 100688 580172 100700
rect 436796 100660 580172 100688
rect 436796 100648 436802 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 284294 99968 284300 100020
rect 284352 100008 284358 100020
rect 345014 100008 345020 100020
rect 284352 99980 345020 100008
rect 284352 99968 284358 99980
rect 345014 99968 345020 99980
rect 345072 99968 345078 100020
rect 230934 99560 230940 99612
rect 230992 99600 230998 99612
rect 232774 99600 232780 99612
rect 230992 99572 232780 99600
rect 230992 99560 230998 99572
rect 232774 99560 232780 99572
rect 232832 99560 232838 99612
rect 254670 99492 254676 99544
rect 254728 99532 254734 99544
rect 265526 99532 265532 99544
rect 254728 99504 265532 99532
rect 254728 99492 254734 99504
rect 265526 99492 265532 99504
rect 265584 99492 265590 99544
rect 169294 99424 169300 99476
rect 169352 99464 169358 99476
rect 213914 99464 213920 99476
rect 169352 99436 213920 99464
rect 169352 99424 169358 99436
rect 213914 99424 213920 99436
rect 213972 99424 213978 99476
rect 238110 99424 238116 99476
rect 238168 99464 238174 99476
rect 265710 99464 265716 99476
rect 238168 99436 265716 99464
rect 238168 99424 238174 99436
rect 265710 99424 265716 99436
rect 265768 99424 265774 99476
rect 164878 99356 164884 99408
rect 164936 99396 164942 99408
rect 214006 99396 214012 99408
rect 164936 99368 214012 99396
rect 164936 99356 164942 99368
rect 214006 99356 214012 99368
rect 214064 99356 214070 99408
rect 236730 99356 236736 99408
rect 236788 99396 236794 99408
rect 265986 99396 265992 99408
rect 236788 99368 265992 99396
rect 236788 99356 236794 99368
rect 265986 99356 265992 99368
rect 266044 99356 266050 99408
rect 230474 98200 230480 98252
rect 230532 98240 230538 98252
rect 232682 98240 232688 98252
rect 230532 98212 232688 98240
rect 230532 98200 230538 98212
rect 232682 98200 232688 98212
rect 232740 98200 232746 98252
rect 248966 98132 248972 98184
rect 249024 98172 249030 98184
rect 266078 98172 266084 98184
rect 249024 98144 266084 98172
rect 249024 98132 249030 98144
rect 266078 98132 266084 98144
rect 266136 98132 266142 98184
rect 167914 98064 167920 98116
rect 167972 98104 167978 98116
rect 214006 98104 214012 98116
rect 167972 98076 214012 98104
rect 167972 98064 167978 98076
rect 214006 98064 214012 98076
rect 214064 98064 214070 98116
rect 232498 98064 232504 98116
rect 232556 98104 232562 98116
rect 264606 98104 264612 98116
rect 232556 98076 264612 98104
rect 232556 98064 232562 98076
rect 264606 98064 264612 98076
rect 264664 98064 264670 98116
rect 166442 97996 166448 98048
rect 166500 98036 166506 98048
rect 213914 98036 213920 98048
rect 166500 98008 213920 98036
rect 166500 97996 166506 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 231210 97996 231216 98048
rect 231268 98036 231274 98048
rect 265618 98036 265624 98048
rect 231268 98008 265624 98036
rect 231268 97996 231274 98008
rect 265618 97996 265624 98008
rect 265676 97996 265682 98048
rect 316678 97928 316684 97980
rect 316736 97968 316742 97980
rect 347498 97968 347504 97980
rect 316736 97940 347504 97968
rect 316736 97928 316742 97940
rect 347498 97928 347504 97940
rect 347556 97928 347562 97980
rect 430574 97928 430580 97980
rect 430632 97968 430638 97980
rect 443086 97968 443092 97980
rect 430632 97940 443092 97968
rect 430632 97928 430638 97940
rect 443086 97928 443092 97940
rect 443144 97928 443150 97980
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 166534 97248 166540 97300
rect 166592 97288 166598 97300
rect 214650 97288 214656 97300
rect 166592 97260 214656 97288
rect 166592 97248 166598 97260
rect 214650 97248 214656 97260
rect 214708 97248 214714 97300
rect 231762 96704 231768 96756
rect 231820 96744 231826 96756
rect 239674 96744 239680 96756
rect 231820 96716 239680 96744
rect 231820 96704 231826 96716
rect 239674 96704 239680 96716
rect 239732 96704 239738 96756
rect 260374 96704 260380 96756
rect 260432 96744 260438 96756
rect 264606 96744 264612 96756
rect 260432 96716 264612 96744
rect 260432 96704 260438 96716
rect 264606 96704 264612 96716
rect 264664 96704 264670 96756
rect 210602 96636 210608 96688
rect 210660 96676 210666 96688
rect 213914 96676 213920 96688
rect 210660 96648 213920 96676
rect 210660 96636 210666 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 230474 96636 230480 96688
rect 230532 96676 230538 96688
rect 233970 96676 233976 96688
rect 230532 96648 233976 96676
rect 230532 96636 230538 96648
rect 233970 96636 233976 96648
rect 234028 96636 234034 96688
rect 235350 96636 235356 96688
rect 235408 96676 235414 96688
rect 261386 96676 261392 96688
rect 235408 96648 261392 96676
rect 235408 96636 235414 96648
rect 261386 96636 261392 96648
rect 261444 96636 261450 96688
rect 348878 96568 348884 96620
rect 348936 96608 348942 96620
rect 580350 96608 580356 96620
rect 348936 96580 580356 96608
rect 348936 96568 348942 96580
rect 580350 96568 580356 96580
rect 580408 96568 580414 96620
rect 329098 96500 329104 96552
rect 329156 96540 329162 96552
rect 428090 96540 428096 96552
rect 329156 96512 428096 96540
rect 329156 96500 329162 96512
rect 428090 96500 428096 96512
rect 428148 96500 428154 96552
rect 188430 96364 188436 96416
rect 188488 96404 188494 96416
rect 281534 96404 281540 96416
rect 188488 96376 281540 96404
rect 188488 96364 188494 96376
rect 281534 96364 281540 96376
rect 281592 96364 281598 96416
rect 226978 95888 226984 95940
rect 227036 95928 227042 95940
rect 248966 95928 248972 95940
rect 227036 95900 248972 95928
rect 227036 95888 227042 95900
rect 248966 95888 248972 95900
rect 249024 95888 249030 95940
rect 204990 95208 204996 95260
rect 205048 95248 205054 95260
rect 213914 95248 213920 95260
rect 205048 95220 213920 95248
rect 205048 95208 205054 95220
rect 213914 95208 213920 95220
rect 213972 95208 213978 95260
rect 228358 95208 228364 95260
rect 228416 95248 228422 95260
rect 265526 95248 265532 95260
rect 228416 95220 265532 95248
rect 228416 95208 228422 95220
rect 265526 95208 265532 95220
rect 265584 95208 265590 95260
rect 318058 95208 318064 95260
rect 318116 95248 318122 95260
rect 389450 95248 389456 95260
rect 318116 95220 389456 95248
rect 318116 95208 318122 95220
rect 389450 95208 389456 95220
rect 389508 95208 389514 95260
rect 209038 95140 209044 95192
rect 209096 95180 209102 95192
rect 427630 95180 427636 95192
rect 209096 95152 427636 95180
rect 209096 95140 209102 95152
rect 427630 95140 427636 95152
rect 427688 95140 427694 95192
rect 196710 95072 196716 95124
rect 196768 95112 196774 95124
rect 280154 95112 280160 95124
rect 196768 95084 280160 95112
rect 196768 95072 196774 95084
rect 280154 95072 280160 95084
rect 280212 95072 280218 95124
rect 326338 95072 326344 95124
rect 326396 95112 326402 95124
rect 428182 95112 428188 95124
rect 326396 95084 428188 95112
rect 326396 95072 326402 95084
rect 428182 95072 428188 95084
rect 428240 95072 428246 95124
rect 203610 95004 203616 95056
rect 203668 95044 203674 95056
rect 280246 95044 280252 95056
rect 203668 95016 280252 95044
rect 203668 95004 203674 95016
rect 280246 95004 280252 95016
rect 280304 95004 280310 95056
rect 342898 95004 342904 95056
rect 342956 95044 342962 95056
rect 400214 95044 400220 95056
rect 342956 95016 400220 95044
rect 342956 95004 342962 95016
rect 400214 95004 400220 95016
rect 400272 95044 400278 95056
rect 400858 95044 400864 95056
rect 400272 95016 400864 95044
rect 400272 95004 400278 95016
rect 400858 95004 400864 95016
rect 400916 95004 400922 95056
rect 340138 94936 340144 94988
rect 340196 94976 340202 94988
rect 396166 94976 396172 94988
rect 340196 94948 396172 94976
rect 340196 94936 340202 94948
rect 396166 94936 396172 94948
rect 396224 94976 396230 94988
rect 397086 94976 397092 94988
rect 396224 94948 397092 94976
rect 396224 94936 396230 94948
rect 397086 94936 397092 94948
rect 397144 94936 397150 94988
rect 222838 94528 222844 94580
rect 222896 94568 222902 94580
rect 233602 94568 233608 94580
rect 222896 94540 233608 94568
rect 222896 94528 222902 94540
rect 233602 94528 233608 94540
rect 233660 94528 233666 94580
rect 130378 94460 130384 94512
rect 130436 94500 130442 94512
rect 214558 94500 214564 94512
rect 130436 94472 214564 94500
rect 130436 94460 130442 94472
rect 214558 94460 214564 94472
rect 214616 94460 214622 94512
rect 224218 94460 224224 94512
rect 224276 94500 224282 94512
rect 267274 94500 267280 94512
rect 224276 94472 267280 94500
rect 224276 94460 224282 94472
rect 267274 94460 267280 94472
rect 267332 94460 267338 94512
rect 120626 94052 120632 94104
rect 120684 94092 120690 94104
rect 167822 94092 167828 94104
rect 120684 94064 167828 94092
rect 120684 94052 120690 94064
rect 167822 94052 167828 94064
rect 167880 94052 167886 94104
rect 118234 93984 118240 94036
rect 118292 94024 118298 94036
rect 172054 94024 172060 94036
rect 118292 93996 172060 94024
rect 118292 93984 118298 93996
rect 172054 93984 172060 93996
rect 172112 93984 172118 94036
rect 106642 93916 106648 93968
rect 106700 93956 106706 93968
rect 170582 93956 170588 93968
rect 106700 93928 170588 93956
rect 106700 93916 106706 93928
rect 170582 93916 170588 93928
rect 170640 93916 170646 93968
rect 93854 93848 93860 93900
rect 93912 93888 93918 93900
rect 174722 93888 174728 93900
rect 93912 93860 174728 93888
rect 93912 93848 93918 93860
rect 174722 93848 174728 93860
rect 174780 93848 174786 93900
rect 67634 93780 67640 93832
rect 67692 93820 67698 93832
rect 199378 93820 199384 93832
rect 67692 93792 199384 93820
rect 67692 93780 67698 93792
rect 199378 93780 199384 93792
rect 199436 93780 199442 93832
rect 239674 93780 239680 93832
rect 239732 93820 239738 93832
rect 270954 93820 270960 93832
rect 239732 93792 270960 93820
rect 239732 93780 239738 93792
rect 270954 93780 270960 93792
rect 271012 93780 271018 93832
rect 347682 93780 347688 93832
rect 347740 93820 347746 93832
rect 582374 93820 582380 93832
rect 347740 93792 582380 93820
rect 347740 93780 347746 93792
rect 582374 93780 582380 93792
rect 582432 93780 582438 93832
rect 195330 93712 195336 93764
rect 195388 93752 195394 93764
rect 281902 93752 281908 93764
rect 195388 93724 281908 93752
rect 195388 93712 195394 93724
rect 281902 93712 281908 93724
rect 281960 93712 281966 93764
rect 349798 93712 349804 93764
rect 349856 93752 349862 93764
rect 360194 93752 360200 93764
rect 349856 93724 360200 93752
rect 349856 93712 349862 93724
rect 360194 93712 360200 93724
rect 360252 93712 360258 93764
rect 233970 93644 233976 93696
rect 234028 93684 234034 93696
rect 276934 93684 276940 93696
rect 234028 93656 276940 93684
rect 234028 93644 234034 93656
rect 276934 93644 276940 93656
rect 276992 93644 276998 93696
rect 345658 93644 345664 93696
rect 345716 93684 345722 93696
rect 356514 93684 356520 93696
rect 345716 93656 356520 93684
rect 345716 93644 345722 93656
rect 356514 93644 356520 93656
rect 356572 93644 356578 93696
rect 349890 93576 349896 93628
rect 349948 93616 349954 93628
rect 358814 93616 358820 93628
rect 349948 93588 358820 93616
rect 349948 93576 349954 93588
rect 358814 93576 358820 93588
rect 358872 93576 358878 93628
rect 270954 93440 270960 93492
rect 271012 93480 271018 93492
rect 351454 93480 351460 93492
rect 271012 93452 351460 93480
rect 271012 93440 271018 93452
rect 351454 93440 351460 93452
rect 351512 93440 351518 93492
rect 151722 93372 151728 93424
rect 151780 93412 151786 93424
rect 187050 93412 187056 93424
rect 151780 93384 187056 93412
rect 151780 93372 151786 93384
rect 187050 93372 187056 93384
rect 187108 93372 187114 93424
rect 114370 93304 114376 93356
rect 114428 93344 114434 93356
rect 173250 93344 173256 93356
rect 114428 93316 173256 93344
rect 114428 93304 114434 93316
rect 173250 93304 173256 93316
rect 173308 93304 173314 93356
rect 129458 93236 129464 93288
rect 129516 93276 129522 93288
rect 176010 93276 176016 93288
rect 129516 93248 176016 93276
rect 129516 93236 129522 93248
rect 176010 93236 176016 93248
rect 176068 93236 176074 93288
rect 113818 93168 113824 93220
rect 113876 93208 113882 93220
rect 185578 93208 185584 93220
rect 113876 93180 185584 93208
rect 113876 93168 113882 93180
rect 185578 93168 185584 93180
rect 185636 93168 185642 93220
rect 118694 93100 118700 93152
rect 118752 93140 118758 93152
rect 214742 93140 214748 93152
rect 118752 93112 214748 93140
rect 118752 93100 118758 93112
rect 214742 93100 214748 93112
rect 214800 93100 214806 93152
rect 399478 93100 399484 93152
rect 399536 93140 399542 93152
rect 406010 93140 406016 93152
rect 399536 93112 406016 93140
rect 399536 93100 399542 93112
rect 406010 93100 406016 93112
rect 406068 93100 406074 93152
rect 410518 93100 410524 93152
rect 410576 93140 410582 93152
rect 427446 93140 427452 93152
rect 410576 93112 427452 93140
rect 410576 93100 410582 93112
rect 427446 93100 427452 93112
rect 427504 93100 427510 93152
rect 348418 92692 348424 92744
rect 348476 92732 348482 92744
rect 353294 92732 353300 92744
rect 348476 92704 353300 92732
rect 348476 92692 348482 92704
rect 353294 92692 353300 92704
rect 353352 92732 353358 92744
rect 354030 92732 354036 92744
rect 353352 92704 354036 92732
rect 353352 92692 353358 92704
rect 354030 92692 354036 92704
rect 354088 92692 354094 92744
rect 356054 92488 356060 92540
rect 356112 92528 356118 92540
rect 356514 92528 356520 92540
rect 356112 92500 356520 92528
rect 356112 92488 356118 92500
rect 356514 92488 356520 92500
rect 356572 92488 356578 92540
rect 395338 92488 395344 92540
rect 395396 92528 395402 92540
rect 396074 92528 396080 92540
rect 395396 92500 396080 92528
rect 395396 92488 395402 92500
rect 396074 92488 396080 92500
rect 396132 92488 396138 92540
rect 396718 92488 396724 92540
rect 396776 92528 396782 92540
rect 399570 92528 399576 92540
rect 396776 92500 399576 92528
rect 396776 92488 396782 92500
rect 399570 92488 399576 92500
rect 399628 92488 399634 92540
rect 406378 92488 406384 92540
rect 406436 92528 406442 92540
rect 408494 92528 408500 92540
rect 406436 92500 408500 92528
rect 406436 92488 406442 92500
rect 408494 92488 408500 92500
rect 408552 92488 408558 92540
rect 88978 92420 88984 92472
rect 89036 92460 89042 92472
rect 164878 92460 164884 92472
rect 89036 92432 164884 92460
rect 89036 92420 89042 92432
rect 164878 92420 164884 92432
rect 164936 92420 164942 92472
rect 192478 92420 192484 92472
rect 192536 92460 192542 92472
rect 357434 92460 357440 92472
rect 192536 92432 357440 92460
rect 192536 92420 192542 92432
rect 357434 92420 357440 92432
rect 357492 92420 357498 92472
rect 202230 92352 202236 92404
rect 202288 92392 202294 92404
rect 281626 92392 281632 92404
rect 202288 92364 281632 92392
rect 202288 92352 202294 92364
rect 281626 92352 281632 92364
rect 281684 92352 281690 92404
rect 337470 92352 337476 92404
rect 337528 92392 337534 92404
rect 394694 92392 394700 92404
rect 337528 92364 394700 92392
rect 337528 92352 337534 92364
rect 394694 92352 394700 92364
rect 394752 92352 394758 92404
rect 98178 92284 98184 92336
rect 98236 92324 98242 92336
rect 118694 92324 118700 92336
rect 98236 92296 118700 92324
rect 98236 92284 98242 92296
rect 118694 92284 118700 92296
rect 118752 92284 118758 92336
rect 133138 92284 133144 92336
rect 133196 92324 133202 92336
rect 169018 92324 169024 92336
rect 133196 92296 169024 92324
rect 133196 92284 133202 92296
rect 169018 92284 169024 92296
rect 169076 92284 169082 92336
rect 178678 92284 178684 92336
rect 178736 92324 178742 92336
rect 281718 92324 281724 92336
rect 178736 92296 281724 92324
rect 178736 92284 178742 92296
rect 281718 92284 281724 92296
rect 281776 92284 281782 92336
rect 298738 92284 298744 92336
rect 298796 92324 298802 92336
rect 352006 92324 352012 92336
rect 298796 92296 352012 92324
rect 298796 92284 298802 92296
rect 352006 92284 352012 92296
rect 352064 92284 352070 92336
rect 125962 92216 125968 92268
rect 126020 92256 126026 92268
rect 195422 92256 195428 92268
rect 126020 92228 195428 92256
rect 126020 92216 126026 92228
rect 195422 92216 195428 92228
rect 195480 92216 195486 92268
rect 216214 92216 216220 92268
rect 216272 92256 216278 92268
rect 280338 92256 280344 92268
rect 216272 92228 280344 92256
rect 216272 92216 216278 92228
rect 280338 92216 280344 92228
rect 280396 92216 280402 92268
rect 115842 92148 115848 92200
rect 115900 92188 115906 92200
rect 130378 92188 130384 92200
rect 115900 92160 130384 92188
rect 115900 92148 115906 92160
rect 130378 92148 130384 92160
rect 130436 92148 130442 92200
rect 136082 92148 136088 92200
rect 136140 92188 136146 92200
rect 191190 92188 191196 92200
rect 136140 92160 191196 92188
rect 136140 92148 136146 92160
rect 191190 92148 191196 92160
rect 191248 92148 191254 92200
rect 152090 92080 152096 92132
rect 152148 92120 152154 92132
rect 189718 92120 189724 92132
rect 152148 92092 189724 92120
rect 152148 92080 152154 92092
rect 189718 92080 189724 92092
rect 189776 92080 189782 92132
rect 84378 92012 84384 92064
rect 84436 92052 84442 92064
rect 203702 92052 203708 92064
rect 84436 92024 203708 92052
rect 84436 92012 84442 92024
rect 203702 92012 203708 92024
rect 203760 92012 203766 92064
rect 352006 91740 352012 91792
rect 352064 91780 352070 91792
rect 352742 91780 352748 91792
rect 352064 91752 352748 91780
rect 352064 91740 352070 91752
rect 352742 91740 352748 91752
rect 352800 91740 352806 91792
rect 74810 91060 74816 91112
rect 74868 91100 74874 91112
rect 135898 91100 135904 91112
rect 74868 91072 135904 91100
rect 74868 91060 74874 91072
rect 135898 91060 135904 91072
rect 135956 91060 135962 91112
rect 105906 90992 105912 91044
rect 105964 91032 105970 91044
rect 193858 91032 193864 91044
rect 105964 91004 193864 91032
rect 105964 90992 105970 91004
rect 193858 90992 193864 91004
rect 193916 90992 193922 91044
rect 316862 90992 316868 91044
rect 316920 91032 316926 91044
rect 391934 91032 391940 91044
rect 316920 91004 391940 91032
rect 316920 90992 316926 91004
rect 391934 90992 391940 91004
rect 391992 90992 391998 91044
rect 111610 90924 111616 90976
rect 111668 90964 111674 90976
rect 166350 90964 166356 90976
rect 111668 90936 166356 90964
rect 111668 90924 111674 90936
rect 166350 90924 166356 90936
rect 166408 90924 166414 90976
rect 126514 90856 126520 90908
rect 126572 90896 126578 90908
rect 180334 90896 180340 90908
rect 126572 90868 180340 90896
rect 126572 90856 126578 90868
rect 180334 90856 180340 90868
rect 180392 90856 180398 90908
rect 122834 90788 122840 90840
rect 122892 90828 122898 90840
rect 170674 90828 170680 90840
rect 122892 90800 170680 90828
rect 122892 90788 122898 90800
rect 170674 90788 170680 90800
rect 170732 90788 170738 90840
rect 124582 90720 124588 90772
rect 124640 90760 124646 90772
rect 171870 90760 171876 90772
rect 124640 90732 171876 90760
rect 124640 90720 124646 90732
rect 171870 90720 171876 90732
rect 171928 90720 171934 90772
rect 151538 90652 151544 90704
rect 151596 90692 151602 90704
rect 198090 90692 198096 90704
rect 151596 90664 198096 90692
rect 151596 90652 151602 90664
rect 198090 90652 198096 90664
rect 198148 90652 198154 90704
rect 298094 90312 298100 90364
rect 298152 90352 298158 90364
rect 366634 90352 366640 90364
rect 298152 90324 366640 90352
rect 298152 90312 298158 90324
rect 366634 90312 366640 90324
rect 366692 90312 366698 90364
rect 65978 89632 65984 89684
rect 66036 89672 66042 89684
rect 210602 89672 210608 89684
rect 66036 89644 210608 89672
rect 66036 89632 66042 89644
rect 210602 89632 210608 89644
rect 210660 89632 210666 89684
rect 100570 89564 100576 89616
rect 100628 89604 100634 89616
rect 207750 89604 207756 89616
rect 100628 89576 207756 89604
rect 100628 89564 100634 89576
rect 207750 89564 207756 89576
rect 207808 89564 207814 89616
rect 102870 89496 102876 89548
rect 102928 89536 102934 89548
rect 198182 89536 198188 89548
rect 102928 89508 198188 89536
rect 102928 89496 102934 89508
rect 198182 89496 198188 89508
rect 198240 89496 198246 89548
rect 115842 89428 115848 89480
rect 115900 89468 115906 89480
rect 178954 89468 178960 89480
rect 115900 89440 178960 89468
rect 115900 89428 115906 89440
rect 178954 89428 178960 89440
rect 179012 89428 179018 89480
rect 132402 89360 132408 89412
rect 132460 89400 132466 89412
rect 171778 89400 171784 89412
rect 132460 89372 171784 89400
rect 132460 89360 132466 89372
rect 171778 89360 171784 89372
rect 171836 89360 171842 89412
rect 291838 89020 291844 89072
rect 291896 89060 291902 89072
rect 327074 89060 327080 89072
rect 291896 89032 327080 89060
rect 291896 89020 291902 89032
rect 327074 89020 327080 89032
rect 327132 89060 327138 89072
rect 355318 89060 355324 89072
rect 327132 89032 355324 89060
rect 327132 89020 327138 89032
rect 355318 89020 355324 89032
rect 355376 89020 355382 89072
rect 198090 88952 198096 89004
rect 198148 88992 198154 89004
rect 265894 88992 265900 89004
rect 198148 88964 265900 88992
rect 198148 88952 198154 88964
rect 265894 88952 265900 88964
rect 265952 88952 265958 89004
rect 300210 88952 300216 89004
rect 300268 88992 300274 89004
rect 351914 88992 351920 89004
rect 300268 88964 351920 88992
rect 300268 88952 300274 88964
rect 351914 88952 351920 88964
rect 351972 88992 351978 89004
rect 388162 88992 388168 89004
rect 351972 88964 388168 88992
rect 351972 88952 351978 88964
rect 388162 88952 388168 88964
rect 388220 88952 388226 89004
rect 411254 88952 411260 89004
rect 411312 88992 411318 89004
rect 412266 88992 412272 89004
rect 411312 88964 412272 88992
rect 411312 88952 411318 88964
rect 412266 88952 412272 88964
rect 412324 88952 412330 89004
rect 101858 88272 101864 88324
rect 101916 88312 101922 88324
rect 181530 88312 181536 88324
rect 101916 88284 181536 88312
rect 101916 88272 101922 88284
rect 181530 88272 181536 88284
rect 181588 88272 181594 88324
rect 230566 88272 230572 88324
rect 230624 88312 230630 88324
rect 233970 88312 233976 88324
rect 230624 88284 233976 88312
rect 230624 88272 230630 88284
rect 233970 88272 233976 88284
rect 234028 88272 234034 88324
rect 85850 88204 85856 88256
rect 85908 88244 85914 88256
rect 166442 88244 166448 88256
rect 85908 88216 166448 88244
rect 85908 88204 85914 88216
rect 166442 88204 166448 88216
rect 166500 88204 166506 88256
rect 107194 88136 107200 88188
rect 107252 88176 107258 88188
rect 169202 88176 169208 88188
rect 107252 88148 169208 88176
rect 107252 88136 107258 88148
rect 169202 88136 169208 88148
rect 169260 88136 169266 88188
rect 117130 88068 117136 88120
rect 117188 88108 117194 88120
rect 178770 88108 178776 88120
rect 117188 88080 178776 88108
rect 117188 88068 117194 88080
rect 178770 88068 178776 88080
rect 178828 88068 178834 88120
rect 151630 88000 151636 88052
rect 151688 88040 151694 88052
rect 211798 88040 211804 88052
rect 151688 88012 211804 88040
rect 151688 88000 151694 88012
rect 211798 88000 211804 88012
rect 211856 88000 211862 88052
rect 135070 87932 135076 87984
rect 135128 87972 135134 87984
rect 167638 87972 167644 87984
rect 135128 87944 167644 87972
rect 135128 87932 135134 87944
rect 167638 87932 167644 87944
rect 167696 87932 167702 87984
rect 197998 87592 198004 87644
rect 198056 87632 198062 87644
rect 302234 87632 302240 87644
rect 198056 87604 302240 87632
rect 198056 87592 198062 87604
rect 302234 87592 302240 87604
rect 302292 87632 302298 87644
rect 365714 87632 365720 87644
rect 302292 87604 365720 87632
rect 302292 87592 302298 87604
rect 365714 87592 365720 87604
rect 365772 87592 365778 87644
rect 67726 86912 67732 86964
rect 67784 86952 67790 86964
rect 214926 86952 214932 86964
rect 67784 86924 214932 86952
rect 67784 86912 67790 86924
rect 214926 86912 214932 86924
rect 214984 86912 214990 86964
rect 439498 86912 439504 86964
rect 439556 86952 439562 86964
rect 580166 86952 580172 86964
rect 439556 86924 580172 86952
rect 439556 86912 439562 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 100662 86844 100668 86896
rect 100720 86884 100726 86896
rect 188522 86884 188528 86896
rect 100720 86856 188528 86884
rect 100720 86844 100726 86856
rect 188522 86844 188528 86856
rect 188580 86844 188586 86896
rect 128170 86776 128176 86828
rect 128228 86816 128234 86828
rect 210418 86816 210424 86828
rect 128228 86788 210424 86816
rect 128228 86776 128234 86788
rect 210418 86776 210424 86788
rect 210476 86776 210482 86828
rect 88058 86708 88064 86760
rect 88116 86748 88122 86760
rect 169294 86748 169300 86760
rect 88116 86720 169300 86748
rect 88116 86708 88122 86720
rect 169294 86708 169300 86720
rect 169352 86708 169358 86760
rect 110138 86640 110144 86692
rect 110196 86680 110202 86692
rect 177574 86680 177580 86692
rect 110196 86652 177580 86680
rect 110196 86640 110202 86652
rect 177574 86640 177580 86652
rect 177632 86640 177638 86692
rect 115750 86572 115756 86624
rect 115808 86612 115814 86624
rect 173434 86612 173440 86624
rect 115808 86584 173440 86612
rect 115808 86572 115814 86584
rect 173434 86572 173440 86584
rect 173492 86572 173498 86624
rect 276014 86232 276020 86284
rect 276072 86272 276078 86284
rect 342346 86272 342352 86284
rect 276072 86244 342352 86272
rect 276072 86232 276078 86244
rect 342346 86232 342352 86244
rect 342404 86232 342410 86284
rect 345014 86232 345020 86284
rect 345072 86272 345078 86284
rect 427998 86272 428004 86284
rect 345072 86244 428004 86272
rect 345072 86232 345078 86244
rect 427998 86232 428004 86244
rect 428056 86232 428062 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 46934 85524 46940 85536
rect 3200 85496 46940 85524
rect 3200 85484 3206 85496
rect 46934 85484 46940 85496
rect 46992 85484 46998 85536
rect 67542 85484 67548 85536
rect 67600 85524 67606 85536
rect 200850 85524 200856 85536
rect 67600 85496 200856 85524
rect 67600 85484 67606 85496
rect 200850 85484 200856 85496
rect 200908 85484 200914 85536
rect 304258 85484 304264 85536
rect 304316 85524 304322 85536
rect 304994 85524 305000 85536
rect 304316 85496 305000 85524
rect 304316 85484 304322 85496
rect 304994 85484 305000 85496
rect 305052 85484 305058 85536
rect 90634 85416 90640 85468
rect 90692 85456 90698 85468
rect 213454 85456 213460 85468
rect 90692 85428 213460 85456
rect 90692 85416 90698 85428
rect 213454 85416 213460 85428
rect 213512 85416 213518 85468
rect 118234 85348 118240 85400
rect 118292 85388 118298 85400
rect 213362 85388 213368 85400
rect 118292 85360 213368 85388
rect 118292 85348 118298 85360
rect 213362 85348 213368 85360
rect 213420 85348 213426 85400
rect 92290 85280 92296 85332
rect 92348 85320 92354 85332
rect 170398 85320 170404 85332
rect 92348 85292 170404 85320
rect 92348 85280 92354 85292
rect 170398 85280 170404 85292
rect 170456 85280 170462 85332
rect 125410 85212 125416 85264
rect 125468 85252 125474 85264
rect 176102 85252 176108 85264
rect 125468 85224 176108 85252
rect 125468 85212 125474 85224
rect 176102 85212 176108 85224
rect 176160 85212 176166 85264
rect 304994 84804 305000 84856
rect 305052 84844 305058 84856
rect 404354 84844 404360 84856
rect 305052 84816 404360 84844
rect 305052 84804 305058 84816
rect 404354 84804 404360 84816
rect 404412 84804 404418 84856
rect 67450 84124 67456 84176
rect 67508 84164 67514 84176
rect 214834 84164 214840 84176
rect 67508 84136 214840 84164
rect 67508 84124 67514 84136
rect 214834 84124 214840 84136
rect 214892 84124 214898 84176
rect 122650 84056 122656 84108
rect 122708 84096 122714 84108
rect 209130 84096 209136 84108
rect 122708 84068 209136 84096
rect 122708 84056 122714 84068
rect 209130 84056 209136 84068
rect 209188 84056 209194 84108
rect 108850 83988 108856 84040
rect 108908 84028 108914 84040
rect 180150 84028 180156 84040
rect 108908 84000 180156 84028
rect 108908 83988 108914 84000
rect 180150 83988 180156 84000
rect 180208 83988 180214 84040
rect 99190 83920 99196 83972
rect 99248 83960 99254 83972
rect 166258 83960 166264 83972
rect 99248 83932 166264 83960
rect 99248 83920 99254 83932
rect 166258 83920 166264 83932
rect 166316 83920 166322 83972
rect 104710 83852 104716 83904
rect 104768 83892 104774 83904
rect 167730 83892 167736 83904
rect 104768 83864 167736 83892
rect 104768 83852 104774 83864
rect 167730 83852 167736 83864
rect 167788 83852 167794 83904
rect 119982 83784 119988 83836
rect 120040 83824 120046 83836
rect 170490 83824 170496 83836
rect 120040 83796 170496 83824
rect 120040 83784 120046 83796
rect 170490 83784 170496 83796
rect 170548 83784 170554 83836
rect 291194 83512 291200 83564
rect 291252 83552 291258 83564
rect 332042 83552 332048 83564
rect 291252 83524 332048 83552
rect 291252 83512 291258 83524
rect 332042 83512 332048 83524
rect 332100 83512 332106 83564
rect 325142 83444 325148 83496
rect 325200 83484 325206 83496
rect 331214 83484 331220 83496
rect 325200 83456 331220 83484
rect 325200 83444 325206 83456
rect 331214 83444 331220 83456
rect 331272 83484 331278 83496
rect 397454 83484 397460 83496
rect 331272 83456 397460 83484
rect 331272 83444 331278 83456
rect 397454 83444 397460 83456
rect 397512 83444 397518 83496
rect 106090 82764 106096 82816
rect 106148 82804 106154 82816
rect 209222 82804 209228 82816
rect 106148 82776 209228 82804
rect 106148 82764 106154 82776
rect 209222 82764 209228 82776
rect 209280 82764 209286 82816
rect 124030 82696 124036 82748
rect 124088 82736 124094 82748
rect 206370 82736 206376 82748
rect 124088 82708 206376 82736
rect 124088 82696 124094 82708
rect 206370 82696 206376 82708
rect 206428 82696 206434 82748
rect 96522 82628 96528 82680
rect 96580 82668 96586 82680
rect 171962 82668 171968 82680
rect 96580 82640 171968 82668
rect 96580 82628 96586 82640
rect 171962 82628 171968 82640
rect 172020 82628 172026 82680
rect 122742 82560 122748 82612
rect 122800 82600 122806 82612
rect 177390 82600 177396 82612
rect 122800 82572 177396 82600
rect 122800 82560 122806 82572
rect 177390 82560 177396 82572
rect 177448 82560 177454 82612
rect 324314 82084 324320 82136
rect 324372 82124 324378 82136
rect 396074 82124 396080 82136
rect 324372 82096 396080 82124
rect 324372 82084 324378 82096
rect 396074 82084 396080 82096
rect 396132 82084 396138 82136
rect 112990 81336 112996 81388
rect 113048 81376 113054 81388
rect 210510 81376 210516 81388
rect 113048 81348 210516 81376
rect 113048 81336 113054 81348
rect 210510 81336 210516 81348
rect 210568 81336 210574 81388
rect 93762 81268 93768 81320
rect 93820 81308 93826 81320
rect 177482 81308 177488 81320
rect 93820 81280 177488 81308
rect 93820 81268 93826 81280
rect 177482 81268 177488 81280
rect 177540 81268 177546 81320
rect 131022 81200 131028 81252
rect 131080 81240 131086 81252
rect 196802 81240 196808 81252
rect 131080 81212 196808 81240
rect 131080 81200 131086 81212
rect 196802 81200 196808 81212
rect 196860 81200 196866 81252
rect 273254 80656 273260 80708
rect 273312 80696 273318 80708
rect 340874 80696 340880 80708
rect 273312 80668 340880 80696
rect 273312 80656 273318 80668
rect 340874 80656 340880 80668
rect 340932 80656 340938 80708
rect 342254 80656 342260 80708
rect 342312 80696 342318 80708
rect 390554 80696 390560 80708
rect 342312 80668 390560 80696
rect 342312 80656 342318 80668
rect 390554 80656 390560 80668
rect 390612 80656 390618 80708
rect 97902 79976 97908 80028
rect 97960 80016 97966 80028
rect 206462 80016 206468 80028
rect 97960 79988 206468 80016
rect 97960 79976 97966 79988
rect 206462 79976 206468 79988
rect 206520 79976 206526 80028
rect 338114 79976 338120 80028
rect 338172 80016 338178 80028
rect 393314 80016 393320 80028
rect 338172 79988 393320 80016
rect 338172 79976 338178 79988
rect 393314 79976 393320 79988
rect 393372 79976 393378 80028
rect 126882 79908 126888 79960
rect 126940 79948 126946 79960
rect 213270 79948 213276 79960
rect 126940 79920 213276 79948
rect 126940 79908 126946 79920
rect 213270 79908 213276 79920
rect 213328 79908 213334 79960
rect 102042 79840 102048 79892
rect 102100 79880 102106 79892
rect 173158 79880 173164 79892
rect 102100 79852 173164 79880
rect 102100 79840 102106 79852
rect 173158 79840 173164 79852
rect 173216 79840 173222 79892
rect 108942 79772 108948 79824
rect 109000 79812 109006 79824
rect 176194 79812 176200 79824
rect 109000 79784 176200 79812
rect 109000 79772 109006 79784
rect 176194 79772 176200 79784
rect 176252 79772 176258 79824
rect 124122 79704 124128 79756
rect 124180 79744 124186 79756
rect 169110 79744 169116 79756
rect 124180 79716 169116 79744
rect 124180 79704 124186 79716
rect 169110 79704 169116 79716
rect 169168 79704 169174 79756
rect 335354 79568 335360 79620
rect 335412 79608 335418 79620
rect 338114 79608 338120 79620
rect 335412 79580 338120 79608
rect 335412 79568 335418 79580
rect 338114 79568 338120 79580
rect 338172 79568 338178 79620
rect 99282 78616 99288 78668
rect 99340 78656 99346 78668
rect 207658 78656 207664 78668
rect 99340 78628 207664 78656
rect 99340 78616 99346 78628
rect 207658 78616 207664 78628
rect 207716 78616 207722 78668
rect 95142 78548 95148 78600
rect 95200 78588 95206 78600
rect 178862 78588 178868 78600
rect 95200 78560 178868 78588
rect 95200 78548 95206 78560
rect 178862 78548 178868 78560
rect 178920 78548 178926 78600
rect 86862 78480 86868 78532
rect 86920 78520 86926 78532
rect 167914 78520 167920 78532
rect 86920 78492 167920 78520
rect 86920 78480 86926 78492
rect 167914 78480 167920 78492
rect 167972 78480 167978 78532
rect 113082 78412 113088 78464
rect 113140 78452 113146 78464
rect 184290 78452 184296 78464
rect 113140 78424 184296 78452
rect 113140 78412 113146 78424
rect 184290 78412 184296 78424
rect 184348 78412 184354 78464
rect 135898 78344 135904 78396
rect 135956 78384 135962 78396
rect 204990 78384 204996 78396
rect 135956 78356 204996 78384
rect 135956 78344 135962 78356
rect 204990 78344 204996 78356
rect 205048 78344 205054 78396
rect 278038 77936 278044 77988
rect 278096 77976 278102 77988
rect 372614 77976 372620 77988
rect 278096 77948 372620 77976
rect 278096 77936 278102 77948
rect 372614 77936 372620 77948
rect 372672 77936 372678 77988
rect 110230 77188 110236 77240
rect 110288 77228 110294 77240
rect 181438 77228 181444 77240
rect 110288 77200 181444 77228
rect 110288 77188 110294 77200
rect 181438 77188 181444 77200
rect 181496 77188 181502 77240
rect 110322 77120 110328 77172
rect 110380 77160 110386 77172
rect 173342 77160 173348 77172
rect 110380 77132 173348 77160
rect 110380 77120 110386 77132
rect 173342 77120 173348 77132
rect 173400 77120 173406 77172
rect 122834 76576 122840 76628
rect 122892 76616 122898 76628
rect 254854 76616 254860 76628
rect 122892 76588 254860 76616
rect 122892 76576 122898 76588
rect 254854 76576 254860 76588
rect 254912 76576 254918 76628
rect 37274 76508 37280 76560
rect 37332 76548 37338 76560
rect 240962 76548 240968 76560
rect 37332 76520 240968 76548
rect 37332 76508 37338 76520
rect 240962 76508 240968 76520
rect 241020 76508 241026 76560
rect 314102 76508 314108 76560
rect 314160 76548 314166 76560
rect 328454 76548 328460 76560
rect 314160 76520 328460 76548
rect 314160 76508 314166 76520
rect 328454 76508 328460 76520
rect 328512 76548 328518 76560
rect 395338 76548 395344 76560
rect 328512 76520 395344 76548
rect 328512 76508 328518 76520
rect 395338 76508 395344 76520
rect 395396 76508 395402 76560
rect 59262 75828 59268 75880
rect 59320 75868 59326 75880
rect 202322 75868 202328 75880
rect 59320 75840 202328 75868
rect 59320 75828 59326 75840
rect 202322 75828 202328 75840
rect 202380 75828 202386 75880
rect 317414 75828 317420 75880
rect 317472 75868 317478 75880
rect 322934 75868 322940 75880
rect 317472 75840 322940 75868
rect 317472 75828 317478 75840
rect 322934 75828 322940 75840
rect 322992 75868 322998 75880
rect 396718 75868 396724 75880
rect 322992 75840 396724 75868
rect 322992 75828 322998 75840
rect 396718 75828 396724 75840
rect 396776 75828 396782 75880
rect 104894 75216 104900 75268
rect 104952 75256 104958 75268
rect 256142 75256 256148 75268
rect 104952 75228 256148 75256
rect 104952 75216 104958 75228
rect 256142 75216 256148 75228
rect 256200 75216 256206 75268
rect 11054 75148 11060 75200
rect 11112 75188 11118 75200
rect 260374 75188 260380 75200
rect 11112 75160 260380 75188
rect 11112 75148 11118 75160
rect 260374 75148 260380 75160
rect 260432 75148 260438 75200
rect 269114 75148 269120 75200
rect 269172 75188 269178 75200
rect 318150 75188 318156 75200
rect 269172 75160 318156 75188
rect 269172 75148 269178 75160
rect 318150 75148 318156 75160
rect 318208 75148 318214 75200
rect 75914 73788 75920 73840
rect 75972 73828 75978 73840
rect 249242 73828 249248 73840
rect 75972 73800 249248 73828
rect 75972 73788 75978 73800
rect 249242 73788 249248 73800
rect 249300 73788 249306 73840
rect 314654 73788 314660 73840
rect 314712 73828 314718 73840
rect 400214 73828 400220 73840
rect 314712 73800 400220 73828
rect 314712 73788 314718 73800
rect 400214 73788 400220 73800
rect 400272 73788 400278 73840
rect 349982 73108 349988 73160
rect 350040 73148 350046 73160
rect 579982 73148 579988 73160
rect 350040 73120 579988 73148
rect 350040 73108 350046 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 64414 72428 64420 72480
rect 64472 72468 64478 72480
rect 311802 72468 311808 72480
rect 64472 72440 311808 72468
rect 64472 72428 64478 72440
rect 311802 72428 311808 72440
rect 311860 72428 311866 72480
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 57882 71720 57888 71732
rect 3476 71692 57888 71720
rect 3476 71680 3482 71692
rect 57882 71680 57888 71692
rect 57940 71720 57946 71732
rect 436094 71720 436100 71732
rect 57940 71692 436100 71720
rect 57940 71680 57946 71692
rect 436094 71680 436100 71692
rect 436152 71680 436158 71732
rect 60734 71000 60740 71052
rect 60792 71040 60798 71052
rect 253382 71040 253388 71052
rect 60792 71012 253388 71040
rect 60792 71000 60798 71012
rect 253382 71000 253388 71012
rect 253440 71000 253446 71052
rect 110414 69708 110420 69760
rect 110472 69748 110478 69760
rect 247770 69748 247776 69760
rect 110472 69720 247776 69748
rect 110472 69708 110478 69720
rect 247770 69708 247776 69720
rect 247828 69708 247834 69760
rect 97994 69640 98000 69692
rect 98052 69680 98058 69692
rect 263134 69680 263140 69692
rect 98052 69652 263140 69680
rect 98052 69640 98058 69652
rect 263134 69640 263140 69652
rect 263192 69640 263198 69692
rect 311158 69640 311164 69692
rect 311216 69680 311222 69692
rect 311802 69680 311808 69692
rect 311216 69652 311808 69680
rect 311216 69640 311222 69652
rect 311802 69640 311808 69652
rect 311860 69680 311866 69692
rect 401594 69680 401600 69692
rect 311860 69652 401600 69680
rect 311860 69640 311866 69652
rect 401594 69640 401600 69652
rect 401652 69640 401658 69692
rect 74534 68280 74540 68332
rect 74592 68320 74598 68332
rect 245102 68320 245108 68332
rect 74592 68292 245108 68320
rect 74592 68280 74598 68292
rect 245102 68280 245108 68292
rect 245160 68280 245166 68332
rect 322198 68280 322204 68332
rect 322256 68320 322262 68332
rect 402974 68320 402980 68332
rect 322256 68292 402980 68320
rect 322256 68280 322262 68292
rect 402974 68280 402980 68292
rect 403032 68280 403038 68332
rect 81434 66920 81440 66972
rect 81492 66960 81498 66972
rect 236822 66960 236828 66972
rect 81492 66932 236828 66960
rect 81492 66920 81498 66932
rect 236822 66920 236828 66932
rect 236880 66920 236886 66972
rect 6914 66852 6920 66904
rect 6972 66892 6978 66904
rect 226978 66892 226984 66904
rect 6972 66864 226984 66892
rect 6972 66852 6978 66864
rect 226978 66852 226984 66864
rect 227036 66852 227042 66904
rect 299658 66852 299664 66904
rect 299716 66892 299722 66904
rect 399478 66892 399484 66904
rect 299716 66864 399484 66892
rect 299716 66852 299722 66864
rect 399478 66852 399484 66864
rect 399536 66852 399542 66904
rect 296714 66172 296720 66224
rect 296772 66212 296778 66224
rect 297358 66212 297364 66224
rect 296772 66184 297364 66212
rect 296772 66172 296778 66184
rect 297358 66172 297364 66184
rect 297416 66212 297422 66224
rect 407114 66212 407120 66224
rect 297416 66184 407120 66212
rect 297416 66172 297422 66184
rect 407114 66172 407120 66184
rect 407172 66172 407178 66224
rect 46934 65560 46940 65612
rect 46992 65600 46998 65612
rect 222838 65600 222844 65612
rect 46992 65572 222844 65600
rect 46992 65560 46998 65572
rect 222838 65560 222844 65572
rect 222896 65560 222902 65612
rect 85574 65492 85580 65544
rect 85632 65532 85638 65544
rect 261662 65532 261668 65544
rect 85632 65504 261668 65532
rect 85632 65492 85638 65504
rect 261662 65492 261668 65504
rect 261720 65492 261726 65544
rect 215938 64268 215944 64320
rect 215996 64308 216002 64320
rect 295334 64308 295340 64320
rect 215996 64280 295340 64308
rect 215996 64268 216002 64280
rect 295334 64268 295340 64280
rect 295392 64308 295398 64320
rect 295392 64280 296714 64308
rect 295392 64268 295398 64280
rect 87598 64200 87604 64252
rect 87656 64240 87662 64252
rect 265802 64240 265808 64252
rect 87656 64212 265808 64240
rect 87656 64200 87662 64212
rect 265802 64200 265808 64212
rect 265860 64200 265866 64252
rect 51166 64132 51172 64184
rect 51224 64172 51230 64184
rect 242434 64172 242440 64184
rect 51224 64144 242440 64172
rect 51224 64132 51230 64144
rect 242434 64132 242440 64144
rect 242492 64132 242498 64184
rect 296686 64172 296714 64280
rect 409874 64172 409880 64184
rect 296686 64144 409880 64172
rect 409874 64132 409880 64144
rect 409932 64132 409938 64184
rect 88334 62840 88340 62892
rect 88392 62880 88398 62892
rect 254762 62880 254768 62892
rect 88392 62852 254768 62880
rect 88392 62840 88398 62852
rect 254762 62840 254768 62852
rect 254820 62840 254826 62892
rect 57974 62772 57980 62824
rect 58032 62812 58038 62824
rect 264514 62812 264520 62824
rect 58032 62784 264520 62812
rect 58032 62772 58038 62784
rect 264514 62772 264520 62784
rect 264572 62772 264578 62824
rect 286318 62772 286324 62824
rect 286376 62812 286382 62824
rect 411346 62812 411352 62824
rect 286376 62784 411352 62812
rect 286376 62772 286382 62784
rect 411346 62772 411352 62784
rect 411404 62772 411410 62824
rect 92474 61412 92480 61464
rect 92532 61452 92538 61464
rect 246574 61452 246580 61464
rect 92532 61424 246580 61452
rect 92532 61412 92538 61424
rect 246574 61412 246580 61424
rect 246632 61412 246638 61464
rect 64874 61344 64880 61396
rect 64932 61384 64938 61396
rect 239582 61384 239588 61396
rect 64932 61356 239588 61384
rect 64932 61344 64938 61356
rect 239582 61344 239588 61356
rect 239640 61344 239646 61396
rect 267090 61344 267096 61396
rect 267148 61384 267154 61396
rect 280246 61384 280252 61396
rect 267148 61356 280252 61384
rect 267148 61344 267154 61356
rect 280246 61344 280252 61356
rect 280304 61384 280310 61396
rect 412634 61384 412640 61396
rect 280304 61356 412640 61384
rect 280304 61344 280310 61356
rect 412634 61344 412640 61356
rect 412692 61344 412698 61396
rect 113174 60120 113180 60172
rect 113232 60160 113238 60172
rect 243630 60160 243636 60172
rect 113232 60132 243636 60160
rect 113232 60120 113238 60132
rect 243630 60120 243636 60132
rect 243688 60120 243694 60172
rect 69014 60052 69020 60104
rect 69072 60092 69078 60104
rect 261754 60092 261760 60104
rect 69072 60064 261760 60092
rect 69072 60052 69078 60064
rect 261754 60052 261760 60064
rect 261812 60052 261818 60104
rect 4246 59984 4252 60036
rect 4304 60024 4310 60036
rect 228358 60024 228364 60036
rect 4304 59996 228364 60024
rect 4304 59984 4310 59996
rect 228358 59984 228364 59996
rect 228416 59984 228422 60036
rect 276658 59984 276664 60036
rect 276716 60024 276722 60036
rect 414014 60024 414020 60036
rect 276716 59996 414020 60024
rect 276716 59984 276722 59996
rect 414014 59984 414020 59996
rect 414072 59984 414078 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 51074 59344 51080 59356
rect 3108 59316 51080 59344
rect 3108 59304 3114 59316
rect 51074 59304 51080 59316
rect 51132 59304 51138 59356
rect 111794 58692 111800 58744
rect 111852 58732 111858 58744
rect 264422 58732 264428 58744
rect 111852 58704 264428 58732
rect 111852 58692 111858 58704
rect 264422 58692 264428 58704
rect 264480 58692 264486 58744
rect 71774 58624 71780 58676
rect 71832 58664 71838 58676
rect 245194 58664 245200 58676
rect 71832 58636 245200 58664
rect 71832 58624 71838 58636
rect 245194 58624 245200 58636
rect 245252 58624 245258 58676
rect 267182 58624 267188 58676
rect 267240 58664 267246 58676
rect 271874 58664 271880 58676
rect 267240 58636 271880 58664
rect 267240 58624 267246 58636
rect 271874 58624 271880 58636
rect 271932 58664 271938 58676
rect 415394 58664 415400 58676
rect 271932 58636 415400 58664
rect 271932 58624 271938 58636
rect 415394 58624 415400 58636
rect 415452 58624 415458 58676
rect 85666 57264 85672 57316
rect 85724 57304 85730 57316
rect 240870 57304 240876 57316
rect 85724 57276 240876 57304
rect 85724 57264 85730 57276
rect 240870 57264 240876 57276
rect 240928 57264 240934 57316
rect 13814 57196 13820 57248
rect 13872 57236 13878 57248
rect 252002 57236 252008 57248
rect 13872 57208 252008 57236
rect 13872 57196 13878 57208
rect 252002 57196 252008 57208
rect 252060 57196 252066 57248
rect 268378 57196 268384 57248
rect 268436 57236 268442 57248
rect 416774 57236 416780 57248
rect 268436 57208 416780 57236
rect 268436 57196 268442 57208
rect 416774 57196 416780 57208
rect 416832 57196 416838 57248
rect 124214 55972 124220 56024
rect 124272 56012 124278 56024
rect 257430 56012 257436 56024
rect 124272 55984 257436 56012
rect 124272 55972 124278 55984
rect 257430 55972 257436 55984
rect 257488 55972 257494 56024
rect 52454 55904 52460 55956
rect 52512 55944 52518 55956
rect 258902 55944 258908 55956
rect 52512 55916 258908 55944
rect 52512 55904 52518 55916
rect 258902 55904 258908 55916
rect 258960 55904 258966 55956
rect 2774 55836 2780 55888
rect 2832 55876 2838 55888
rect 229922 55876 229928 55888
rect 2832 55848 229928 55876
rect 2832 55836 2838 55848
rect 229922 55836 229928 55848
rect 229980 55836 229986 55888
rect 264422 55836 264428 55888
rect 264480 55876 264486 55888
rect 419534 55876 419540 55888
rect 264480 55848 419540 55876
rect 264480 55836 264486 55848
rect 419534 55836 419540 55848
rect 419592 55836 419598 55888
rect 60826 54544 60832 54596
rect 60884 54584 60890 54596
rect 256234 54584 256240 54596
rect 60884 54556 256240 54584
rect 60884 54544 60890 54556
rect 256234 54544 256240 54556
rect 256292 54544 256298 54596
rect 15194 54476 15200 54528
rect 15252 54516 15258 54528
rect 235350 54516 235356 54528
rect 15252 54488 235356 54516
rect 15252 54476 15258 54488
rect 235350 54476 235356 54488
rect 235408 54476 235414 54528
rect 254578 54476 254584 54528
rect 254636 54516 254642 54528
rect 422294 54516 422300 54528
rect 254636 54488 422300 54516
rect 254636 54476 254642 54488
rect 422294 54476 422300 54488
rect 422352 54476 422358 54528
rect 177298 53184 177304 53236
rect 177356 53224 177362 53236
rect 251174 53224 251180 53236
rect 177356 53196 251180 53224
rect 177356 53184 177362 53196
rect 251174 53184 251180 53196
rect 251232 53224 251238 53236
rect 251232 53196 267734 53224
rect 251232 53184 251238 53196
rect 107654 53116 107660 53168
rect 107712 53156 107718 53168
rect 260282 53156 260288 53168
rect 107712 53128 260288 53156
rect 107712 53116 107718 53128
rect 260282 53116 260288 53128
rect 260340 53116 260346 53168
rect 30374 53048 30380 53100
rect 30432 53088 30438 53100
rect 247862 53088 247868 53100
rect 30432 53060 247868 53088
rect 30432 53048 30438 53060
rect 247862 53048 247868 53060
rect 247920 53048 247926 53100
rect 267706 53088 267734 53196
rect 423674 53088 423680 53100
rect 267706 53060 423680 53088
rect 423674 53048 423680 53060
rect 423732 53048 423738 53100
rect 118694 51756 118700 51808
rect 118752 51796 118758 51808
rect 249150 51796 249156 51808
rect 118752 51768 249156 51796
rect 118752 51756 118758 51768
rect 249150 51756 249156 51768
rect 249208 51756 249214 51808
rect 425054 51796 425060 51808
rect 258046 51768 425060 51796
rect 17954 51688 17960 51740
rect 18012 51728 18018 51740
rect 18012 51700 238754 51728
rect 18012 51688 18018 51700
rect 238726 51660 238754 51700
rect 248506 51688 248512 51740
rect 248564 51728 248570 51740
rect 258046 51728 258074 51768
rect 425054 51756 425060 51768
rect 425112 51756 425118 51808
rect 248564 51700 258074 51728
rect 248564 51688 248570 51700
rect 252094 51660 252100 51672
rect 238726 51632 252100 51660
rect 252094 51620 252100 51632
rect 252152 51620 252158 51672
rect 313274 50396 313280 50448
rect 313332 50436 313338 50448
rect 360194 50436 360200 50448
rect 313332 50408 360200 50436
rect 313332 50396 313338 50408
rect 360194 50396 360200 50408
rect 360252 50396 360258 50448
rect 19334 50328 19340 50380
rect 19392 50368 19398 50380
rect 250530 50368 250536 50380
rect 19392 50340 250536 50368
rect 19392 50328 19398 50340
rect 250530 50328 250536 50340
rect 250588 50328 250594 50380
rect 259454 50328 259460 50380
rect 259512 50368 259518 50380
rect 314010 50368 314016 50380
rect 259512 50340 314016 50368
rect 259512 50328 259518 50340
rect 314010 50328 314016 50340
rect 314068 50328 314074 50380
rect 347774 50328 347780 50380
rect 347832 50368 347838 50380
rect 432046 50368 432052 50380
rect 347832 50340 432052 50368
rect 347832 50328 347838 50340
rect 432046 50328 432052 50340
rect 432104 50328 432110 50380
rect 96614 49036 96620 49088
rect 96672 49076 96678 49088
rect 234062 49076 234068 49088
rect 96672 49048 234068 49076
rect 96672 49036 96678 49048
rect 234062 49036 234068 49048
rect 234120 49036 234126 49088
rect 309226 49036 309232 49088
rect 309284 49076 309290 49088
rect 361574 49076 361580 49088
rect 309284 49048 361580 49076
rect 309284 49036 309290 49048
rect 361574 49036 361580 49048
rect 361632 49036 361638 49088
rect 56594 48968 56600 49020
rect 56652 49008 56658 49020
rect 258810 49008 258816 49020
rect 56652 48980 258816 49008
rect 56652 48968 56658 48980
rect 258810 48968 258816 48980
rect 258868 48968 258874 49020
rect 340138 48968 340144 49020
rect 340196 49008 340202 49020
rect 394694 49008 394700 49020
rect 340196 48980 394700 49008
rect 340196 48968 340202 48980
rect 394694 48968 394700 48980
rect 394752 48968 394758 49020
rect 93854 47608 93860 47660
rect 93912 47648 93918 47660
rect 263042 47648 263048 47660
rect 93912 47620 263048 47648
rect 93912 47608 93918 47620
rect 263042 47608 263048 47620
rect 263100 47608 263106 47660
rect 44174 47540 44180 47592
rect 44232 47580 44238 47592
rect 242250 47580 242256 47592
rect 44232 47552 242256 47580
rect 44232 47540 44238 47552
rect 242250 47540 242256 47552
rect 242308 47540 242314 47592
rect 302878 47540 302884 47592
rect 302936 47580 302942 47592
rect 364334 47580 364340 47592
rect 302936 47552 364340 47580
rect 302936 47540 302942 47552
rect 364334 47540 364340 47552
rect 364392 47540 364398 47592
rect 464338 46860 464344 46912
rect 464396 46900 464402 46912
rect 580166 46900 580172 46912
rect 464396 46872 580172 46900
rect 464396 46860 464402 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 117314 46316 117320 46368
rect 117372 46356 117378 46368
rect 238018 46356 238024 46368
rect 117372 46328 238024 46356
rect 117372 46316 117378 46328
rect 238018 46316 238024 46328
rect 238076 46316 238082 46368
rect 106274 46248 106280 46300
rect 106332 46288 106338 46300
rect 229830 46288 229836 46300
rect 106332 46260 229836 46288
rect 106332 46248 106338 46260
rect 229830 46248 229836 46260
rect 229888 46248 229894 46300
rect 244274 46248 244280 46300
rect 244332 46288 244338 46300
rect 426526 46288 426532 46300
rect 244332 46260 426532 46288
rect 244332 46248 244338 46260
rect 426526 46248 426532 46260
rect 426584 46248 426590 46300
rect 40034 46180 40040 46232
rect 40092 46220 40098 46232
rect 253474 46220 253480 46232
rect 40092 46192 253480 46220
rect 40092 46180 40098 46192
rect 253474 46180 253480 46192
rect 253532 46180 253538 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 25498 45540 25504 45552
rect 3476 45512 25504 45540
rect 3476 45500 3482 45512
rect 25498 45500 25504 45512
rect 25556 45500 25562 45552
rect 48314 44888 48320 44940
rect 48372 44928 48378 44940
rect 256050 44928 256056 44940
rect 48372 44900 256056 44928
rect 48372 44888 48378 44900
rect 256050 44888 256056 44900
rect 256108 44888 256114 44940
rect 31754 44820 31760 44872
rect 31812 44860 31818 44872
rect 247678 44860 247684 44872
rect 31812 44832 247684 44860
rect 31812 44820 31818 44832
rect 247678 44820 247684 44832
rect 247736 44820 247742 44872
rect 269758 44820 269764 44872
rect 269816 44860 269822 44872
rect 386414 44860 386420 44872
rect 269816 44832 386420 44860
rect 269816 44820 269822 44832
rect 386414 44820 386420 44832
rect 386472 44820 386478 44872
rect 240410 43528 240416 43580
rect 240468 43568 240474 43580
rect 410518 43568 410524 43580
rect 240468 43540 410524 43568
rect 240468 43528 240474 43540
rect 410518 43528 410524 43540
rect 410576 43528 410582 43580
rect 52546 43460 52552 43512
rect 52604 43500 52610 43512
rect 245010 43500 245016 43512
rect 52604 43472 245016 43500
rect 52604 43460 52610 43472
rect 245010 43460 245016 43472
rect 245068 43460 245074 43512
rect 27614 43392 27620 43444
rect 27672 43432 27678 43444
rect 246390 43432 246396 43444
rect 27672 43404 246396 43432
rect 27672 43392 27678 43404
rect 246390 43392 246396 43404
rect 246448 43392 246454 43444
rect 338114 42168 338120 42220
rect 338172 42208 338178 42220
rect 352006 42208 352012 42220
rect 338172 42180 352012 42208
rect 338172 42168 338178 42180
rect 352006 42168 352012 42180
rect 352064 42168 352070 42220
rect 262214 42100 262220 42152
rect 262272 42140 262278 42152
rect 339494 42140 339500 42152
rect 262272 42112 339500 42140
rect 262272 42100 262278 42112
rect 339494 42100 339500 42112
rect 339552 42100 339558 42152
rect 53834 42032 53840 42084
rect 53892 42072 53898 42084
rect 262858 42072 262864 42084
rect 53892 42044 262864 42072
rect 53892 42032 53898 42044
rect 262858 42032 262864 42044
rect 262916 42032 262922 42084
rect 349246 42032 349252 42084
rect 349304 42072 349310 42084
rect 430666 42072 430672 42084
rect 349304 42044 430672 42072
rect 349304 42032 349310 42044
rect 430666 42032 430672 42044
rect 430724 42032 430730 42084
rect 340874 41352 340880 41404
rect 340932 41392 340938 41404
rect 341518 41392 341524 41404
rect 340932 41364 341524 41392
rect 340932 41352 340938 41364
rect 341518 41352 341524 41364
rect 341576 41392 341582 41404
rect 427906 41392 427912 41404
rect 341576 41364 427912 41392
rect 341576 41352 341582 41364
rect 427906 41352 427912 41364
rect 427964 41352 427970 41404
rect 100754 40740 100760 40792
rect 100812 40780 100818 40792
rect 235258 40780 235264 40792
rect 100812 40752 235264 40780
rect 100812 40740 100818 40752
rect 235258 40740 235264 40752
rect 235316 40740 235322 40792
rect 41414 40672 41420 40724
rect 41472 40712 41478 40724
rect 265710 40712 265716 40724
rect 41472 40684 265716 40712
rect 41472 40672 41478 40684
rect 265710 40672 265716 40684
rect 265768 40672 265774 40724
rect 298094 40672 298100 40724
rect 298152 40712 298158 40724
rect 338206 40712 338212 40724
rect 298152 40684 338212 40712
rect 298152 40672 298158 40684
rect 338206 40672 338212 40684
rect 338264 40672 338270 40724
rect 333974 39992 333980 40044
rect 334032 40032 334038 40044
rect 334618 40032 334624 40044
rect 334032 40004 334624 40032
rect 334032 39992 334038 40004
rect 334618 39992 334624 40004
rect 334676 40032 334682 40044
rect 429286 40032 429292 40044
rect 334676 40004 429292 40032
rect 334676 39992 334682 40004
rect 429286 39992 429292 40004
rect 429344 39992 429350 40044
rect 110506 39380 110512 39432
rect 110564 39420 110570 39432
rect 264330 39420 264336 39432
rect 110564 39392 264336 39420
rect 110564 39380 110570 39392
rect 264330 39380 264336 39392
rect 264388 39380 264394 39432
rect 27706 39312 27712 39364
rect 27764 39352 27770 39364
rect 240778 39352 240784 39364
rect 27764 39324 240784 39352
rect 27764 39312 27770 39324
rect 240778 39312 240784 39324
rect 240836 39312 240842 39364
rect 255314 39312 255320 39364
rect 255372 39352 255378 39364
rect 327810 39352 327816 39364
rect 255372 39324 327816 39352
rect 255372 39312 255378 39324
rect 327810 39312 327816 39324
rect 327868 39312 327874 39364
rect 35894 37952 35900 38004
rect 35952 37992 35958 38004
rect 232590 37992 232596 38004
rect 35952 37964 232596 37992
rect 35952 37952 35958 37964
rect 232590 37952 232596 37964
rect 232648 37952 232654 38004
rect 324406 37952 324412 38004
rect 324464 37992 324470 38004
rect 356054 37992 356060 38004
rect 324464 37964 356060 37992
rect 324464 37952 324470 37964
rect 356054 37952 356060 37964
rect 356112 37952 356118 38004
rect 24854 37884 24860 37936
rect 24912 37924 24918 37936
rect 231210 37924 231216 37936
rect 24912 37896 231216 37924
rect 24912 37884 24918 37896
rect 231210 37884 231216 37896
rect 231268 37884 231274 37936
rect 248506 37884 248512 37936
rect 248564 37924 248570 37936
rect 325050 37924 325056 37936
rect 248564 37896 325056 37924
rect 248564 37884 248570 37896
rect 325050 37884 325056 37896
rect 325108 37884 325114 37936
rect 356698 37884 356704 37936
rect 356756 37924 356762 37936
rect 389174 37924 389180 37936
rect 356756 37896 389180 37924
rect 356756 37884 356762 37896
rect 389174 37884 389180 37896
rect 389232 37884 389238 37936
rect 337378 37204 337384 37256
rect 337436 37244 337442 37256
rect 429194 37244 429200 37256
rect 337436 37216 429200 37244
rect 337436 37204 337442 37216
rect 429194 37204 429200 37216
rect 429252 37204 429258 37256
rect 336734 36864 336740 36916
rect 336792 36904 336798 36916
rect 337378 36904 337384 36916
rect 336792 36876 337384 36904
rect 336792 36864 336798 36876
rect 337378 36864 337384 36876
rect 337436 36864 337442 36916
rect 266354 36524 266360 36576
rect 266412 36564 266418 36576
rect 336182 36564 336188 36576
rect 266412 36536 336188 36564
rect 266412 36524 266418 36536
rect 336182 36524 336188 36536
rect 336240 36524 336246 36576
rect 103514 35232 103520 35284
rect 103572 35272 103578 35284
rect 257614 35272 257620 35284
rect 103572 35244 257620 35272
rect 103572 35232 103578 35244
rect 257614 35232 257620 35244
rect 257672 35232 257678 35284
rect 320174 35232 320180 35284
rect 320232 35272 320238 35284
rect 357434 35272 357440 35284
rect 320232 35244 357440 35272
rect 320232 35232 320238 35244
rect 357434 35232 357440 35244
rect 357492 35232 357498 35284
rect 34514 35164 34520 35216
rect 34572 35204 34578 35216
rect 238294 35204 238300 35216
rect 34572 35176 238300 35204
rect 34572 35164 34578 35176
rect 238294 35164 238300 35176
rect 238352 35164 238358 35216
rect 241882 35164 241888 35216
rect 241940 35204 241946 35216
rect 322290 35204 322296 35216
rect 241940 35176 322296 35204
rect 241940 35164 241946 35176
rect 322290 35164 322296 35176
rect 322348 35164 322354 35216
rect 340966 35164 340972 35216
rect 341024 35204 341030 35216
rect 433610 35204 433616 35216
rect 341024 35176 433616 35204
rect 341024 35164 341030 35176
rect 433610 35164 433616 35176
rect 433668 35164 433674 35216
rect 22002 34416 22008 34468
rect 22060 34456 22066 34468
rect 429378 34456 429384 34468
rect 22060 34428 429384 34456
rect 22060 34416 22066 34428
rect 429378 34416 429384 34428
rect 429436 34416 429442 34468
rect 3234 33736 3240 33788
rect 3292 33776 3298 33788
rect 22002 33776 22008 33788
rect 3292 33748 22008 33776
rect 3292 33736 3298 33748
rect 22002 33736 22008 33748
rect 22060 33736 22066 33788
rect 45554 33736 45560 33788
rect 45612 33776 45618 33788
rect 251818 33776 251824 33788
rect 45612 33748 251824 33776
rect 45612 33736 45618 33748
rect 251818 33736 251824 33748
rect 251876 33736 251882 33788
rect 349154 33056 349160 33108
rect 349212 33096 349218 33108
rect 580166 33096 580172 33108
rect 349212 33068 580172 33096
rect 349212 33056 349218 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 174538 32444 174544 32496
rect 174596 32484 174602 32496
rect 244274 32484 244280 32496
rect 174596 32456 244280 32484
rect 174596 32444 174602 32456
rect 244274 32444 244280 32456
rect 244332 32484 244338 32496
rect 244332 32456 248414 32484
rect 244332 32444 244338 32456
rect 55214 32376 55220 32428
rect 55272 32416 55278 32428
rect 239490 32416 239496 32428
rect 55272 32388 239496 32416
rect 55272 32376 55278 32388
rect 239490 32376 239496 32388
rect 239548 32376 239554 32428
rect 248386 32416 248414 32456
rect 316126 32444 316132 32496
rect 316184 32484 316190 32496
rect 358814 32484 358820 32496
rect 316184 32456 358820 32484
rect 316184 32444 316190 32456
rect 358814 32444 358820 32456
rect 358872 32444 358878 32496
rect 320910 32416 320916 32428
rect 248386 32388 320916 32416
rect 320910 32376 320916 32388
rect 320968 32376 320974 32428
rect 95234 31152 95240 31204
rect 95292 31192 95298 31204
rect 236638 31192 236644 31204
rect 95292 31164 236644 31192
rect 95292 31152 95298 31164
rect 236638 31152 236644 31164
rect 236696 31152 236702 31204
rect 121454 31084 121460 31136
rect 121512 31124 121518 31136
rect 264238 31124 264244 31136
rect 121512 31096 264244 31124
rect 121512 31084 121518 31096
rect 264238 31084 264244 31096
rect 264296 31084 264302 31136
rect 22094 31016 22100 31068
rect 22152 31056 22158 31068
rect 251910 31056 251916 31068
rect 22152 31028 251916 31056
rect 22152 31016 22158 31028
rect 251910 31016 251916 31028
rect 251968 31016 251974 31068
rect 294138 31016 294144 31068
rect 294196 31056 294202 31068
rect 367094 31056 367100 31068
rect 294196 31028 367100 31056
rect 294196 31016 294202 31028
rect 367094 31016 367100 31028
rect 367152 31016 367158 31068
rect 204898 29792 204904 29844
rect 204956 29832 204962 29844
rect 283558 29832 283564 29844
rect 204956 29804 283564 29832
rect 204956 29792 204962 29804
rect 283558 29792 283564 29804
rect 283616 29792 283622 29844
rect 200758 29724 200764 29776
rect 200816 29764 200822 29776
rect 200816 29736 277394 29764
rect 200816 29724 200822 29736
rect 114554 29656 114560 29708
rect 114612 29696 114618 29708
rect 238202 29696 238208 29708
rect 114612 29668 238208 29696
rect 114612 29656 114618 29668
rect 238202 29656 238208 29668
rect 238260 29656 238266 29708
rect 59354 29588 59360 29640
rect 59412 29628 59418 29640
rect 244918 29628 244924 29640
rect 59412 29600 244924 29628
rect 59412 29588 59418 29600
rect 244918 29588 244924 29600
rect 244976 29588 244982 29640
rect 277366 29628 277394 29736
rect 288434 29628 288440 29640
rect 277366 29600 288440 29628
rect 288434 29588 288440 29600
rect 288492 29628 288498 29640
rect 368474 29628 368480 29640
rect 288492 29600 368480 29628
rect 288492 29588 288498 29600
rect 368474 29588 368480 29600
rect 368532 29588 368538 29640
rect 196618 28908 196624 28960
rect 196676 28948 196682 28960
rect 276106 28948 276112 28960
rect 196676 28920 276112 28948
rect 196676 28908 196682 28920
rect 276106 28908 276112 28920
rect 276164 28948 276170 28960
rect 276658 28948 276664 28960
rect 276164 28920 276664 28948
rect 276164 28908 276170 28920
rect 276658 28908 276664 28920
rect 276716 28908 276722 28960
rect 73154 28296 73160 28348
rect 73212 28336 73218 28348
rect 253198 28336 253204 28348
rect 73212 28308 253204 28336
rect 73212 28296 73218 28308
rect 253198 28296 253204 28308
rect 253256 28296 253262 28348
rect 44266 28228 44272 28280
rect 44324 28268 44330 28280
rect 231118 28268 231124 28280
rect 44324 28240 231124 28268
rect 44324 28228 44330 28240
rect 231118 28228 231124 28240
rect 231176 28228 231182 28280
rect 287698 28228 287704 28280
rect 287756 28268 287762 28280
rect 369854 28268 369860 28280
rect 287756 28240 369860 28268
rect 287756 28228 287762 28240
rect 369854 28228 369860 28240
rect 369912 28228 369918 28280
rect 206278 26936 206284 26988
rect 206336 26976 206342 26988
rect 206336 26948 259592 26976
rect 206336 26936 206342 26948
rect 259564 26920 259592 26948
rect 28994 26868 29000 26920
rect 29052 26908 29058 26920
rect 258994 26908 259000 26920
rect 29052 26880 259000 26908
rect 29052 26868 29058 26880
rect 258994 26868 259000 26880
rect 259052 26868 259058 26920
rect 259546 26868 259552 26920
rect 259604 26908 259610 26920
rect 379514 26908 379520 26920
rect 259604 26880 379520 26908
rect 259604 26868 259610 26880
rect 379514 26868 379520 26880
rect 379572 26868 379578 26920
rect 33134 25508 33140 25560
rect 33192 25548 33198 25560
rect 257522 25548 257528 25560
rect 33192 25520 257528 25548
rect 33192 25508 33198 25520
rect 257522 25508 257528 25520
rect 257580 25508 257586 25560
rect 289078 25508 289084 25560
rect 289136 25548 289142 25560
rect 373994 25548 374000 25560
rect 289136 25520 374000 25548
rect 289136 25508 289142 25520
rect 373994 25508 374000 25520
rect 374052 25508 374058 25560
rect 252922 24216 252928 24268
rect 252980 24256 252986 24268
rect 380986 24256 380992 24268
rect 252980 24228 380992 24256
rect 252980 24216 252986 24228
rect 380986 24216 380992 24228
rect 381044 24216 381050 24268
rect 36538 24148 36544 24200
rect 36596 24188 36602 24200
rect 263594 24188 263600 24200
rect 36596 24160 263600 24188
rect 36596 24148 36602 24160
rect 263594 24148 263600 24160
rect 263652 24148 263658 24200
rect 11146 24080 11152 24132
rect 11204 24120 11210 24132
rect 254670 24120 254676 24132
rect 11204 24092 254676 24120
rect 11204 24080 11210 24092
rect 254670 24080 254676 24092
rect 254728 24080 254734 24132
rect 115934 22788 115940 22840
rect 115992 22828 115998 22840
rect 224218 22828 224224 22840
rect 115992 22800 224224 22828
rect 115992 22788 115998 22800
rect 224218 22788 224224 22800
rect 224276 22788 224282 22840
rect 26234 22720 26240 22772
rect 26292 22760 26298 22772
rect 246482 22760 246488 22772
rect 26292 22732 246488 22760
rect 26292 22720 26298 22732
rect 246482 22720 246488 22732
rect 246540 22720 246546 22772
rect 383654 22760 383660 22772
rect 248386 22732 383660 22760
rect 245746 22652 245752 22704
rect 245804 22692 245810 22704
rect 248386 22692 248414 22732
rect 383654 22720 383660 22732
rect 383712 22720 383718 22772
rect 245804 22664 248414 22692
rect 245804 22652 245810 22664
rect 203518 21496 203524 21548
rect 203576 21536 203582 21548
rect 203576 21508 267734 21536
rect 203576 21496 203582 21508
rect 89714 21428 89720 21480
rect 89772 21468 89778 21480
rect 261570 21468 261576 21480
rect 89772 21440 261576 21468
rect 89772 21428 89778 21440
rect 261570 21428 261576 21440
rect 261628 21428 261634 21480
rect 67634 21360 67640 21412
rect 67692 21400 67698 21412
rect 243538 21400 243544 21412
rect 67692 21372 243544 21400
rect 67692 21360 67698 21372
rect 243538 21360 243544 21372
rect 243596 21360 243602 21412
rect 267706 21400 267734 21508
rect 270494 21400 270500 21412
rect 267706 21372 270500 21400
rect 270494 21360 270500 21372
rect 270552 21400 270558 21412
rect 375374 21400 375380 21412
rect 270552 21372 375380 21400
rect 270552 21360 270558 21372
rect 375374 21360 375380 21372
rect 375432 21360 375438 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 29638 20652 29644 20664
rect 3476 20624 29644 20652
rect 3476 20612 3482 20624
rect 29638 20612 29644 20624
rect 29696 20612 29702 20664
rect 191098 20612 191104 20664
rect 191156 20652 191162 20664
rect 267734 20652 267740 20664
rect 191156 20624 267740 20652
rect 191156 20612 191162 20624
rect 267734 20612 267740 20624
rect 267792 20652 267798 20664
rect 268378 20652 268384 20664
rect 267792 20624 268384 20652
rect 267792 20612 267798 20624
rect 268378 20612 268384 20624
rect 268436 20612 268442 20664
rect 493318 20612 493324 20664
rect 493376 20652 493382 20664
rect 579982 20652 579988 20664
rect 493376 20624 579988 20652
rect 493376 20612 493382 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 84194 20000 84200 20052
rect 84252 20040 84258 20052
rect 233878 20040 233884 20052
rect 84252 20012 233884 20040
rect 84252 20000 84258 20012
rect 233878 20000 233884 20012
rect 233936 20000 233942 20052
rect 77294 19932 77300 19984
rect 77352 19972 77358 19984
rect 260190 19972 260196 19984
rect 77352 19944 260196 19972
rect 77352 19932 77358 19944
rect 260190 19932 260196 19944
rect 260248 19932 260254 19984
rect 273346 19932 273352 19984
rect 273404 19972 273410 19984
rect 376754 19972 376760 19984
rect 273404 19944 376760 19972
rect 273404 19932 273410 19944
rect 376754 19932 376760 19944
rect 376812 19932 376818 19984
rect 263594 19252 263600 19304
rect 263652 19292 263658 19304
rect 378134 19292 378140 19304
rect 263652 19264 378140 19292
rect 263652 19252 263658 19264
rect 378134 19252 378140 19264
rect 378192 19252 378198 19304
rect 195238 19184 195244 19236
rect 195296 19224 195302 19236
rect 273346 19224 273352 19236
rect 195296 19196 273352 19224
rect 195296 19184 195302 19196
rect 273346 19184 273352 19196
rect 273404 19184 273410 19236
rect 82814 18640 82820 18692
rect 82872 18680 82878 18692
rect 253290 18680 253296 18692
rect 82872 18652 253296 18680
rect 82872 18640 82878 18652
rect 253290 18640 253296 18652
rect 253348 18640 253354 18692
rect 70394 18572 70400 18624
rect 70452 18612 70458 18624
rect 250438 18612 250444 18624
rect 70452 18584 250444 18612
rect 70452 18572 70458 18584
rect 250438 18572 250444 18584
rect 250496 18572 250502 18624
rect 180058 17212 180064 17264
rect 180116 17252 180122 17264
rect 249794 17252 249800 17264
rect 180116 17224 249800 17252
rect 180116 17212 180122 17224
rect 249794 17212 249800 17224
rect 249852 17252 249858 17264
rect 382274 17252 382280 17264
rect 249852 17224 382280 17252
rect 249852 17212 249858 17224
rect 382274 17212 382280 17224
rect 382332 17212 382338 17264
rect 102134 15920 102140 15972
rect 102192 15960 102198 15972
rect 262950 15960 262956 15972
rect 102192 15932 262956 15960
rect 102192 15920 102198 15932
rect 262950 15920 262956 15932
rect 263008 15920 263014 15972
rect 21818 15852 21824 15904
rect 21876 15892 21882 15904
rect 238110 15892 238116 15904
rect 21876 15864 238116 15892
rect 21876 15852 21882 15864
rect 238110 15852 238116 15864
rect 238168 15852 238174 15904
rect 243538 15852 243544 15904
rect 243596 15892 243602 15904
rect 385034 15892 385040 15904
rect 243596 15864 385040 15892
rect 243596 15852 243602 15864
rect 385034 15852 385040 15864
rect 385092 15852 385098 15904
rect 87506 14492 87512 14544
rect 87564 14532 87570 14544
rect 257338 14532 257344 14544
rect 87564 14504 257344 14532
rect 87564 14492 87570 14504
rect 257338 14492 257344 14504
rect 257396 14492 257402 14544
rect 339494 14492 339500 14544
rect 339552 14532 339558 14544
rect 391934 14532 391940 14544
rect 339552 14504 391940 14532
rect 339552 14492 339558 14504
rect 391934 14492 391940 14504
rect 391992 14492 391998 14544
rect 164418 14424 164424 14476
rect 164476 14464 164482 14476
rect 350626 14464 350632 14476
rect 164476 14436 350632 14464
rect 164476 14424 164482 14436
rect 350626 14424 350632 14436
rect 350684 14424 350690 14476
rect 293218 13744 293224 13796
rect 293276 13784 293282 13796
rect 406378 13784 406384 13796
rect 293276 13756 406384 13784
rect 293276 13744 293282 13756
rect 406378 13744 406384 13756
rect 406436 13744 406442 13796
rect 188338 13200 188344 13252
rect 188396 13240 188402 13252
rect 261754 13240 261760 13252
rect 188396 13212 261760 13240
rect 188396 13200 188402 13212
rect 261754 13200 261760 13212
rect 261812 13240 261818 13252
rect 264422 13240 264428 13252
rect 261812 13212 264428 13240
rect 261812 13200 261818 13212
rect 264422 13200 264428 13212
rect 264480 13200 264486 13252
rect 80882 13132 80888 13184
rect 80940 13172 80946 13184
rect 239398 13172 239404 13184
rect 80940 13144 239404 13172
rect 80940 13132 80946 13144
rect 239398 13132 239404 13144
rect 239456 13132 239462 13184
rect 94682 13064 94688 13116
rect 94740 13104 94746 13116
rect 260098 13104 260104 13116
rect 94740 13076 260104 13104
rect 94740 13064 94746 13076
rect 260098 13064 260104 13076
rect 260156 13064 260162 13116
rect 283098 12384 283104 12436
rect 283156 12424 283162 12436
rect 283558 12424 283564 12436
rect 283156 12396 283564 12424
rect 283156 12384 283162 12396
rect 283558 12384 283564 12396
rect 283616 12424 283622 12436
rect 411254 12424 411260 12436
rect 283616 12396 411260 12424
rect 283616 12384 283622 12396
rect 411254 12384 411260 12396
rect 411312 12384 411318 12436
rect 20162 11772 20168 11824
rect 20220 11812 20226 11824
rect 232498 11812 232504 11824
rect 20220 11784 232504 11812
rect 20220 11772 20226 11784
rect 232498 11772 232504 11784
rect 232556 11772 232562 11824
rect 63402 11704 63408 11756
rect 63460 11744 63466 11756
rect 281902 11744 281908 11756
rect 63460 11716 281908 11744
rect 63460 11704 63466 11716
rect 281902 11704 281908 11716
rect 281960 11704 281966 11756
rect 33134 10956 33140 11008
rect 33192 10996 33198 11008
rect 34330 10996 34336 11008
rect 33192 10968 34336 10996
rect 33192 10956 33198 10968
rect 34330 10956 34336 10968
rect 34388 10996 34394 11008
rect 230474 10996 230480 11008
rect 34388 10968 230480 10996
rect 34388 10956 34394 10968
rect 230474 10956 230480 10968
rect 230532 10956 230538 11008
rect 258442 10888 258448 10940
rect 258500 10928 258506 10940
rect 259362 10928 259368 10940
rect 258500 10900 259368 10928
rect 258500 10888 258506 10900
rect 259362 10888 259368 10900
rect 259420 10888 259426 10940
rect 5442 10276 5448 10328
rect 5500 10316 5506 10328
rect 33134 10316 33140 10328
rect 5500 10288 33140 10316
rect 5500 10276 5506 10288
rect 33134 10276 33140 10288
rect 33192 10276 33198 10328
rect 78122 10276 78128 10328
rect 78180 10316 78186 10328
rect 255958 10316 255964 10328
rect 78180 10288 255964 10316
rect 78180 10276 78186 10288
rect 255958 10276 255964 10288
rect 256016 10276 256022 10328
rect 259362 10276 259368 10328
rect 259420 10316 259426 10328
rect 420914 10316 420920 10328
rect 259420 10288 420920 10316
rect 259420 10276 259426 10288
rect 420914 10276 420920 10288
rect 420972 10276 420978 10328
rect 186958 9596 186964 9648
rect 187016 9636 187022 9648
rect 278038 9636 278044 9648
rect 187016 9608 278044 9636
rect 187016 9596 187022 9608
rect 278038 9596 278044 9608
rect 278096 9636 278102 9648
rect 278314 9636 278320 9648
rect 278096 9608 278320 9636
rect 278096 9596 278102 9608
rect 278314 9596 278320 9608
rect 278372 9596 278378 9648
rect 102226 8984 102232 9036
rect 102284 9024 102290 9036
rect 261478 9024 261484 9036
rect 102284 8996 261484 9024
rect 102284 8984 102290 8996
rect 261478 8984 261484 8996
rect 261536 8984 261542 9036
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 229738 8956 229744 8968
rect 13596 8928 229744 8956
rect 13596 8916 13602 8928
rect 229738 8916 229744 8928
rect 229796 8916 229802 8968
rect 264974 8916 264980 8968
rect 265032 8956 265038 8968
rect 418154 8956 418160 8968
rect 265032 8928 418160 8956
rect 265032 8916 265038 8928
rect 418154 8916 418160 8928
rect 418212 8916 418218 8968
rect 251266 8168 251272 8220
rect 251324 8208 251330 8220
rect 252370 8208 252376 8220
rect 251324 8180 252376 8208
rect 251324 8168 251330 8180
rect 252370 8168 252376 8180
rect 252428 8168 252434 8220
rect 202138 7692 202144 7744
rect 202196 7732 202202 7744
rect 256694 7732 256700 7744
rect 202196 7704 256700 7732
rect 202196 7692 202202 7704
rect 256694 7692 256700 7704
rect 256752 7692 256758 7744
rect 70302 7624 70308 7676
rect 70360 7664 70366 7676
rect 246298 7664 246304 7676
rect 70360 7636 246304 7664
rect 70360 7624 70366 7636
rect 246298 7624 246304 7636
rect 246356 7624 246362 7676
rect 307018 7664 307024 7676
rect 296686 7636 307024 7664
rect 17034 7556 17040 7608
rect 17092 7596 17098 7608
rect 236730 7596 236736 7608
rect 17092 7568 236736 7596
rect 17092 7556 17098 7568
rect 236730 7556 236736 7568
rect 236788 7556 236794 7608
rect 252370 7556 252376 7608
rect 252428 7596 252434 7608
rect 296686 7596 296714 7636
rect 307018 7624 307024 7636
rect 307076 7624 307082 7676
rect 252428 7568 296714 7596
rect 252428 7556 252434 7568
rect 306742 7556 306748 7608
rect 306800 7596 306806 7608
rect 362954 7596 362960 7608
rect 306800 7568 362960 7596
rect 306800 7556 306806 7568
rect 362954 7556 362960 7568
rect 363012 7556 363018 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 15838 6848 15844 6860
rect 3476 6820 15844 6848
rect 3476 6808 3482 6820
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 281902 6808 281908 6860
rect 281960 6848 281966 6860
rect 371234 6848 371240 6860
rect 281960 6820 371240 6848
rect 281960 6808 281966 6820
rect 371234 6808 371240 6820
rect 371292 6808 371298 6860
rect 471238 6808 471244 6860
rect 471296 6848 471302 6860
rect 580166 6848 580172 6860
rect 471296 6820 580172 6848
rect 471296 6808 471302 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 38562 6264 38568 6316
rect 38620 6304 38626 6316
rect 136450 6304 136456 6316
rect 38620 6276 136456 6304
rect 38620 6264 38626 6276
rect 136450 6264 136456 6276
rect 136508 6264 136514 6316
rect 34422 6196 34428 6248
rect 34480 6236 34486 6248
rect 132954 6236 132960 6248
rect 34480 6208 132960 6236
rect 34480 6196 34486 6208
rect 132954 6196 132960 6208
rect 133012 6196 133018 6248
rect 15194 6128 15200 6180
rect 15252 6168 15258 6180
rect 265618 6168 265624 6180
rect 15252 6140 265624 6168
rect 15252 6128 15258 6140
rect 265618 6128 265624 6140
rect 265676 6128 265682 6180
rect 256694 5448 256700 5500
rect 256752 5488 256758 5500
rect 257062 5488 257068 5500
rect 256752 5460 257068 5488
rect 256752 5448 256758 5460
rect 257062 5448 257068 5460
rect 257120 5488 257126 5500
rect 380894 5488 380900 5500
rect 257120 5460 380900 5488
rect 257120 5448 257126 5460
rect 380894 5448 380900 5460
rect 380952 5448 380958 5500
rect 184198 4904 184204 4956
rect 184256 4944 184262 4956
rect 239122 4944 239128 4956
rect 184256 4916 239128 4944
rect 184256 4904 184262 4916
rect 239122 4904 239128 4916
rect 239180 4904 239186 4956
rect 91554 4836 91560 4888
rect 91612 4876 91618 4888
rect 249058 4876 249064 4888
rect 91612 4848 249064 4876
rect 91612 4836 91618 4848
rect 249058 4836 249064 4848
rect 249116 4836 249122 4888
rect 63218 4768 63224 4820
rect 63276 4808 63282 4820
rect 258718 4808 258724 4820
rect 63276 4780 258724 4808
rect 63276 4768 63282 4780
rect 258718 4768 258724 4780
rect 258776 4768 258782 4820
rect 349154 4224 349160 4276
rect 349212 4264 349218 4276
rect 353294 4264 353300 4276
rect 349212 4236 353300 4264
rect 349212 4224 349218 4236
rect 353294 4224 353300 4236
rect 353352 4224 353358 4276
rect 239122 4088 239128 4140
rect 239180 4128 239186 4140
rect 239306 4128 239312 4140
rect 239180 4100 239312 4128
rect 239180 4088 239186 4100
rect 239306 4088 239312 4100
rect 239364 4128 239370 4140
rect 269758 4128 269764 4140
rect 239364 4100 269764 4128
rect 239364 4088 239370 4100
rect 269758 4088 269764 4100
rect 269816 4088 269822 4140
rect 308398 4088 308404 4140
rect 308456 4128 308462 4140
rect 322198 4128 322204 4140
rect 308456 4100 322204 4128
rect 308456 4088 308462 4100
rect 322198 4088 322204 4100
rect 322256 4088 322262 4140
rect 216030 4020 216036 4072
rect 216088 4060 216094 4072
rect 242894 4060 242900 4072
rect 216088 4032 242900 4060
rect 216088 4020 216094 4032
rect 242894 4020 242900 4032
rect 242952 4060 242958 4072
rect 243538 4060 243544 4072
rect 242952 4032 243544 4060
rect 242952 4020 242958 4032
rect 243538 4020 243544 4032
rect 243596 4020 243602 4072
rect 125870 3612 125876 3664
rect 125928 3652 125934 3664
rect 173894 3652 173900 3664
rect 125928 3624 173900 3652
rect 125928 3612 125934 3624
rect 173894 3612 173900 3624
rect 173952 3612 173958 3664
rect 35802 3544 35808 3596
rect 35860 3584 35866 3596
rect 129366 3584 129372 3596
rect 35860 3556 129372 3584
rect 35860 3544 35866 3556
rect 129366 3544 129372 3556
rect 129424 3544 129430 3596
rect 244090 3544 244096 3596
rect 244148 3584 244154 3596
rect 245102 3584 245108 3596
rect 244148 3556 245108 3584
rect 244148 3544 244154 3556
rect 245102 3544 245108 3556
rect 245160 3544 245166 3596
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 276750 3584 276756 3596
rect 276072 3556 276756 3584
rect 276072 3544 276078 3556
rect 276750 3544 276756 3556
rect 276808 3544 276814 3596
rect 292574 3544 292580 3596
rect 292632 3584 292638 3596
rect 294046 3584 294052 3596
rect 292632 3556 294052 3584
rect 292632 3544 292638 3556
rect 294046 3544 294052 3556
rect 294104 3544 294110 3596
rect 316126 3544 316132 3596
rect 316184 3584 316190 3596
rect 317322 3584 317328 3596
rect 316184 3556 317328 3584
rect 316184 3544 316190 3556
rect 317322 3544 317328 3556
rect 317380 3544 317386 3596
rect 322106 3544 322112 3596
rect 322164 3584 322170 3596
rect 331214 3584 331220 3596
rect 322164 3556 331220 3584
rect 322164 3544 322170 3556
rect 331214 3544 331220 3556
rect 331272 3544 331278 3596
rect 346946 3544 346952 3596
rect 347004 3584 347010 3596
rect 356698 3584 356704 3596
rect 347004 3556 356704 3584
rect 347004 3544 347010 3556
rect 356698 3544 356704 3556
rect 356756 3544 356762 3596
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 28534 3516 28540 3528
rect 27672 3488 28540 3516
rect 27672 3476 27678 3488
rect 28534 3476 28540 3488
rect 28592 3476 28598 3528
rect 44174 3476 44180 3528
rect 44232 3516 44238 3528
rect 45094 3516 45100 3528
rect 44232 3488 45100 3516
rect 44232 3476 44238 3488
rect 45094 3476 45100 3488
rect 45152 3476 45158 3528
rect 52454 3476 52460 3528
rect 52512 3516 52518 3528
rect 53374 3516 53380 3528
rect 52512 3488 53380 3516
rect 52512 3476 52518 3488
rect 53374 3476 53380 3488
rect 53432 3476 53438 3528
rect 64322 3476 64328 3528
rect 64380 3516 64386 3528
rect 87598 3516 87604 3528
rect 64380 3488 87604 3516
rect 64380 3476 64386 3488
rect 87598 3476 87604 3488
rect 87656 3476 87662 3528
rect 102134 3476 102140 3528
rect 102192 3516 102198 3528
rect 103330 3516 103336 3528
rect 102192 3488 103336 3516
rect 102192 3476 102198 3488
rect 103330 3476 103336 3488
rect 103388 3476 103394 3528
rect 103422 3476 103428 3528
rect 103480 3516 103486 3528
rect 198090 3516 198096 3528
rect 103480 3488 198096 3516
rect 103480 3476 103486 3488
rect 198090 3476 198096 3488
rect 198148 3476 198154 3528
rect 266998 3476 267004 3528
rect 267056 3516 267062 3528
rect 274818 3516 274824 3528
rect 267056 3488 274824 3516
rect 267056 3476 267062 3488
rect 274818 3476 274824 3488
rect 274876 3516 274882 3528
rect 289078 3516 289084 3528
rect 274876 3488 289084 3516
rect 274876 3476 274882 3488
rect 289078 3476 289084 3488
rect 289136 3476 289142 3528
rect 290182 3476 290188 3528
rect 290240 3516 290246 3528
rect 295334 3516 295340 3528
rect 290240 3488 295340 3516
rect 290240 3476 290246 3488
rect 295334 3476 295340 3488
rect 295392 3476 295398 3528
rect 304350 3476 304356 3528
rect 304408 3516 304414 3528
rect 304994 3516 305000 3528
rect 304408 3488 305000 3516
rect 304408 3476 304414 3488
rect 304994 3476 305000 3488
rect 305052 3476 305058 3528
rect 309042 3476 309048 3528
rect 309100 3516 309106 3528
rect 309778 3516 309784 3528
rect 309100 3488 309784 3516
rect 309100 3476 309106 3488
rect 309778 3476 309784 3488
rect 309836 3476 309842 3528
rect 324314 3476 324320 3528
rect 324372 3516 324378 3528
rect 325602 3516 325608 3528
rect 324372 3488 325608 3516
rect 324372 3476 324378 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 332594 3476 332600 3528
rect 332652 3516 332658 3528
rect 333882 3516 333888 3528
rect 332652 3488 333888 3516
rect 332652 3476 332658 3488
rect 333882 3476 333888 3488
rect 333940 3476 333946 3528
rect 340138 3516 340144 3528
rect 334084 3488 340144 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 15194 3448 15200 3460
rect 6512 3420 15200 3448
rect 6512 3408 6518 3420
rect 15194 3408 15200 3420
rect 15252 3408 15258 3460
rect 35986 3408 35992 3460
rect 36044 3448 36050 3460
rect 214558 3448 214564 3460
rect 36044 3420 214564 3448
rect 36044 3408 36050 3420
rect 214558 3408 214564 3420
rect 214616 3408 214622 3460
rect 216122 3408 216128 3460
rect 216180 3448 216186 3460
rect 285398 3448 285404 3460
rect 216180 3420 285404 3448
rect 216180 3408 216186 3420
rect 285398 3408 285404 3420
rect 285456 3448 285462 3460
rect 287698 3448 287704 3460
rect 285456 3420 287704 3448
rect 285456 3408 285462 3420
rect 287698 3408 287704 3420
rect 287756 3408 287762 3460
rect 332686 3408 332692 3460
rect 332744 3448 332750 3460
rect 334084 3448 334112 3488
rect 340138 3476 340144 3488
rect 340196 3476 340202 3528
rect 340874 3476 340880 3528
rect 340932 3516 340938 3528
rect 342162 3516 342168 3528
rect 340932 3488 342168 3516
rect 340932 3476 340938 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 350442 3476 350448 3528
rect 350500 3516 350506 3528
rect 351914 3516 351920 3528
rect 350500 3488 351920 3516
rect 350500 3476 350506 3488
rect 351914 3476 351920 3488
rect 351972 3476 351978 3528
rect 349154 3448 349160 3460
rect 332744 3420 334112 3448
rect 335326 3420 349160 3448
rect 332744 3408 332750 3420
rect 99834 3340 99840 3392
rect 99892 3380 99898 3392
rect 103422 3380 103428 3392
rect 99892 3352 103428 3380
rect 99892 3340 99898 3352
rect 103422 3340 103428 3352
rect 103480 3340 103486 3392
rect 331582 3340 331588 3392
rect 331640 3380 331646 3392
rect 335326 3380 335354 3420
rect 349154 3408 349160 3420
rect 349212 3408 349218 3460
rect 351638 3408 351644 3460
rect 351696 3448 351702 3460
rect 388438 3448 388444 3460
rect 351696 3420 388444 3448
rect 351696 3408 351702 3420
rect 388438 3408 388444 3420
rect 388496 3408 388502 3460
rect 331640 3352 335354 3380
rect 331640 3340 331646 3352
rect 267734 3272 267740 3324
rect 267792 3312 267798 3324
rect 273346 3312 273352 3324
rect 267792 3284 273352 3312
rect 267792 3272 267798 3284
rect 273346 3272 273352 3284
rect 273404 3272 273410 3324
rect 1670 3204 1676 3256
rect 1728 3244 1734 3256
rect 5442 3244 5448 3256
rect 1728 3216 5448 3244
rect 1728 3204 1734 3216
rect 5442 3204 5448 3216
rect 5500 3204 5506 3256
rect 299658 3136 299664 3188
rect 299716 3176 299722 3188
rect 302234 3176 302240 3188
rect 299716 3148 302240 3176
rect 299716 3136 299722 3148
rect 302234 3136 302240 3148
rect 302292 3136 302298 3188
rect 233970 3000 233976 3052
rect 234028 3040 234034 3052
rect 235810 3040 235816 3052
rect 234028 3012 235816 3040
rect 234028 3000 234034 3012
rect 235810 3000 235816 3012
rect 235868 3000 235874 3052
rect 279510 2932 279516 2984
rect 279568 2972 279574 2984
rect 280246 2972 280252 2984
rect 279568 2944 280252 2972
rect 279568 2932 279574 2944
rect 280246 2932 280252 2944
rect 280304 2932 280310 2984
rect 109310 2048 109316 2100
rect 109368 2088 109374 2100
rect 242158 2088 242164 2100
rect 109368 2060 242164 2088
rect 109368 2048 109374 2060
rect 242158 2048 242164 2060
rect 242216 2048 242222 2100
<< via1 >>
rect 201500 703264 201552 703316
rect 202788 703264 202840 703316
rect 77944 703196 77996 703248
rect 267648 703196 267700 703248
rect 95148 703128 95200 703180
rect 332508 703128 332560 703180
rect 110328 703060 110380 703112
rect 348792 703060 348844 703112
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 76564 702992 76616 703044
rect 364984 702992 365036 703044
rect 104808 702924 104860 702976
rect 413652 702924 413704 702976
rect 111708 702856 111760 702908
rect 462320 702856 462372 702908
rect 75184 702788 75236 702840
rect 381544 702788 381596 702840
rect 386420 702788 386472 702840
rect 424968 702788 425020 702840
rect 429844 702788 429896 702840
rect 117228 702720 117280 702772
rect 478512 702720 478564 702772
rect 113088 702652 113140 702704
rect 494796 702652 494848 702704
rect 79324 702584 79376 702636
rect 527180 702584 527232 702636
rect 108948 702516 109000 702568
rect 465724 702516 465776 702568
rect 550548 702516 550600 702568
rect 559656 702516 559708 702568
rect 68928 702448 68980 702500
rect 543464 702448 543516 702500
rect 69664 700340 69716 700392
rect 154120 700340 154172 700392
rect 155224 700340 155276 700392
rect 218980 700340 219032 700392
rect 62028 700272 62080 700324
rect 235172 700272 235224 700324
rect 238024 700272 238076 700324
rect 283840 700272 283892 700324
rect 386420 700272 386472 700324
rect 424968 700272 425020 700324
rect 465724 700272 465776 700324
rect 550548 700272 550600 700324
rect 24308 698912 24360 698964
rect 106280 698912 106332 698964
rect 159364 683136 159416 683188
rect 579620 683136 579672 683188
rect 3516 670692 3568 670744
rect 54484 670692 54536 670744
rect 90364 670692 90416 670744
rect 579620 670692 579672 670744
rect 579988 670692 580040 670744
rect 3516 656888 3568 656940
rect 11704 656888 11756 656940
rect 457444 643696 457496 643748
rect 579620 643696 579672 643748
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 130384 630640 130436 630692
rect 580172 630640 580224 630692
rect 3516 618264 3568 618316
rect 86960 618264 87012 618316
rect 3516 605820 3568 605872
rect 35164 605820 35216 605872
rect 6920 598204 6972 598256
rect 52368 598204 52420 598256
rect 52368 597524 52420 597576
rect 85580 597524 85632 597576
rect 68744 596776 68796 596828
rect 136640 596776 136692 596828
rect 3424 595416 3476 595468
rect 42800 595416 42852 595468
rect 42800 594804 42852 594856
rect 44088 594804 44140 594856
rect 71872 594804 71924 594856
rect 69020 594056 69072 594108
rect 580264 594056 580316 594108
rect 81808 591268 81860 591320
rect 90364 591268 90416 591320
rect 40040 590656 40092 590708
rect 48228 590656 48280 590708
rect 74632 590656 74684 590708
rect 556804 590656 556856 590708
rect 580172 590656 580224 590708
rect 91468 589296 91520 589348
rect 124220 589296 124272 589348
rect 86960 588956 87012 589008
rect 88248 588956 88300 589008
rect 11704 588548 11756 588600
rect 87696 588548 87748 588600
rect 88340 588548 88392 588600
rect 116124 588548 116176 588600
rect 56416 587868 56468 587920
rect 86960 587868 87012 587920
rect 121460 587120 121512 587172
rect 155224 587120 155276 587172
rect 59176 586644 59228 586696
rect 83188 586644 83240 586696
rect 94872 586644 94924 586696
rect 125600 586644 125652 586696
rect 39764 586576 39816 586628
rect 79324 586576 79376 586628
rect 87696 586576 87748 586628
rect 120172 586576 120224 586628
rect 42616 586508 42668 586560
rect 83004 586508 83056 586560
rect 85304 586508 85356 586560
rect 118700 586508 118752 586560
rect 68836 585760 68888 585812
rect 238024 585760 238076 585812
rect 103520 585420 103572 585472
rect 104808 585420 104860 585472
rect 122840 585420 122892 585472
rect 102416 585352 102468 585404
rect 121460 585352 121512 585404
rect 52276 585284 52328 585336
rect 76564 585284 76616 585336
rect 95148 585284 95200 585336
rect 114560 585284 114612 585336
rect 53472 585216 53524 585268
rect 78036 585216 78088 585268
rect 94136 585216 94188 585268
rect 116216 585216 116268 585268
rect 41144 585148 41196 585200
rect 80612 585148 80664 585200
rect 89628 585148 89680 585200
rect 121552 585148 121604 585200
rect 88248 585080 88300 585132
rect 95424 585080 95476 585132
rect 98736 585012 98788 585064
rect 102416 585012 102468 585064
rect 57796 583992 57848 584044
rect 73344 584060 73396 584112
rect 102600 584060 102652 584112
rect 106648 584060 106700 584112
rect 53748 583924 53800 583976
rect 70400 583992 70452 584044
rect 77852 583992 77904 584044
rect 79232 583992 79284 584044
rect 104624 583992 104676 584044
rect 136640 583992 136692 584044
rect 68468 583924 68520 583976
rect 69664 583924 69716 583976
rect 101312 583924 101364 583976
rect 113364 583924 113416 583976
rect 60648 583856 60700 583908
rect 81900 583856 81952 583908
rect 96528 583856 96580 583908
rect 110512 583856 110564 583908
rect 45376 583788 45428 583840
rect 78680 583788 78732 583840
rect 99288 583788 99340 583840
rect 128360 583788 128412 583840
rect 41328 583720 41380 583772
rect 77852 583720 77904 583772
rect 105544 583720 105596 583772
rect 114652 583720 114704 583772
rect 59084 582972 59136 583024
rect 71780 582972 71832 583024
rect 97448 582700 97500 582752
rect 120264 582700 120316 582752
rect 92848 582632 92900 582684
rect 117412 582632 117464 582684
rect 43996 582564 44048 582616
rect 76748 582564 76800 582616
rect 90272 582564 90324 582616
rect 118792 582564 118844 582616
rect 46664 582496 46716 582548
rect 84476 582496 84528 582548
rect 91008 582496 91060 582548
rect 122932 582496 122984 582548
rect 3424 582428 3476 582480
rect 107660 582428 107712 582480
rect 69204 582360 69256 582412
rect 580172 582360 580224 582412
rect 66168 581816 66220 581868
rect 70952 581816 71004 581868
rect 37096 581272 37148 581324
rect 75460 581748 75512 581800
rect 104440 581748 104492 581800
rect 108672 581748 108724 581800
rect 68744 581680 68796 581732
rect 72240 581680 72292 581732
rect 50344 581204 50396 581256
rect 67640 581204 67692 581256
rect 57888 581136 57940 581188
rect 84016 581680 84068 581732
rect 97908 581680 97960 581732
rect 35808 581068 35860 581120
rect 68744 581068 68796 581120
rect 103888 581680 103940 581732
rect 113272 581136 113324 581188
rect 108672 581068 108724 581120
rect 128452 581068 128504 581120
rect 128636 581000 128688 581052
rect 106648 580932 106700 580984
rect 114836 580932 114888 580984
rect 39948 580252 40000 580304
rect 67824 580252 67876 580304
rect 108948 579708 109000 579760
rect 126980 579708 127032 579760
rect 3332 579640 3384 579692
rect 53104 579640 53156 579692
rect 69112 579028 69164 579080
rect 69756 579028 69808 579080
rect 59268 578280 59320 578332
rect 67640 578280 67692 578332
rect 108396 578280 108448 578332
rect 111892 578280 111944 578332
rect 108948 578212 109000 578264
rect 131120 578212 131172 578264
rect 108856 577464 108908 577516
rect 115940 577464 115992 577516
rect 66076 577396 66128 577448
rect 68192 577396 68244 577448
rect 108948 576852 109000 576904
rect 138020 576852 138072 576904
rect 108948 576104 109000 576156
rect 123116 576104 123168 576156
rect 38568 575492 38620 575544
rect 67640 575492 67692 575544
rect 108488 575492 108540 575544
rect 117320 575492 117372 575544
rect 123116 575492 123168 575544
rect 429844 575492 429896 575544
rect 52184 574064 52236 574116
rect 67640 574064 67692 574116
rect 126888 573996 126940 574048
rect 159364 573996 159416 574048
rect 108948 573316 109000 573368
rect 126152 573316 126204 573368
rect 126888 573316 126940 573368
rect 105636 572840 105688 572892
rect 110604 572840 110656 572892
rect 65984 572772 66036 572824
rect 67732 572772 67784 572824
rect 61936 572704 61988 572756
rect 67640 572704 67692 572756
rect 107660 572704 107712 572756
rect 110420 572704 110472 572756
rect 55036 572024 55088 572076
rect 67824 572024 67876 572076
rect 49516 571956 49568 572008
rect 67916 571956 67968 572008
rect 108948 571344 109000 571396
rect 130016 571344 130068 571396
rect 66168 571276 66220 571328
rect 68284 571276 68336 571328
rect 108856 569984 108908 570036
rect 136732 569984 136784 570036
rect 63224 569916 63276 569968
rect 67640 569916 67692 569968
rect 108948 569916 109000 569968
rect 139400 569916 139452 569968
rect 66168 568624 66220 568676
rect 67732 568624 67784 568676
rect 34244 568556 34296 568608
rect 67640 568556 67692 568608
rect 108948 568556 109000 568608
rect 124864 568556 124916 568608
rect 108948 567536 109000 567588
rect 113824 567536 113876 567588
rect 64604 567264 64656 567316
rect 67640 567264 67692 567316
rect 60464 567196 60516 567248
rect 67732 567196 67784 567248
rect 108948 567196 109000 567248
rect 117964 567196 118016 567248
rect 106924 566448 106976 566500
rect 121644 566448 121696 566500
rect 108396 565904 108448 565956
rect 111984 565904 112036 565956
rect 3240 565836 3292 565888
rect 25504 565836 25556 565888
rect 64696 565836 64748 565888
rect 67640 565836 67692 565888
rect 108948 565836 109000 565888
rect 140872 565836 140924 565888
rect 48044 564476 48096 564528
rect 67640 564476 67692 564528
rect 117228 564476 117280 564528
rect 132592 564476 132644 564528
rect 108948 564408 109000 564460
rect 143448 564408 143500 564460
rect 204904 564408 204956 564460
rect 108396 564340 108448 564392
rect 117228 564340 117280 564392
rect 374644 563660 374696 563712
rect 429844 563660 429896 563712
rect 580172 563660 580224 563712
rect 63132 563116 63184 563168
rect 67640 563116 67692 563168
rect 56508 563048 56560 563100
rect 67732 563048 67784 563100
rect 60740 562300 60792 562352
rect 62028 562300 62080 562352
rect 67640 562300 67692 562352
rect 61752 561688 61804 561740
rect 67640 561688 67692 561740
rect 108948 561688 109000 561740
rect 135444 561688 135496 561740
rect 53564 560940 53616 560992
rect 60740 560940 60792 560992
rect 58992 560328 59044 560380
rect 67732 560328 67784 560380
rect 108212 560328 108264 560380
rect 131396 560328 131448 560380
rect 55128 560260 55180 560312
rect 67640 560260 67692 560312
rect 108948 560260 109000 560312
rect 133972 560260 134024 560312
rect 135168 559512 135220 559564
rect 201500 559512 201552 559564
rect 108948 558968 109000 559020
rect 132776 558968 132828 559020
rect 41236 558900 41288 558952
rect 67640 558900 67692 558952
rect 108856 558900 108908 558952
rect 133880 558900 133932 558952
rect 135168 558900 135220 558952
rect 64788 558220 64840 558272
rect 68836 558220 68888 558272
rect 59176 558152 59228 558204
rect 69756 558152 69808 558204
rect 108948 557540 109000 557592
rect 116032 557540 116084 557592
rect 48136 556248 48188 556300
rect 67640 556248 67692 556300
rect 42708 556180 42760 556232
rect 67732 556180 67784 556232
rect 108948 556180 109000 556232
rect 136824 556180 136876 556232
rect 108856 556112 108908 556164
rect 110604 556112 110656 556164
rect 110604 555432 110656 555484
rect 125968 555432 126020 555484
rect 57612 554820 57664 554872
rect 67640 554820 67692 554872
rect 36544 554752 36596 554804
rect 67732 554752 67784 554804
rect 140964 554004 141016 554056
rect 556804 554004 556856 554056
rect 58624 553392 58676 553444
rect 67640 553392 67692 553444
rect 108948 553392 109000 553444
rect 140964 553392 141016 553444
rect 54944 552032 54996 552084
rect 67640 552032 67692 552084
rect 35716 550604 35768 550656
rect 67640 550604 67692 550656
rect 108948 550604 109000 550656
rect 120080 550604 120132 550656
rect 63316 549312 63368 549364
rect 67640 549312 67692 549364
rect 108856 549312 108908 549364
rect 134248 549312 134300 549364
rect 61844 549244 61896 549296
rect 67732 549244 67784 549296
rect 108948 549244 109000 549296
rect 142160 549244 142212 549296
rect 34336 547884 34388 547936
rect 67640 547884 67692 547936
rect 108948 547884 109000 547936
rect 139584 547884 139636 547936
rect 60556 546456 60608 546508
rect 67640 546456 67692 546508
rect 108948 546456 109000 546508
rect 135352 546456 135404 546508
rect 108948 545708 109000 545760
rect 113088 545708 113140 545760
rect 119344 545708 119396 545760
rect 108948 545096 109000 545148
rect 138204 545096 138256 545148
rect 25504 544348 25556 544400
rect 67732 544348 67784 544400
rect 60280 542444 60332 542496
rect 67640 542444 67692 542496
rect 49608 542376 49660 542428
rect 68008 542376 68060 542428
rect 108948 542376 109000 542428
rect 134156 542376 134208 542428
rect 60648 541628 60700 541680
rect 69664 541628 69716 541680
rect 128544 541628 128596 541680
rect 299480 541628 299532 541680
rect 64144 541016 64196 541068
rect 67732 541016 67784 541068
rect 63408 540948 63460 541000
rect 67640 540948 67692 541000
rect 109684 540948 109736 541000
rect 128544 540948 128596 541000
rect 108948 539656 109000 539708
rect 110328 539656 110380 539708
rect 114744 539656 114796 539708
rect 62028 539588 62080 539640
rect 67640 539588 67692 539640
rect 107844 539588 107896 539640
rect 127072 539588 127124 539640
rect 35164 539520 35216 539572
rect 105820 539520 105872 539572
rect 54484 538908 54536 538960
rect 73160 538908 73212 538960
rect 95056 538908 95108 538960
rect 109132 538908 109184 538960
rect 4804 538840 4856 538892
rect 82268 538840 82320 538892
rect 95148 538840 95200 538892
rect 116216 538840 116268 538892
rect 122104 538840 122156 538892
rect 580356 538840 580408 538892
rect 53104 538160 53156 538212
rect 98368 538160 98420 538212
rect 103520 538160 103572 538212
rect 109684 538160 109736 538212
rect 88064 538092 88116 538144
rect 122104 538228 122156 538280
rect 204904 538160 204956 538212
rect 580172 538160 580224 538212
rect 73160 538024 73212 538076
rect 91284 538024 91336 538076
rect 82268 537956 82320 538008
rect 99012 537956 99064 538008
rect 57888 537752 57940 537804
rect 79324 537752 79376 537804
rect 94504 537684 94556 537736
rect 104716 537684 104768 537736
rect 57888 537616 57940 537668
rect 81624 537616 81676 537668
rect 95792 537616 95844 537668
rect 123024 537616 123076 537668
rect 43812 537548 43864 537600
rect 72608 537548 72660 537600
rect 102232 537548 102284 537600
rect 129832 537548 129884 537600
rect 50988 537480 51040 537532
rect 82912 537480 82964 537532
rect 102876 537480 102928 537532
rect 132684 537480 132736 537532
rect 73160 536868 73212 536920
rect 73804 536868 73856 536920
rect 84844 536868 84896 536920
rect 90364 536868 90416 536920
rect 70124 536800 70176 536852
rect 75920 536800 75972 536852
rect 82268 536800 82320 536852
rect 82728 536800 82780 536852
rect 84108 536800 84160 536852
rect 85488 536800 85540 536852
rect 102048 536800 102100 536852
rect 105544 536800 105596 536852
rect 59084 536732 59136 536784
rect 73896 536732 73948 536784
rect 57612 536188 57664 536240
rect 65892 536188 65944 536240
rect 45468 536120 45520 536172
rect 59084 536120 59136 536172
rect 104716 536120 104768 536172
rect 109132 536120 109184 536172
rect 116124 536120 116176 536172
rect 37188 536052 37240 536104
rect 71320 536052 71372 536104
rect 97908 536052 97960 536104
rect 114836 536052 114888 536104
rect 56324 535440 56376 535492
rect 57612 535440 57664 535492
rect 65892 535372 65944 535424
rect 169760 535372 169812 535424
rect 72424 534896 72476 534948
rect 77760 534896 77812 534948
rect 99288 534896 99340 534948
rect 113272 534896 113324 534948
rect 53656 534828 53708 534880
rect 75184 534828 75236 534880
rect 98644 534828 98696 534880
rect 117412 534828 117464 534880
rect 46848 534760 46900 534812
rect 78404 534760 78456 534812
rect 93860 534760 93912 534812
rect 125784 534760 125836 534812
rect 39856 534692 39908 534744
rect 73252 534692 73304 534744
rect 89996 534692 90048 534744
rect 124404 534692 124456 534744
rect 69296 533332 69348 533384
rect 69756 533332 69808 533384
rect 49332 532108 49384 532160
rect 76472 532108 76524 532160
rect 52000 532040 52052 532092
rect 83556 532040 83608 532092
rect 89352 532040 89404 532092
rect 113272 532040 113324 532092
rect 47952 531972 48004 532024
rect 79048 531972 79100 532024
rect 93768 531972 93820 532024
rect 124220 531972 124272 532024
rect 54852 529320 54904 529372
rect 77116 529320 77168 529372
rect 41052 529252 41104 529304
rect 70400 529252 70452 529304
rect 42524 529184 42576 529236
rect 74540 529184 74592 529236
rect 3148 528504 3200 528556
rect 107016 528572 107068 528624
rect 124956 528572 125008 528624
rect 39672 526396 39724 526448
rect 71964 526396 72016 526448
rect 34152 525784 34204 525836
rect 64144 525784 64196 525836
rect 579804 525716 579856 525768
rect 3424 514768 3476 514820
rect 7564 514768 7616 514820
rect 59268 511980 59320 512032
rect 67456 511980 67508 512032
rect 67456 511232 67508 511284
rect 405740 511232 405792 511284
rect 405740 510620 405792 510672
rect 580172 510620 580224 510672
rect 93216 500420 93268 500472
rect 116124 500420 116176 500472
rect 84108 500352 84160 500404
rect 110604 500352 110656 500404
rect 91100 500284 91152 500336
rect 128636 500284 128688 500336
rect 7564 500216 7616 500268
rect 91744 500216 91796 500268
rect 91928 500216 91980 500268
rect 124312 500216 124364 500268
rect 135260 500216 135312 500268
rect 84200 498788 84252 498840
rect 118884 498788 118936 498840
rect 81440 498176 81492 498228
rect 114928 498176 114980 498228
rect 87420 497564 87472 497616
rect 112076 497564 112128 497616
rect 90640 497496 90692 497548
rect 120448 497496 120500 497548
rect 69664 497428 69716 497480
rect 75828 497428 75880 497480
rect 81440 497428 81492 497480
rect 83832 497428 83884 497480
rect 118792 497428 118844 497480
rect 131212 497428 131264 497480
rect 88248 496136 88300 496188
rect 121644 496136 121696 496188
rect 129004 496136 129056 496188
rect 50712 496068 50764 496120
rect 80980 496068 81032 496120
rect 93216 496068 93268 496120
rect 128360 496068 128412 496120
rect 136916 496068 136968 496120
rect 42616 495592 42668 495644
rect 76104 495592 76156 495644
rect 39764 495524 39816 495576
rect 73252 495524 73304 495576
rect 41144 495456 41196 495508
rect 74540 495456 74592 495508
rect 3424 495388 3476 495440
rect 83832 495388 83884 495440
rect 96436 494980 96488 495032
rect 113180 494980 113232 495032
rect 98736 494912 98788 494964
rect 121644 494912 121696 494964
rect 82268 494844 82320 494896
rect 111800 494844 111852 494896
rect 82728 494776 82780 494828
rect 120356 494776 120408 494828
rect 80980 494708 81032 494760
rect 120172 494708 120224 494760
rect 128360 494708 128412 494760
rect 85488 494164 85540 494216
rect 89628 494164 89680 494216
rect 79324 494028 79376 494080
rect 79968 494028 80020 494080
rect 123116 494028 123168 494080
rect 97724 493960 97776 494012
rect 102140 493960 102192 494012
rect 70860 493688 70912 493740
rect 72424 493688 72476 493740
rect 95240 493484 95292 493536
rect 81624 493416 81676 493468
rect 88248 493416 88300 493468
rect 90272 493416 90324 493468
rect 110512 493416 110564 493468
rect 113364 493416 113416 493468
rect 132500 493416 132552 493468
rect 57704 493348 57756 493400
rect 74816 493348 74868 493400
rect 82912 493348 82964 493400
rect 121552 493348 121604 493400
rect 127164 493348 127216 493400
rect 43720 493280 43772 493332
rect 53472 493280 53524 493332
rect 71780 493280 71832 493332
rect 79692 493280 79744 493332
rect 118700 493280 118752 493332
rect 125876 493280 125928 493332
rect 51908 492804 51960 492856
rect 52276 492804 52328 492856
rect 70032 492804 70084 492856
rect 58900 492736 58952 492788
rect 90272 492736 90324 492788
rect 56416 492668 56468 492720
rect 89720 492668 89772 492720
rect 77760 492600 77812 492652
rect 79968 492600 80020 492652
rect 91284 492600 91336 492652
rect 91744 492600 91796 492652
rect 120264 492600 120316 492652
rect 120264 492328 120316 492380
rect 121552 492328 121604 492380
rect 97724 492260 97776 492312
rect 99288 492260 99340 492312
rect 96436 492056 96488 492108
rect 97908 492056 97960 492108
rect 38476 491988 38528 492040
rect 43996 491988 44048 492040
rect 70400 491988 70452 492040
rect 43904 491920 43956 491972
rect 45376 491920 45428 491972
rect 72240 491920 72292 491972
rect 99288 491988 99340 492040
rect 111064 491988 111116 492040
rect 109776 491920 109828 491972
rect 88708 491580 88760 491632
rect 100668 491580 100720 491632
rect 84844 491512 84896 491564
rect 122932 491512 122984 491564
rect 99012 491444 99064 491496
rect 110512 491444 110564 491496
rect 41328 491376 41380 491428
rect 52368 491376 52420 491428
rect 80060 491376 80112 491428
rect 86776 491376 86828 491428
rect 70952 491308 71004 491360
rect 86132 491308 86184 491360
rect 93768 491308 93820 491360
rect 58624 491240 58676 491292
rect 63500 491240 63552 491292
rect 99656 491376 99708 491428
rect 114652 491376 114704 491428
rect 115480 491376 115532 491428
rect 98644 491240 98696 491292
rect 101404 491240 101456 491292
rect 110512 491240 110564 491292
rect 111708 491240 111760 491292
rect 136640 491240 136692 491292
rect 100668 491172 100720 491224
rect 114560 491172 114612 491224
rect 115480 491172 115532 491224
rect 118792 491172 118844 491224
rect 59084 490764 59136 490816
rect 73804 490764 73856 490816
rect 93860 490764 93912 490816
rect 100024 490764 100076 490816
rect 56232 490696 56284 490748
rect 79600 490696 79652 490748
rect 45376 490628 45428 490680
rect 46664 490628 46716 490680
rect 78036 490628 78088 490680
rect 92848 490628 92900 490680
rect 106280 490628 106332 490680
rect 35532 490560 35584 490612
rect 37096 490560 37148 490612
rect 69756 490560 69808 490612
rect 94136 490560 94188 490612
rect 94964 490560 95016 490612
rect 109684 490560 109736 490612
rect 114836 490560 114888 490612
rect 125600 490560 125652 490612
rect 75920 490152 75972 490204
rect 77070 490152 77122 490204
rect 88248 489948 88300 490000
rect 114836 489948 114888 490000
rect 77300 489880 77352 489932
rect 111800 489880 111852 489932
rect 69848 489812 69900 489864
rect 70860 489812 70912 489864
rect 98736 489812 98788 489864
rect 99288 489812 99340 489864
rect 106280 489812 106332 489864
rect 107384 489812 107436 489864
rect 121460 489812 121512 489864
rect 115848 489132 115900 489184
rect 126980 489132 127032 489184
rect 103428 488588 103480 488640
rect 115848 488588 115900 488640
rect 99288 488520 99340 488572
rect 103336 488452 103388 488504
rect 111892 488452 111944 488504
rect 122932 488520 122984 488572
rect 131488 488520 131540 488572
rect 114376 488452 114428 488504
rect 128452 488452 128504 488504
rect 102876 488384 102928 488436
rect 109040 488384 109092 488436
rect 111892 487908 111944 487960
rect 116216 487908 116268 487960
rect 48228 487840 48280 487892
rect 57244 487840 57296 487892
rect 109040 487840 109092 487892
rect 122932 487840 122984 487892
rect 50804 487772 50856 487824
rect 67640 487772 67692 487824
rect 106280 487772 106332 487824
rect 138020 487772 138072 487824
rect 147680 487772 147732 487824
rect 56600 487160 56652 487212
rect 57244 487160 57296 487212
rect 67640 487160 67692 487212
rect 35808 487092 35860 487144
rect 68100 487092 68152 487144
rect 103336 487092 103388 487144
rect 131120 487092 131172 487144
rect 131304 487092 131356 487144
rect 131304 486412 131356 486464
rect 142344 486412 142396 486464
rect 103428 486004 103480 486056
rect 106280 486004 106332 486056
rect 57796 485732 57848 485784
rect 65524 485800 65576 485852
rect 67640 485800 67692 485852
rect 102232 485732 102284 485784
rect 115940 485732 115992 485784
rect 117228 485732 117280 485784
rect 131304 485052 131356 485104
rect 131488 485052 131540 485104
rect 64512 484508 64564 484560
rect 68376 484508 68428 484560
rect 44088 484304 44140 484356
rect 53288 484372 53340 484424
rect 67640 484372 67692 484424
rect 102232 484372 102284 484424
rect 113088 484304 113140 484356
rect 117320 484304 117372 484356
rect 102232 483624 102284 483676
rect 123208 483624 123260 483676
rect 37096 483012 37148 483064
rect 50344 483012 50396 483064
rect 104716 483012 104768 483064
rect 125692 483012 125744 483064
rect 67640 482944 67692 482996
rect 102324 482944 102376 482996
rect 106372 482944 106424 482996
rect 107568 482944 107620 482996
rect 115848 482944 115900 482996
rect 117688 482944 117740 482996
rect 102232 482604 102284 482656
rect 104716 482604 104768 482656
rect 107568 481720 107620 481772
rect 115296 481720 115348 481772
rect 102232 481584 102284 481636
rect 106188 481652 106240 481704
rect 150624 481652 150676 481704
rect 110420 481584 110472 481636
rect 111156 481584 111208 481636
rect 102324 481516 102376 481568
rect 106188 481448 106240 481500
rect 39948 480904 40000 480956
rect 67640 480904 67692 480956
rect 101956 480904 102008 480956
rect 130016 480904 130068 480956
rect 147864 480904 147916 480956
rect 59268 480224 59320 480276
rect 67548 480224 67600 480276
rect 111156 480224 111208 480276
rect 113364 480224 113416 480276
rect 102232 480156 102284 480208
rect 104900 480156 104952 480208
rect 66076 479680 66128 479732
rect 68376 479680 68428 479732
rect 124864 478864 124916 478916
rect 137008 478864 137060 478916
rect 105544 477572 105596 477624
rect 107936 477572 107988 477624
rect 102876 477504 102928 477556
rect 111892 477504 111944 477556
rect 102324 477436 102376 477488
rect 113824 477504 113876 477556
rect 118700 477504 118752 477556
rect 102232 477368 102284 477420
rect 124864 477368 124916 477420
rect 111892 477300 111944 477352
rect 113088 477300 113140 477352
rect 136732 477300 136784 477352
rect 34428 476076 34480 476128
rect 67640 476076 67692 476128
rect 117964 476076 118016 476128
rect 128452 476076 128504 476128
rect 102416 476008 102468 476060
rect 103336 476008 103388 476060
rect 139400 476008 139452 476060
rect 102232 475940 102284 475992
rect 117964 475940 118016 475992
rect 102324 475872 102376 475924
rect 111892 475872 111944 475924
rect 51080 475396 51132 475448
rect 52184 475396 52236 475448
rect 67640 475396 67692 475448
rect 35624 475328 35676 475380
rect 65984 475328 66036 475380
rect 67732 475328 67784 475380
rect 111892 475328 111944 475380
rect 121460 475328 121512 475380
rect 3424 474716 3476 474768
rect 25504 474716 25556 474768
rect 60372 474648 60424 474700
rect 61936 474648 61988 474700
rect 67640 474648 67692 474700
rect 102232 474648 102284 474700
rect 140872 474648 140924 474700
rect 141240 474648 141292 474700
rect 44088 473968 44140 474020
rect 51080 473968 51132 474020
rect 113088 473968 113140 474020
rect 117320 473968 117372 474020
rect 141240 473968 141292 474020
rect 144920 473968 144972 474020
rect 49516 473288 49568 473340
rect 65616 473356 65668 473408
rect 67640 473356 67692 473408
rect 100300 473288 100352 473340
rect 100760 473288 100812 473340
rect 102324 472676 102376 472728
rect 103428 472676 103480 472728
rect 109040 472676 109092 472728
rect 55036 472608 55088 472660
rect 67640 472608 67692 472660
rect 102232 472608 102284 472660
rect 143540 472608 143592 472660
rect 61936 471928 61988 471980
rect 63224 471928 63276 471980
rect 67640 471928 67692 471980
rect 102232 471928 102284 471980
rect 132592 471996 132644 472048
rect 102784 471316 102836 471368
rect 135444 471316 135496 471368
rect 143632 471316 143684 471368
rect 109040 471248 109092 471300
rect 146300 471248 146352 471300
rect 146300 470568 146352 470620
rect 579988 470568 580040 470620
rect 66168 469888 66220 469940
rect 67640 469888 67692 469940
rect 103520 469888 103572 469940
rect 131396 469888 131448 469940
rect 139492 469888 139544 469940
rect 46664 469820 46716 469872
rect 102232 469820 102284 469872
rect 134064 469820 134116 469872
rect 34244 469140 34296 469192
rect 66996 469140 67048 469192
rect 67548 469140 67600 469192
rect 64604 467848 64656 467900
rect 65984 467848 66036 467900
rect 67640 467848 67692 467900
rect 125508 467100 125560 467152
rect 133880 467100 133932 467152
rect 108396 466556 108448 466608
rect 113272 466556 113324 466608
rect 105636 466488 105688 466540
rect 107844 466488 107896 466540
rect 64696 466420 64748 466472
rect 67640 466420 67692 466472
rect 102232 466420 102284 466472
rect 125508 466420 125560 466472
rect 102324 465808 102376 465860
rect 107752 465808 107804 465860
rect 116584 465808 116636 465860
rect 102232 465740 102284 465792
rect 116032 465740 116084 465792
rect 116676 465740 116728 465792
rect 103520 465672 103572 465724
rect 136824 465672 136876 465724
rect 138112 465672 138164 465724
rect 67640 465060 67692 465112
rect 48044 464992 48096 465044
rect 50344 464992 50396 465044
rect 59176 464992 59228 465044
rect 63132 464992 63184 465044
rect 67732 464992 67784 465044
rect 104716 464108 104768 464160
rect 107660 464108 107712 464160
rect 67640 463700 67692 463752
rect 56508 463632 56560 463684
rect 57244 463632 57296 463684
rect 125600 463632 125652 463684
rect 125968 463632 126020 463684
rect 52460 462952 52512 463004
rect 53564 462952 53616 463004
rect 67640 462952 67692 463004
rect 102232 462952 102284 463004
rect 125600 462952 125652 463004
rect 2780 462544 2832 462596
rect 4804 462544 4856 462596
rect 61752 462340 61804 462392
rect 64604 462340 64656 462392
rect 67640 462340 67692 462392
rect 107568 462340 107620 462392
rect 140964 462340 141016 462392
rect 48228 462272 48280 462324
rect 52460 462272 52512 462324
rect 58992 462272 59044 462324
rect 63132 462272 63184 462324
rect 102324 462272 102376 462324
rect 129924 462272 129976 462324
rect 130384 462272 130436 462324
rect 102232 462204 102284 462256
rect 107568 462204 107620 462256
rect 116676 462204 116728 462256
rect 120724 462204 120776 462256
rect 63132 460912 63184 460964
rect 67640 460912 67692 460964
rect 102324 460844 102376 460896
rect 106648 460844 106700 460896
rect 102140 460300 102192 460352
rect 105544 460300 105596 460352
rect 54208 460232 54260 460284
rect 55128 460232 55180 460284
rect 67640 460232 67692 460284
rect 41236 460164 41288 460216
rect 67732 460164 67784 460216
rect 40960 459552 41012 459604
rect 41236 459552 41288 459604
rect 107016 459552 107068 459604
rect 114744 459552 114796 459604
rect 124956 459552 125008 459604
rect 133972 459552 134024 459604
rect 102140 459484 102192 459536
rect 108212 458804 108264 458856
rect 134248 458804 134300 458856
rect 149244 458804 149296 458856
rect 48044 458192 48096 458244
rect 54208 458192 54260 458244
rect 64788 458192 64840 458244
rect 67640 458192 67692 458244
rect 102140 458192 102192 458244
rect 102324 458124 102376 458176
rect 108212 458124 108264 458176
rect 115848 458124 115900 458176
rect 120080 458124 120132 458176
rect 103520 457444 103572 457496
rect 139584 457444 139636 457496
rect 142252 457444 142304 457496
rect 52460 456832 52512 456884
rect 53196 456832 53248 456884
rect 67640 456832 67692 456884
rect 42708 456696 42760 456748
rect 44824 456696 44876 456748
rect 67732 456764 67784 456816
rect 377404 456764 377456 456816
rect 580172 456764 580224 456816
rect 48136 456696 48188 456748
rect 52460 456696 52512 456748
rect 102140 456696 102192 456748
rect 142160 456696 142212 456748
rect 143448 456696 143500 456748
rect 143448 456016 143500 456068
rect 151912 456016 151964 456068
rect 30288 455404 30340 455456
rect 36544 455336 36596 455388
rect 67640 455404 67692 455456
rect 102876 455336 102928 455388
rect 105636 455336 105688 455388
rect 56324 455268 56376 455320
rect 56508 455268 56560 455320
rect 106188 454792 106240 454844
rect 114836 454792 114888 454844
rect 108212 454724 108264 454776
rect 138204 454724 138256 454776
rect 150532 454724 150584 454776
rect 56508 454656 56560 454708
rect 67640 454656 67692 454708
rect 102140 454656 102192 454708
rect 135352 454656 135404 454708
rect 102140 453976 102192 454028
rect 118976 453976 119028 454028
rect 102324 453908 102376 453960
rect 108212 453908 108264 453960
rect 55128 453364 55180 453416
rect 57704 453364 57756 453416
rect 67640 453364 67692 453416
rect 54944 453296 54996 453348
rect 67732 453296 67784 453348
rect 52092 451936 52144 451988
rect 54944 451936 54996 451988
rect 102140 451936 102192 451988
rect 115940 451936 115992 451988
rect 102508 451868 102560 451920
rect 134156 451868 134208 451920
rect 147772 451868 147824 451920
rect 101956 451188 102008 451240
rect 105728 451188 105780 451240
rect 100116 450508 100168 450560
rect 109132 450508 109184 450560
rect 61844 449896 61896 449948
rect 64420 449896 64472 449948
rect 67640 449896 67692 449948
rect 106924 449896 106976 449948
rect 122840 449896 122892 449948
rect 102324 449828 102376 449880
rect 102140 449760 102192 449812
rect 105360 449760 105412 449812
rect 63316 448536 63368 448588
rect 64696 448536 64748 448588
rect 67640 448536 67692 448588
rect 102140 447924 102192 447976
rect 107016 447924 107068 447976
rect 104716 447856 104768 447908
rect 114928 447856 114980 447908
rect 102324 447788 102376 447840
rect 127072 447788 127124 447840
rect 61384 447108 61436 447160
rect 67640 447108 67692 447160
rect 34336 446972 34388 447024
rect 60740 445748 60792 445800
rect 61752 445748 61804 445800
rect 67640 445748 67692 445800
rect 101036 445748 101088 445800
rect 102048 445748 102100 445800
rect 146392 445748 146444 445800
rect 102140 445680 102192 445732
rect 103704 445680 103756 445732
rect 104164 445680 104216 445732
rect 102324 445272 102376 445324
rect 104900 445272 104952 445324
rect 105636 445272 105688 445324
rect 104808 445068 104860 445120
rect 128544 445068 128596 445120
rect 37004 445000 37056 445052
rect 67640 445000 67692 445052
rect 102140 445000 102192 445052
rect 132684 445000 132736 445052
rect 142160 445000 142212 445052
rect 102324 443980 102376 444032
rect 104808 443980 104860 444032
rect 34336 443640 34388 443692
rect 67640 443640 67692 443692
rect 113088 443640 113140 443692
rect 123116 443640 123168 443692
rect 33048 442892 33100 442944
rect 34152 442892 34204 442944
rect 67640 442892 67692 442944
rect 49608 442824 49660 442876
rect 66260 442824 66312 442876
rect 60280 442756 60332 442808
rect 61844 442756 61896 442808
rect 67732 442756 67784 442808
rect 64420 442280 64472 442332
rect 64788 442280 64840 442332
rect 102140 441600 102192 441652
rect 62028 441532 62080 441584
rect 63316 441532 63368 441584
rect 63408 441532 63460 441584
rect 66168 441532 66220 441584
rect 129832 441532 129884 441584
rect 66168 441124 66220 441176
rect 67640 441124 67692 441176
rect 63316 440988 63368 441040
rect 67640 440988 67692 441040
rect 56232 440920 56284 440972
rect 43812 440852 43864 440904
rect 116124 440852 116176 440904
rect 129832 440852 129884 440904
rect 139584 440852 139636 440904
rect 71780 440648 71832 440700
rect 72332 440648 72384 440700
rect 79324 440648 79376 440700
rect 94136 440648 94188 440700
rect 97448 440648 97500 440700
rect 99932 440648 99984 440700
rect 100760 440308 100812 440360
rect 131120 440308 131172 440360
rect 99472 440240 99524 440292
rect 100852 440240 100904 440292
rect 136824 440240 136876 440292
rect 95332 440172 95384 440224
rect 100116 440172 100168 440224
rect 97908 440104 97960 440156
rect 103612 440104 103664 440156
rect 97264 439900 97316 439952
rect 69204 439560 69256 439612
rect 76564 439560 76616 439612
rect 95148 439560 95200 439612
rect 110604 439560 110656 439612
rect 50712 439492 50764 439544
rect 79324 439492 79376 439544
rect 81440 439492 81492 439544
rect 96528 439492 96580 439544
rect 120448 439492 120500 439544
rect 69112 439016 69164 439068
rect 73804 439016 73856 439068
rect 79784 439016 79836 439068
rect 82820 439016 82872 439068
rect 46756 438948 46808 439000
rect 80980 438948 81032 439000
rect 88708 438948 88760 439000
rect 121644 438948 121696 439000
rect 25504 438880 25556 438932
rect 96620 438880 96672 438932
rect 97724 438880 97776 438932
rect 75184 438812 75236 438864
rect 82268 438812 82320 438864
rect 86132 438812 86184 438864
rect 94504 438812 94556 438864
rect 95148 438812 95200 438864
rect 96436 438812 96488 438864
rect 50896 438744 50948 438796
rect 82912 438744 82964 438796
rect 84200 438744 84252 438796
rect 85580 438744 85632 438796
rect 91284 438744 91336 438796
rect 95240 438744 95292 438796
rect 96528 438744 96580 438796
rect 99012 438812 99064 438864
rect 121736 438812 121788 438864
rect 124220 438812 124272 438864
rect 123024 438744 123076 438796
rect 52000 438676 52052 438728
rect 83556 438676 83608 438728
rect 70400 438608 70452 438660
rect 77116 438608 77168 438660
rect 88248 438608 88300 438660
rect 105728 438608 105780 438660
rect 3424 438540 3476 438592
rect 99380 438540 99432 438592
rect 93584 438472 93636 438524
rect 93952 438472 94004 438524
rect 87420 438268 87472 438320
rect 88248 438268 88300 438320
rect 56324 438200 56376 438252
rect 73896 438200 73948 438252
rect 4804 438132 4856 438184
rect 49516 438132 49568 438184
rect 52000 438132 52052 438184
rect 52460 438132 52512 438184
rect 71320 438132 71372 438184
rect 85580 438132 85632 438184
rect 118884 438132 118936 438184
rect 98368 437996 98420 438048
rect 99288 437996 99340 438048
rect 102232 437996 102284 438048
rect 69112 437452 69164 437504
rect 73252 437452 73304 437504
rect 85028 437452 85080 437504
rect 86776 437452 86828 437504
rect 88064 437452 88116 437504
rect 89628 437452 89680 437504
rect 47952 437384 48004 437436
rect 78680 437384 78732 437436
rect 79048 437384 79100 437436
rect 89996 437384 90048 437436
rect 90364 437384 90416 437436
rect 124404 437384 124456 437436
rect 39856 437316 39908 437368
rect 69112 437316 69164 437368
rect 94964 437316 95016 437368
rect 125784 437316 125836 437368
rect 37188 437248 37240 437300
rect 52460 437248 52512 437300
rect 53104 437248 53156 437300
rect 53656 437248 53708 437300
rect 74632 437248 74684 437300
rect 75828 437248 75880 437300
rect 89352 437248 89404 437300
rect 89536 437248 89588 437300
rect 108396 437248 108448 437300
rect 54852 437180 54904 437232
rect 70400 437180 70452 437232
rect 93216 437180 93268 437232
rect 93676 437180 93728 437232
rect 108488 437180 108540 437232
rect 45468 437112 45520 437164
rect 55864 437112 55916 437164
rect 56324 437112 56376 437164
rect 64512 436704 64564 436756
rect 75184 436704 75236 436756
rect 59084 436024 59136 436076
rect 91744 436024 91796 436076
rect 92572 436024 92624 436076
rect 93768 436024 93820 436076
rect 124312 436024 124364 436076
rect 46848 435956 46900 436008
rect 78588 435956 78640 436008
rect 89628 435956 89680 436008
rect 112076 435956 112128 436008
rect 65524 435344 65576 435396
rect 77944 435344 77996 435396
rect 41052 434664 41104 434716
rect 41236 434664 41288 434716
rect 42524 434664 42576 434716
rect 74540 434664 74592 434716
rect 70676 434596 70728 434648
rect 49332 434528 49384 434580
rect 49608 434528 49660 434580
rect 76472 434528 76524 434580
rect 45284 433984 45336 434036
rect 49608 433984 49660 434036
rect 78588 431944 78640 431996
rect 80152 431944 80204 431996
rect 580908 431944 580960 431996
rect 39672 431876 39724 431928
rect 71872 431876 71924 431928
rect 100760 430584 100812 430636
rect 101956 430584 102008 430636
rect 104256 430584 104308 430636
rect 3424 429836 3476 429888
rect 100760 429836 100812 429888
rect 3516 422288 3568 422340
rect 118792 422220 118844 422272
rect 121644 404336 121696 404388
rect 579620 404336 579672 404388
rect 70400 404268 70452 404320
rect 71044 404268 71096 404320
rect 93584 403656 93636 403708
rect 129924 403656 129976 403708
rect 104164 403588 104216 403640
rect 141056 403588 141108 403640
rect 70400 402976 70452 403028
rect 341524 402976 341576 403028
rect 74816 401616 74868 401668
rect 304264 401616 304316 401668
rect 96620 400868 96672 400920
rect 132684 400868 132736 400920
rect 89536 399576 89588 399628
rect 125968 399576 126020 399628
rect 41144 399508 41196 399560
rect 86224 399508 86276 399560
rect 93676 399508 93728 399560
rect 127256 399508 127308 399560
rect 39764 399440 39816 399492
rect 85120 399440 85172 399492
rect 92664 399440 92716 399492
rect 125876 399440 125928 399492
rect 198004 399440 198056 399492
rect 65984 398828 66036 398880
rect 170404 398828 170456 398880
rect 100668 398760 100720 398812
rect 104164 398760 104216 398812
rect 104256 398216 104308 398268
rect 135444 398216 135496 398268
rect 97264 398148 97316 398200
rect 130016 398148 130068 398200
rect 43996 398080 44048 398132
rect 77300 398080 77352 398132
rect 91744 398080 91796 398132
rect 128544 398080 128596 398132
rect 128360 397672 128412 397724
rect 128728 397672 128780 397724
rect 128360 397536 128412 397588
rect 129004 397536 129056 397588
rect 215944 397536 215996 397588
rect 61936 397468 61988 397520
rect 291844 397468 291896 397520
rect 77944 397400 77996 397452
rect 121644 397400 121696 397452
rect 39856 396788 39908 396840
rect 56416 396856 56468 396908
rect 89720 396856 89772 396908
rect 93768 396856 93820 396908
rect 128636 396856 128688 396908
rect 84108 396788 84160 396840
rect 120816 396788 120868 396840
rect 42616 396720 42668 396772
rect 88340 396720 88392 396772
rect 94136 396720 94188 396772
rect 128360 396720 128412 396772
rect 88340 396040 88392 396092
rect 195244 396040 195296 396092
rect 43904 395428 43956 395480
rect 50988 395428 51040 395480
rect 59268 395428 59320 395480
rect 84200 395428 84252 395480
rect 89720 395428 89772 395480
rect 103796 395428 103848 395480
rect 43720 395360 43772 395412
rect 82820 395360 82872 395412
rect 95148 395360 95200 395412
rect 125784 395360 125836 395412
rect 38476 395292 38528 395344
rect 81440 395292 81492 395344
rect 98000 395292 98052 395344
rect 131304 395292 131356 395344
rect 322940 395292 322992 395344
rect 82820 394748 82872 394800
rect 83096 394748 83148 394800
rect 139400 394748 139452 394800
rect 50988 394680 51040 394732
rect 84200 394680 84252 394732
rect 103520 394680 103572 394732
rect 104716 394680 104768 394732
rect 206284 394680 206336 394732
rect 109776 394612 109828 394664
rect 111984 394612 112036 394664
rect 110880 394136 110932 394188
rect 129740 394136 129792 394188
rect 93860 394068 93912 394120
rect 128728 394068 128780 394120
rect 45376 394000 45428 394052
rect 57612 394000 57664 394052
rect 96712 394000 96764 394052
rect 131212 394000 131264 394052
rect 46572 393932 46624 393984
rect 82912 393932 82964 393984
rect 88248 393932 88300 393984
rect 124312 393932 124364 393984
rect 128728 393932 128780 393984
rect 129740 393932 129792 393984
rect 150440 393932 150492 393984
rect 57612 393456 57664 393508
rect 91100 393456 91152 393508
rect 39764 393388 39816 393440
rect 110880 393388 110932 393440
rect 85120 393320 85172 393372
rect 260104 393320 260156 393372
rect 105544 392776 105596 392828
rect 117596 392776 117648 392828
rect 110328 392708 110380 392760
rect 132500 392708 132552 392760
rect 136640 392708 136692 392760
rect 56416 392640 56468 392692
rect 74540 392640 74592 392692
rect 96528 392640 96580 392692
rect 123024 392640 123076 392692
rect 3424 392572 3476 392624
rect 116124 392436 116176 392488
rect 118700 392436 118752 392488
rect 111064 392028 111116 392080
rect 113640 392028 113692 392080
rect 67456 391960 67508 392012
rect 298744 391960 298796 392012
rect 99288 391280 99340 391332
rect 120172 391280 120224 391332
rect 53288 391212 53340 391264
rect 75460 391212 75512 391264
rect 96528 391212 96580 391264
rect 127164 391212 127216 391264
rect 142436 391212 142488 391264
rect 120080 390736 120132 390788
rect 120724 390736 120776 390788
rect 127164 390736 127216 390788
rect 49608 390668 49660 390720
rect 77944 390668 77996 390720
rect 81440 390668 81492 390720
rect 82544 390668 82596 390720
rect 143724 390668 143776 390720
rect 75460 390600 75512 390652
rect 140780 390600 140832 390652
rect 72424 390532 72476 390584
rect 146576 390532 146628 390584
rect 58900 390056 58952 390108
rect 104532 390056 104584 390108
rect 70308 389988 70360 390040
rect 79324 389988 79376 390040
rect 69848 389920 69900 389972
rect 85580 389920 85632 389972
rect 118792 389920 118844 389972
rect 131212 389920 131264 389972
rect 57336 389852 57388 389904
rect 120080 389852 120132 389904
rect 52184 389784 52236 389836
rect 58900 389784 58952 389836
rect 99380 389784 99432 389836
rect 111800 389784 111852 389836
rect 334716 389784 334768 389836
rect 111708 389580 111760 389632
rect 114836 389580 114888 389632
rect 115572 389444 115624 389496
rect 118792 389444 118844 389496
rect 101312 389308 101364 389360
rect 133880 389308 133932 389360
rect 50804 389240 50856 389292
rect 53748 389240 53800 389292
rect 79324 389240 79376 389292
rect 114284 389240 114336 389292
rect 146484 389240 146536 389292
rect 42984 389172 43036 389224
rect 43444 389172 43496 389224
rect 71780 389172 71832 389224
rect 113640 389172 113692 389224
rect 262864 389172 262916 389224
rect 36636 389104 36688 389156
rect 37096 389104 37148 389156
rect 72424 389104 72476 389156
rect 39948 389036 40000 389088
rect 42984 389036 43036 389088
rect 90272 388560 90324 388612
rect 99380 388560 99432 388612
rect 88248 388492 88300 388544
rect 103520 388492 103572 388544
rect 107016 388492 107068 388544
rect 135260 388492 135312 388544
rect 136548 388492 136600 388544
rect 4804 388424 4856 388476
rect 36636 388424 36688 388476
rect 91008 388424 91060 388476
rect 113088 388424 113140 388476
rect 313924 388424 313976 388476
rect 102600 388356 102652 388408
rect 106188 388356 106240 388408
rect 73528 388084 73580 388136
rect 73804 388084 73856 388136
rect 122196 388084 122248 388136
rect 109684 388016 109736 388068
rect 119436 388016 119488 388068
rect 52276 387948 52328 388000
rect 92940 387948 92992 388000
rect 101404 387948 101456 388000
rect 119344 387948 119396 388000
rect 35532 387880 35584 387932
rect 35716 387880 35768 387932
rect 80060 387880 80112 387932
rect 100024 387880 100076 387932
rect 119528 387880 119580 387932
rect 58532 387812 58584 387864
rect 70216 387812 70268 387864
rect 106188 387812 106240 387864
rect 108764 387812 108816 387864
rect 69664 387336 69716 387388
rect 78680 387336 78732 387388
rect 47952 387268 48004 387320
rect 71872 387268 71924 387320
rect 52368 387200 52420 387252
rect 80612 387200 80664 387252
rect 89628 387200 89680 387252
rect 118700 387200 118752 387252
rect 59084 387132 59136 387184
rect 90364 387132 90416 387184
rect 108304 387132 108356 387184
rect 117412 387132 117464 387184
rect 60648 387064 60700 387116
rect 95240 387064 95292 387116
rect 99288 387064 99340 387116
rect 127348 387064 127400 387116
rect 127532 387064 127584 387116
rect 54944 386452 54996 386504
rect 87052 386452 87104 386504
rect 103704 386452 103756 386504
rect 104164 386452 104216 386504
rect 138204 386452 138256 386504
rect 76656 386384 76708 386436
rect 327724 386384 327776 386436
rect 121368 386316 121420 386368
rect 121552 386316 121604 386368
rect 66076 386248 66128 386300
rect 68744 386248 68796 386300
rect 53564 385704 53616 385756
rect 80152 385976 80204 386028
rect 105636 385704 105688 385756
rect 131304 385704 131356 385756
rect 41328 385636 41380 385688
rect 113364 385636 113416 385688
rect 117228 385636 117280 385688
rect 122288 385636 122340 385688
rect 136916 385636 136968 385688
rect 112168 385364 112220 385416
rect 52368 385024 52420 385076
rect 107108 385296 107160 385348
rect 108948 385296 109000 385348
rect 122104 385296 122156 385348
rect 122288 385296 122340 385348
rect 324964 385024 325016 385076
rect 116032 384344 116084 384396
rect 122932 384344 122984 384396
rect 118608 384276 118660 384328
rect 249064 384276 249116 384328
rect 34244 383664 34296 383716
rect 68744 383664 68796 383716
rect 35808 382236 35860 382288
rect 67640 382236 67692 382288
rect 116216 382236 116268 382288
rect 145012 382236 145064 382288
rect 118608 382168 118660 382220
rect 142344 382168 142396 382220
rect 143448 382168 143500 382220
rect 118608 381556 118660 381608
rect 147680 381556 147732 381608
rect 143448 381488 143500 381540
rect 204904 381488 204956 381540
rect 147680 380876 147732 380928
rect 147956 380876 148008 380928
rect 42800 380808 42852 380860
rect 44088 380808 44140 380860
rect 67640 380808 67692 380860
rect 60372 380740 60424 380792
rect 68008 380740 68060 380792
rect 35624 380196 35676 380248
rect 60188 380196 60240 380248
rect 18604 380128 18656 380180
rect 42800 380128 42852 380180
rect 118608 379584 118660 379636
rect 124496 379584 124548 379636
rect 128360 379584 128412 379636
rect 60188 379516 60240 379568
rect 60464 379516 60516 379568
rect 67640 379516 67692 379568
rect 118516 379516 118568 379568
rect 342904 379516 342956 379568
rect 118608 378836 118660 378888
rect 123116 378836 123168 378888
rect 65156 378768 65208 378820
rect 67640 378768 67692 378820
rect 119528 378768 119580 378820
rect 346400 378768 346452 378820
rect 117872 378156 117924 378208
rect 121552 378156 121604 378208
rect 121552 377544 121604 377596
rect 125876 377544 125928 377596
rect 119528 377408 119580 377460
rect 125692 377408 125744 377460
rect 118608 376796 118660 376848
rect 119528 376796 119580 376848
rect 55036 376660 55088 376712
rect 65524 376728 65576 376780
rect 67640 376728 67692 376780
rect 125876 376728 125928 376780
rect 372620 376728 372672 376780
rect 149060 376660 149112 376712
rect 150624 376660 150676 376712
rect 61936 376592 61988 376644
rect 67640 376592 67692 376644
rect 55036 375980 55088 376032
rect 70308 375980 70360 376032
rect 66996 375844 67048 375896
rect 67640 375844 67692 375896
rect 118608 375368 118660 375420
rect 149060 375368 149112 375420
rect 46664 375300 46716 375352
rect 69112 375300 69164 375352
rect 118148 375300 118200 375352
rect 147680 375300 147732 375352
rect 147864 375300 147916 375352
rect 63408 374620 63460 374672
rect 67640 374620 67692 374672
rect 147680 374620 147732 374672
rect 191104 374620 191156 374672
rect 58992 373940 59044 373992
rect 67640 373940 67692 373992
rect 65984 373124 66036 373176
rect 67640 373124 67692 373176
rect 118332 372648 118384 372700
rect 120172 372648 120224 372700
rect 118516 372580 118568 372632
rect 331864 372580 331916 372632
rect 3240 372512 3292 372564
rect 57336 372512 57388 372564
rect 118148 371220 118200 371272
rect 421564 371220 421616 371272
rect 120172 371152 120224 371204
rect 151820 371152 151872 371204
rect 153108 371152 153160 371204
rect 64512 370608 64564 370660
rect 67640 370608 67692 370660
rect 50344 370540 50396 370592
rect 67272 370540 67324 370592
rect 67732 370540 67784 370592
rect 50804 370472 50856 370524
rect 69756 370472 69808 370524
rect 115940 369928 115992 369980
rect 120172 369928 120224 369980
rect 118148 369860 118200 369912
rect 151820 369860 151872 369912
rect 57244 369112 57296 369164
rect 67640 369112 67692 369164
rect 118608 368500 118660 368552
rect 124404 368500 124456 368552
rect 128452 368500 128504 368552
rect 59176 367820 59228 367872
rect 67916 367820 67968 367872
rect 118608 367820 118660 367872
rect 121460 367820 121512 367872
rect 134524 367820 134576 367872
rect 58992 367752 59044 367804
rect 69664 367752 69716 367804
rect 124128 367752 124180 367804
rect 144920 367752 144972 367804
rect 479524 367752 479576 367804
rect 579620 367752 579672 367804
rect 118608 367208 118660 367260
rect 122932 367208 122984 367260
rect 124128 367208 124180 367260
rect 48228 367004 48280 367056
rect 60188 367004 60240 367056
rect 120172 367004 120224 367056
rect 137008 367004 137060 367056
rect 137192 367004 137244 367056
rect 64604 366392 64656 366444
rect 68468 366392 68520 366444
rect 118608 366392 118660 366444
rect 143540 366392 143592 366444
rect 60188 366324 60240 366376
rect 67640 366324 67692 366376
rect 137192 366324 137244 366376
rect 579620 366324 579672 366376
rect 37188 365644 37240 365696
rect 40960 365644 41012 365696
rect 60556 365712 60608 365764
rect 120816 365644 120868 365696
rect 121460 365644 121512 365696
rect 118608 365032 118660 365084
rect 132592 365032 132644 365084
rect 63132 364964 63184 365016
rect 68560 364964 68612 365016
rect 120724 364964 120776 365016
rect 146300 364964 146352 365016
rect 118516 364352 118568 364404
rect 120724 364352 120776 364404
rect 121460 364352 121512 364404
rect 579804 364352 579856 364404
rect 60556 364284 60608 364336
rect 67732 364284 67784 364336
rect 48044 363604 48096 363656
rect 67640 363604 67692 363656
rect 117412 363604 117464 363656
rect 282184 363604 282236 363656
rect 48044 363060 48096 363112
rect 48228 363060 48280 363112
rect 118608 362856 118660 362908
rect 143632 362856 143684 362908
rect 144828 362856 144880 362908
rect 118608 362176 118660 362228
rect 119988 362176 120040 362228
rect 134064 362176 134116 362228
rect 144828 362176 144880 362228
rect 202144 362176 202196 362228
rect 116584 361972 116636 362024
rect 117320 361972 117372 362024
rect 32956 361496 33008 361548
rect 36544 361564 36596 361616
rect 67640 361496 67692 361548
rect 44824 360816 44876 360868
rect 45468 360816 45520 360868
rect 67640 360816 67692 360868
rect 125508 360272 125560 360324
rect 128452 360272 128504 360324
rect 118056 360204 118108 360256
rect 135904 360204 135956 360256
rect 139492 360204 139544 360256
rect 117964 360136 118016 360188
rect 152004 360136 152056 360188
rect 153108 360136 153160 360188
rect 118608 360068 118660 360120
rect 125508 360068 125560 360120
rect 68560 359524 68612 359576
rect 68928 359524 68980 359576
rect 53196 359456 53248 359508
rect 53656 359456 53708 359508
rect 67640 359456 67692 359508
rect 68468 359456 68520 359508
rect 68836 359456 68888 359508
rect 153108 359456 153160 359508
rect 188344 359456 188396 359508
rect 3332 358708 3384 358760
rect 37004 358708 37056 358760
rect 43536 358708 43588 358760
rect 56508 358708 56560 358760
rect 59360 358708 59412 358760
rect 118608 358708 118660 358760
rect 127164 358708 127216 358760
rect 129832 358708 129884 358760
rect 30288 358028 30340 358080
rect 65984 358028 66036 358080
rect 67640 358028 67692 358080
rect 59360 357416 59412 357468
rect 67640 357416 67692 357468
rect 115848 357348 115900 357400
rect 117412 357348 117464 357400
rect 118608 357348 118660 357400
rect 138112 357348 138164 357400
rect 140872 357348 140924 357400
rect 42708 356668 42760 356720
rect 67640 356668 67692 356720
rect 118240 356668 118292 356720
rect 340144 356668 340196 356720
rect 55128 355988 55180 356040
rect 61476 355988 61528 356040
rect 67640 355988 67692 356040
rect 52092 355308 52144 355360
rect 59176 355308 59228 355360
rect 119344 355308 119396 355360
rect 580264 355308 580316 355360
rect 59176 354696 59228 354748
rect 67640 354696 67692 354748
rect 118608 354628 118660 354680
rect 140964 354628 141016 354680
rect 117504 354560 117556 354612
rect 125600 354560 125652 354612
rect 140964 354016 141016 354068
rect 147680 354016 147732 354068
rect 118792 353948 118844 354000
rect 297364 353948 297416 354000
rect 125600 353268 125652 353320
rect 126980 353268 127032 353320
rect 117504 353200 117556 353252
rect 134064 353200 134116 353252
rect 146300 353268 146352 353320
rect 64788 352588 64840 352640
rect 67640 352588 67692 352640
rect 7564 352520 7616 352572
rect 68560 352520 68612 352572
rect 482284 352520 482336 352572
rect 579620 352520 579672 352572
rect 118056 351840 118108 351892
rect 138020 351840 138072 351892
rect 138020 351228 138072 351280
rect 196624 351228 196676 351280
rect 64696 351160 64748 351212
rect 68008 351160 68060 351212
rect 118608 351160 118660 351212
rect 318064 351160 318116 351212
rect 49424 350548 49476 350600
rect 53840 350548 53892 350600
rect 53840 349800 53892 349852
rect 55128 349800 55180 349852
rect 67640 349800 67692 349852
rect 122196 349800 122248 349852
rect 346492 349800 346544 349852
rect 61384 349120 61436 349172
rect 64420 349120 64472 349172
rect 67640 349120 67692 349172
rect 117504 349120 117556 349172
rect 119436 349120 119488 349172
rect 46848 349052 46900 349104
rect 48136 349052 48188 349104
rect 63224 348440 63276 348492
rect 67640 348440 67692 348492
rect 48136 348372 48188 348424
rect 63500 348372 63552 348424
rect 118516 348372 118568 348424
rect 320824 348372 320876 348424
rect 63500 347692 63552 347744
rect 67640 347692 67692 347744
rect 118608 347692 118660 347744
rect 151912 347692 151964 347744
rect 153108 347692 153160 347744
rect 153108 347012 153160 347064
rect 184204 347012 184256 347064
rect 118608 346332 118660 346384
rect 135352 346332 135404 346384
rect 136548 346332 136600 346384
rect 2780 346264 2832 346316
rect 4804 346264 4856 346316
rect 118516 345720 118568 345772
rect 142252 345720 142304 345772
rect 43536 345652 43588 345704
rect 61936 345652 61988 345704
rect 136548 345652 136600 345704
rect 186964 345652 187016 345704
rect 61936 345108 61988 345160
rect 67640 345108 67692 345160
rect 56324 345040 56376 345092
rect 67088 345040 67140 345092
rect 68008 344972 68060 345024
rect 117964 344972 118016 345024
rect 149244 344972 149296 345024
rect 149244 344292 149296 344344
rect 349896 344292 349948 344344
rect 62120 343612 62172 343664
rect 67640 343612 67692 343664
rect 117872 343612 117924 343664
rect 244924 343612 244976 343664
rect 34336 342864 34388 342916
rect 41144 342864 41196 342916
rect 62120 342864 62172 342916
rect 118608 342864 118660 342916
rect 130108 342864 130160 342916
rect 61844 342252 61896 342304
rect 66076 342252 66128 342304
rect 67640 342252 67692 342304
rect 118608 342184 118660 342236
rect 150532 342184 150584 342236
rect 150992 342184 151044 342236
rect 66168 341572 66220 341624
rect 68652 341572 68704 341624
rect 150992 341504 151044 341556
rect 348424 341504 348476 341556
rect 33048 340756 33100 340808
rect 64144 340892 64196 340944
rect 67640 340892 67692 340944
rect 118056 340892 118108 340944
rect 142252 340892 142304 340944
rect 63316 340824 63368 340876
rect 68652 340824 68704 340876
rect 117964 340824 118016 340876
rect 147772 340824 147824 340876
rect 118608 340756 118660 340808
rect 135444 340756 135496 340808
rect 138020 340756 138072 340808
rect 147772 340144 147824 340196
rect 338764 340144 338816 340196
rect 69020 340008 69072 340060
rect 69756 340008 69808 340060
rect 71780 339872 71832 339924
rect 72424 339872 72476 339924
rect 43904 339464 43956 339516
rect 78404 339464 78456 339516
rect 97724 339464 97776 339516
rect 129924 339464 129976 339516
rect 42524 339396 42576 339448
rect 75184 339396 75236 339448
rect 75828 339396 75880 339448
rect 87420 339396 87472 339448
rect 87696 339396 87748 339448
rect 121460 339396 121512 339448
rect 46756 339328 46808 339380
rect 50712 339328 50764 339380
rect 99656 339328 99708 339380
rect 100668 339328 100720 339380
rect 130016 339328 130068 339380
rect 67364 338852 67416 338904
rect 77944 338852 77996 338904
rect 78404 338784 78456 338836
rect 93124 338784 93176 338836
rect 64788 338716 64840 338768
rect 87604 338716 87656 338768
rect 50712 338104 50764 338156
rect 43996 338036 44048 338088
rect 79048 338036 79100 338088
rect 82268 338036 82320 338088
rect 106188 338036 106240 338088
rect 131120 338036 131172 338088
rect 57888 337968 57940 338020
rect 84200 337968 84252 338020
rect 100300 337968 100352 338020
rect 123024 337968 123076 338020
rect 56416 337900 56468 337952
rect 76472 337900 76524 337952
rect 113824 337900 113876 337952
rect 127072 337900 127124 337952
rect 55864 337832 55916 337884
rect 74540 337832 74592 337884
rect 75276 337832 75328 337884
rect 103520 337560 103572 337612
rect 114468 337560 114520 337612
rect 50896 337356 50948 337408
rect 60556 337356 60608 337408
rect 84844 337492 84896 337544
rect 93952 337492 94004 337544
rect 123116 337492 123168 337544
rect 79048 337424 79100 337476
rect 220084 337424 220136 337476
rect 68560 337356 68612 337408
rect 322204 337356 322256 337408
rect 59084 336676 59136 336728
rect 92480 336676 92532 336728
rect 108028 336676 108080 336728
rect 139584 336676 139636 336728
rect 39672 336608 39724 336660
rect 71964 336608 72016 336660
rect 72516 336608 72568 336660
rect 115112 336608 115164 336660
rect 115296 336608 115348 336660
rect 119436 336608 119488 336660
rect 133972 336608 134024 336660
rect 135168 336608 135220 336660
rect 55036 336540 55088 336592
rect 83464 336540 83516 336592
rect 122840 336540 122892 336592
rect 123484 336540 123536 336592
rect 124220 336540 124272 336592
rect 53564 336472 53616 336524
rect 79324 336472 79376 336524
rect 47952 336404 48004 336456
rect 73344 336404 73396 336456
rect 92480 335996 92532 336048
rect 93216 335996 93268 336048
rect 104164 335996 104216 336048
rect 114468 335996 114520 336048
rect 123484 335996 123536 336048
rect 135168 335996 135220 336048
rect 269764 335996 269816 336048
rect 46572 335248 46624 335300
rect 81624 335248 81676 335300
rect 115204 335248 115256 335300
rect 149152 335248 149204 335300
rect 50804 335180 50856 335232
rect 86776 335180 86828 335232
rect 109960 335180 110012 335232
rect 128820 335180 128872 335232
rect 133972 335180 134024 335232
rect 60648 335112 60700 335164
rect 94504 335112 94556 335164
rect 102876 335112 102928 335164
rect 103428 335112 103480 335164
rect 120080 335112 120132 335164
rect 58992 335044 59044 335096
rect 80980 335044 81032 335096
rect 86316 334636 86368 334688
rect 86776 334636 86828 334688
rect 100024 334636 100076 334688
rect 124404 334636 124456 334688
rect 56508 334568 56560 334620
rect 119436 334568 119488 334620
rect 81624 333956 81676 334008
rect 82084 333956 82136 334008
rect 49516 333888 49568 333940
rect 86224 333888 86276 333940
rect 97080 333888 97132 333940
rect 127256 333888 127308 333940
rect 57704 333276 57756 333328
rect 87696 333276 87748 333328
rect 95148 333276 95200 333328
rect 113824 333276 113876 333328
rect 68744 333208 68796 333260
rect 309784 333208 309836 333260
rect 97080 332732 97132 332784
rect 97908 332732 97960 332784
rect 108304 332528 108356 332580
rect 142160 332528 142212 332580
rect 143448 332528 143500 332580
rect 61936 331916 61988 331968
rect 98644 331916 98696 331968
rect 64144 331848 64196 331900
rect 124220 331848 124272 331900
rect 143448 331848 143500 331900
rect 409880 331848 409932 331900
rect 59268 331168 59320 331220
rect 88984 331168 89036 331220
rect 105452 331168 105504 331220
rect 136824 331168 136876 331220
rect 137100 331168 137152 331220
rect 60464 330488 60516 330540
rect 115204 330488 115256 330540
rect 137100 330488 137152 330540
rect 425704 330488 425756 330540
rect 88708 329740 88760 329792
rect 122012 329740 122064 329792
rect 92572 329672 92624 329724
rect 125968 329672 126020 329724
rect 126888 329672 126940 329724
rect 69204 329128 69256 329180
rect 121460 329128 121512 329180
rect 48136 329060 48188 329112
rect 108028 329060 108080 329112
rect 126888 329060 126940 329112
rect 295984 329060 296036 329112
rect 4804 328448 4856 328500
rect 48136 328448 48188 328500
rect 122012 328448 122064 328500
rect 216036 328448 216088 328500
rect 106096 327904 106148 327956
rect 116032 327904 116084 327956
rect 91928 327836 91980 327888
rect 125600 327836 125652 327888
rect 66076 327768 66128 327820
rect 269856 327768 269908 327820
rect 78036 327700 78088 327752
rect 358084 327700 358136 327752
rect 112536 327020 112588 327072
rect 146392 327020 146444 327072
rect 146760 327020 146812 327072
rect 76564 326476 76616 326528
rect 122196 326476 122248 326528
rect 71044 326340 71096 326392
rect 122104 326340 122156 326392
rect 214564 326408 214616 326460
rect 146760 326340 146812 326392
rect 254584 326340 254636 326392
rect 63224 325048 63276 325100
rect 177304 325048 177356 325100
rect 82084 324980 82136 325032
rect 268384 324980 268436 325032
rect 72516 324912 72568 324964
rect 300124 324912 300176 324964
rect 95792 324232 95844 324284
rect 128636 324232 128688 324284
rect 73160 323552 73212 323604
rect 115940 323552 115992 323604
rect 128636 323552 128688 323604
rect 395344 323552 395396 323604
rect 110604 322872 110656 322924
rect 140964 322872 141016 322924
rect 140964 322260 141016 322312
rect 302884 322260 302936 322312
rect 86316 322192 86368 322244
rect 399484 322192 399536 322244
rect 89996 321512 90048 321564
rect 124312 321512 124364 321564
rect 125508 321512 125560 321564
rect 67548 320900 67600 320952
rect 116124 320900 116176 320952
rect 125508 320900 125560 320952
rect 267004 320900 267056 320952
rect 68836 320832 68888 320884
rect 336096 320832 336148 320884
rect 100944 320084 100996 320136
rect 132776 320084 132828 320136
rect 133788 320084 133840 320136
rect 93768 319540 93820 319592
rect 115296 319540 115348 319592
rect 3240 319472 3292 319524
rect 18604 319472 18656 319524
rect 101404 319472 101456 319524
rect 133788 319472 133840 319524
rect 216128 319472 216180 319524
rect 68928 319404 68980 319456
rect 343640 319404 343692 319456
rect 91284 318724 91336 318776
rect 118700 318724 118752 318776
rect 111248 318656 111300 318708
rect 131304 318656 131356 318708
rect 131672 318656 131724 318708
rect 131672 318112 131724 318164
rect 265624 318112 265676 318164
rect 75276 318044 75328 318096
rect 115296 318044 115348 318096
rect 118700 318044 118752 318096
rect 267096 318044 267148 318096
rect 102232 317364 102284 317416
rect 132684 317364 132736 317416
rect 133788 317364 133840 317416
rect 72516 316684 72568 316736
rect 108304 316684 108356 316736
rect 133788 316684 133840 316736
rect 345020 316684 345072 316736
rect 84292 316072 84344 316124
rect 113180 316072 113232 316124
rect 69204 316004 69256 316056
rect 104256 316004 104308 316056
rect 72424 315256 72476 315308
rect 159364 315256 159416 315308
rect 91100 314644 91152 314696
rect 231124 314644 231176 314696
rect 57612 313964 57664 314016
rect 80060 313964 80112 314016
rect 91100 313964 91152 314016
rect 93124 313964 93176 314016
rect 151084 313964 151136 314016
rect 67456 313896 67508 313948
rect 125876 313896 125928 313948
rect 81440 313284 81492 313336
rect 226984 313284 227036 313336
rect 65524 311856 65576 311908
rect 66168 311856 66220 311908
rect 264244 311856 264296 311908
rect 453304 311856 453356 311908
rect 579988 311856 580040 311908
rect 101404 311244 101456 311296
rect 116584 311244 116636 311296
rect 87604 311176 87656 311228
rect 162124 311176 162176 311228
rect 115848 311108 115900 311160
rect 135904 311108 135956 311160
rect 271144 311108 271196 311160
rect 84384 309884 84436 309936
rect 115848 309884 115900 309936
rect 104900 309816 104952 309868
rect 145012 309816 145064 309868
rect 445760 309816 445812 309868
rect 113180 309748 113232 309800
rect 433340 309748 433392 309800
rect 75920 309136 75972 309188
rect 155316 309136 155368 309188
rect 104256 309068 104308 309120
rect 138204 309068 138256 309120
rect 138664 309068 138716 309120
rect 74448 308456 74500 308508
rect 121552 308456 121604 308508
rect 138664 308456 138716 308508
rect 262956 308456 263008 308508
rect 83464 308388 83516 308440
rect 345664 308388 345716 308440
rect 88340 307776 88392 307828
rect 153844 307776 153896 307828
rect 94228 307708 94280 307760
rect 94596 307708 94648 307760
rect 128544 307708 128596 307760
rect 128728 307708 128780 307760
rect 128728 307164 128780 307216
rect 155224 307164 155276 307216
rect 97908 307096 97960 307148
rect 334624 307096 334676 307148
rect 106188 307028 106240 307080
rect 113824 307028 113876 307080
rect 118700 307028 118752 307080
rect 146576 307028 146628 307080
rect 403624 307028 403676 307080
rect 74540 306348 74592 306400
rect 167644 306348 167696 306400
rect 98368 306280 98420 306332
rect 125784 306280 125836 306332
rect 143632 306280 143684 306332
rect 580264 306280 580316 306332
rect 3424 306212 3476 306264
rect 7564 306212 7616 306264
rect 121276 305668 121328 305720
rect 143632 305668 143684 305720
rect 97724 305600 97776 305652
rect 341616 305600 341668 305652
rect 125784 305124 125836 305176
rect 128544 305124 128596 305176
rect 85580 305056 85632 305108
rect 214656 305056 214708 305108
rect 114560 304988 114612 305040
rect 115296 304988 115348 305040
rect 245016 304988 245068 305040
rect 100668 304580 100720 304632
rect 104256 304580 104308 304632
rect 57520 304240 57572 304292
rect 126244 304240 126296 304292
rect 98644 303900 98696 303952
rect 180064 303900 180116 303952
rect 92664 303832 92716 303884
rect 210424 303832 210476 303884
rect 73252 303764 73304 303816
rect 228456 303764 228508 303816
rect 94044 303628 94096 303680
rect 95148 303628 95200 303680
rect 98000 303628 98052 303680
rect 98644 303628 98696 303680
rect 115940 303696 115992 303748
rect 116584 303696 116636 303748
rect 326344 303696 326396 303748
rect 416780 303628 416832 303680
rect 106832 303016 106884 303068
rect 132592 303016 132644 303068
rect 173164 303016 173216 303068
rect 75276 302948 75328 303000
rect 131212 302948 131264 303000
rect 353944 302948 353996 303000
rect 75184 302880 75236 302932
rect 331956 302880 332008 302932
rect 87512 302268 87564 302320
rect 240784 302268 240836 302320
rect 86316 302200 86368 302252
rect 276664 302200 276716 302252
rect 104992 301316 105044 301368
rect 106096 301316 106148 301368
rect 90272 301180 90324 301232
rect 220176 301180 220228 301232
rect 81532 301112 81584 301164
rect 251824 301112 251876 301164
rect 98644 301044 98696 301096
rect 283012 301044 283064 301096
rect 109040 300976 109092 301028
rect 298100 300976 298152 301028
rect 71780 300908 71832 300960
rect 306380 300908 306432 300960
rect 106096 300840 106148 300892
rect 450544 300840 450596 300892
rect 86224 300160 86276 300212
rect 132592 300160 132644 300212
rect 69020 300092 69072 300144
rect 342260 300092 342312 300144
rect 112444 299684 112496 299736
rect 227076 299684 227128 299736
rect 100852 299616 100904 299668
rect 256700 299616 256752 299668
rect 97356 299548 97408 299600
rect 279424 299548 279476 299600
rect 88984 299480 89036 299532
rect 303620 299480 303672 299532
rect 59176 298732 59228 298784
rect 124864 298732 124916 298784
rect 113824 298392 113876 298444
rect 169024 298392 169076 298444
rect 87420 298324 87472 298376
rect 211804 298324 211856 298376
rect 66076 298256 66128 298308
rect 203524 298256 203576 298308
rect 106740 298188 106792 298240
rect 269948 298188 270000 298240
rect 111248 298120 111300 298172
rect 278044 298120 278096 298172
rect 439504 298120 439556 298172
rect 580172 298120 580224 298172
rect 107568 297440 107620 297492
rect 127072 297440 127124 297492
rect 104164 297372 104216 297424
rect 125692 297372 125744 297424
rect 83556 296896 83608 296948
rect 133144 296896 133196 296948
rect 57888 296828 57940 296880
rect 100024 296828 100076 296880
rect 110604 296828 110656 296880
rect 249800 296828 249852 296880
rect 99656 296760 99708 296812
rect 258080 296760 258132 296812
rect 70676 296692 70728 296744
rect 300952 296692 301004 296744
rect 103428 295944 103480 295996
rect 323584 295944 323636 295996
rect 82912 295604 82964 295656
rect 135904 295604 135956 295656
rect 104256 295536 104308 295588
rect 104808 295536 104860 295588
rect 160744 295536 160796 295588
rect 91928 295468 91980 295520
rect 213276 295468 213328 295520
rect 102232 295400 102284 295452
rect 234620 295400 234672 295452
rect 117044 295332 117096 295384
rect 311900 295332 311952 295384
rect 72608 295264 72660 295316
rect 75276 295264 75328 295316
rect 54944 294720 54996 294772
rect 91284 294720 91336 294772
rect 70032 294652 70084 294704
rect 112444 294652 112496 294704
rect 77116 294584 77168 294636
rect 146484 294584 146536 294636
rect 428464 294584 428516 294636
rect 71320 294312 71372 294364
rect 72516 294312 72568 294364
rect 73160 294312 73212 294364
rect 73620 294312 73672 294364
rect 84292 294312 84344 294364
rect 85212 294312 85264 294364
rect 93952 294312 94004 294364
rect 94780 294312 94832 294364
rect 100024 294312 100076 294364
rect 101588 294312 101640 294364
rect 104900 294312 104952 294364
rect 105820 294312 105872 294364
rect 109960 294244 110012 294296
rect 122932 294244 122984 294296
rect 123668 294244 123720 294296
rect 102876 294176 102928 294228
rect 144184 294176 144236 294228
rect 97080 294108 97132 294160
rect 159456 294108 159508 294160
rect 65524 294040 65576 294092
rect 79048 294040 79100 294092
rect 108028 294040 108080 294092
rect 222844 294040 222896 294092
rect 34336 293972 34388 294024
rect 96436 293972 96488 294024
rect 113824 293972 113876 294024
rect 314660 293972 314712 294024
rect 2780 293156 2832 293208
rect 4804 293156 4856 293208
rect 118608 293020 118660 293072
rect 120080 293020 120132 293072
rect 93860 292816 93912 292868
rect 142804 292816 142856 292868
rect 69112 292748 69164 292800
rect 199384 292748 199436 292800
rect 75184 292680 75236 292732
rect 218704 292680 218756 292732
rect 51172 292612 51224 292664
rect 97080 292612 97132 292664
rect 103520 292612 103572 292664
rect 273904 292612 273956 292664
rect 11704 292544 11756 292596
rect 92572 292544 92624 292596
rect 93768 292544 93820 292596
rect 352564 292544 352616 292596
rect 51080 292476 51132 292528
rect 52184 292476 52236 292528
rect 65524 292476 65576 292528
rect 84292 291864 84344 291916
rect 4068 291796 4120 291848
rect 51080 291796 51132 291848
rect 104440 291864 104492 291916
rect 112812 291864 112864 291916
rect 119712 291864 119764 291916
rect 121552 291796 121604 291848
rect 124128 291796 124180 291848
rect 129648 291796 129700 291848
rect 273996 291388 274048 291440
rect 178776 291320 178828 291372
rect 119712 291252 119764 291304
rect 260840 291252 260892 291304
rect 22744 290436 22796 290488
rect 67640 290436 67692 290488
rect 121552 289892 121604 289944
rect 225604 289892 225656 289944
rect 121644 289824 121696 289876
rect 253940 289824 253992 289876
rect 121736 289144 121788 289196
rect 198096 289144 198148 289196
rect 121828 289076 121880 289128
rect 122012 289076 122064 289128
rect 452660 289076 452712 289128
rect 453304 289076 453356 289128
rect 50988 288396 51040 288448
rect 67640 288396 67692 288448
rect 121644 288396 121696 288448
rect 233884 288396 233936 288448
rect 66168 288328 66220 288380
rect 67732 288328 67784 288380
rect 121552 288328 121604 288380
rect 142436 288328 142488 288380
rect 143448 288328 143500 288380
rect 66076 288260 66128 288312
rect 68192 288260 68244 288312
rect 129740 287716 129792 287768
rect 282276 287716 282328 287768
rect 143448 287648 143500 287700
rect 360844 287648 360896 287700
rect 121460 286628 121512 286680
rect 121644 286628 121696 286680
rect 121460 286492 121512 286544
rect 125692 286492 125744 286544
rect 121552 286424 121604 286476
rect 128452 286424 128504 286476
rect 121644 286356 121696 286408
rect 130384 286356 130436 286408
rect 122288 286288 122340 286340
rect 287336 286288 287388 286340
rect 125692 284928 125744 284980
rect 305644 284928 305696 284980
rect 121460 284384 121512 284436
rect 293960 284384 294012 284436
rect 49424 284316 49476 284368
rect 67640 284316 67692 284368
rect 120908 284316 120960 284368
rect 414664 284316 414716 284368
rect 49608 284248 49660 284300
rect 67732 284248 67784 284300
rect 148324 283568 148376 283620
rect 365720 283568 365772 283620
rect 121460 282888 121512 282940
rect 272524 282888 272576 282940
rect 121460 281528 121512 281580
rect 224224 281528 224276 281580
rect 59176 280236 59228 280288
rect 67640 280236 67692 280288
rect 45376 280168 45428 280220
rect 67732 280168 67784 280220
rect 121460 280168 121512 280220
rect 251180 280168 251232 280220
rect 15844 279420 15896 279472
rect 42708 279420 42760 279472
rect 56416 279420 56468 279472
rect 128452 279420 128504 279472
rect 316684 279420 316736 279472
rect 121552 278808 121604 278860
rect 206376 278808 206428 278860
rect 56416 278740 56468 278792
rect 67640 278740 67692 278792
rect 121460 278740 121512 278792
rect 228364 278740 228416 278792
rect 126336 277992 126388 278044
rect 224316 277992 224368 278044
rect 121460 277448 121512 277500
rect 278136 277448 278188 277500
rect 48044 277380 48096 277432
rect 67640 277380 67692 277432
rect 121552 277380 121604 277432
rect 280896 277380 280948 277432
rect 60648 276088 60700 276140
rect 67640 276088 67692 276140
rect 121460 276088 121512 276140
rect 311992 276088 312044 276140
rect 53564 276020 53616 276072
rect 67732 276020 67784 276072
rect 121552 276020 121604 276072
rect 122288 276020 122340 276072
rect 418804 276020 418856 276072
rect 124128 275272 124180 275324
rect 419540 275272 419592 275324
rect 49516 274728 49568 274780
rect 67640 274728 67692 274780
rect 123576 274728 123628 274780
rect 129832 274728 129884 274780
rect 41236 274660 41288 274712
rect 67732 274660 67784 274712
rect 121460 274660 121512 274712
rect 234712 274660 234764 274712
rect 282184 273912 282236 273964
rect 308404 273912 308456 273964
rect 64604 273232 64656 273284
rect 67640 273232 67692 273284
rect 121460 273232 121512 273284
rect 200856 273232 200908 273284
rect 121460 272484 121512 272536
rect 123484 272484 123536 272536
rect 448520 272484 448572 272536
rect 65984 271940 66036 271992
rect 68100 271940 68152 271992
rect 64696 271872 64748 271924
rect 67640 271872 67692 271924
rect 121460 271872 121512 271924
rect 173900 271872 173952 271924
rect 59268 271124 59320 271176
rect 67640 271124 67692 271176
rect 123668 271124 123720 271176
rect 430948 271124 431000 271176
rect 57612 270512 57664 270564
rect 67732 270512 67784 270564
rect 121460 270512 121512 270564
rect 221464 270512 221516 270564
rect 55036 269152 55088 269204
rect 67732 269152 67784 269204
rect 121460 269152 121512 269204
rect 231952 269152 232004 269204
rect 39948 269084 40000 269136
rect 67640 269084 67692 269136
rect 121552 269084 121604 269136
rect 232136 269084 232188 269136
rect 39856 269016 39908 269068
rect 67732 269016 67784 269068
rect 121460 269016 121512 269068
rect 150440 269016 150492 269068
rect 22008 268336 22060 268388
rect 39856 268336 39908 268388
rect 150440 268336 150492 268388
rect 231216 268336 231268 268388
rect 121552 267724 121604 267776
rect 257344 267724 257396 267776
rect 41144 266976 41196 267028
rect 60188 266976 60240 267028
rect 60740 266500 60792 266552
rect 61384 266500 61436 266552
rect 67640 266500 67692 266552
rect 121644 266432 121696 266484
rect 255964 266432 256016 266484
rect 60188 266364 60240 266416
rect 60464 266364 60516 266416
rect 52276 266296 52328 266348
rect 60740 266296 60792 266348
rect 67732 266364 67784 266416
rect 121552 266364 121604 266416
rect 300860 266364 300912 266416
rect 62028 265616 62080 265668
rect 67640 265616 67692 265668
rect 121552 265004 121604 265056
rect 195336 265004 195388 265056
rect 52184 264936 52236 264988
rect 67732 264936 67784 264988
rect 121644 264936 121696 264988
rect 287152 264936 287204 264988
rect 48228 264868 48280 264920
rect 67640 264868 67692 264920
rect 7564 264188 7616 264240
rect 48228 264188 48280 264240
rect 130384 264188 130436 264240
rect 379520 264188 379572 264240
rect 121644 263576 121696 263628
rect 239036 263576 239088 263628
rect 121552 263508 121604 263560
rect 123024 263508 123076 263560
rect 124128 263508 124180 263560
rect 41328 262964 41380 263016
rect 53840 262964 53892 263016
rect 41328 262828 41380 262880
rect 66904 262828 66956 262880
rect 53840 262284 53892 262336
rect 54852 262284 54904 262336
rect 67732 262284 67784 262336
rect 121552 262284 121604 262336
rect 284300 262284 284352 262336
rect 50804 262216 50856 262268
rect 67640 262216 67692 262268
rect 134708 262216 134760 262268
rect 454040 262216 454092 262268
rect 121552 262148 121604 262200
rect 140780 262148 140832 262200
rect 140780 261468 140832 261520
rect 371884 261468 371936 261520
rect 48228 260856 48280 260908
rect 67732 260856 67784 260908
rect 121644 260856 121696 260908
rect 305000 260856 305052 260908
rect 56508 260788 56560 260840
rect 67640 260788 67692 260840
rect 121552 260788 121604 260840
rect 134708 260788 134760 260840
rect 124128 260108 124180 260160
rect 432144 260108 432196 260160
rect 121552 259496 121604 259548
rect 248420 259496 248472 259548
rect 63132 259428 63184 259480
rect 67640 259428 67692 259480
rect 137284 259428 137336 259480
rect 370504 259428 370556 259480
rect 121552 259360 121604 259412
rect 119988 259292 120040 259344
rect 121644 259292 121696 259344
rect 63316 258136 63368 258188
rect 67640 258136 67692 258188
rect 52276 258068 52328 258120
rect 67732 258068 67784 258120
rect 121736 258068 121788 258120
rect 280804 258068 280856 258120
rect 485044 258068 485096 258120
rect 580172 258068 580224 258120
rect 121460 257864 121512 257916
rect 121736 257864 121788 257916
rect 17224 257320 17276 257372
rect 35716 257320 35768 257372
rect 52460 257320 52512 257372
rect 162216 257320 162268 257372
rect 460940 257320 460992 257372
rect 121276 257048 121328 257100
rect 121644 257048 121696 257100
rect 61844 256776 61896 256828
rect 67640 256776 67692 256828
rect 52460 256708 52512 256760
rect 53472 256708 53524 256760
rect 67732 256708 67784 256760
rect 121460 256708 121512 256760
rect 227168 256708 227220 256760
rect 121644 255960 121696 256012
rect 315304 255960 315356 256012
rect 122840 255756 122892 255808
rect 125600 255756 125652 255808
rect 56324 255348 56376 255400
rect 67640 255348 67692 255400
rect 44088 255280 44140 255332
rect 67732 255280 67784 255332
rect 3148 255212 3200 255264
rect 33324 255212 33376 255264
rect 53748 255212 53800 255264
rect 67640 255212 67692 255264
rect 121460 255212 121512 255264
rect 131120 255212 131172 255264
rect 131488 255212 131540 255264
rect 33324 254532 33376 254584
rect 34244 254532 34296 254584
rect 60004 254532 60056 254584
rect 60556 254532 60608 254584
rect 67640 254532 67692 254584
rect 131488 254532 131540 254584
rect 330484 254532 330536 254584
rect 121644 253988 121696 254040
rect 250444 253988 250496 254040
rect 121460 253920 121512 253972
rect 259460 253920 259512 253972
rect 45468 253852 45520 253904
rect 47308 253852 47360 253904
rect 125600 253172 125652 253224
rect 356060 253172 356112 253224
rect 121644 252628 121696 252680
rect 220268 252628 220320 252680
rect 46940 252560 46992 252612
rect 47308 252560 47360 252612
rect 69020 252560 69072 252612
rect 121460 252560 121512 252612
rect 283104 252560 283156 252612
rect 178684 251880 178736 251932
rect 271236 251880 271288 251932
rect 121736 251812 121788 251864
rect 407764 251812 407816 251864
rect 54944 251200 54996 251252
rect 67640 251200 67692 251252
rect 121460 251200 121512 251252
rect 310520 251200 310572 251252
rect 169024 250520 169076 250572
rect 264336 250520 264388 250572
rect 135904 250452 135956 250504
rect 238852 250452 238904 250504
rect 53748 249840 53800 249892
rect 67732 249840 67784 249892
rect 120080 249840 120132 249892
rect 122840 249840 122892 249892
rect 50896 249772 50948 249824
rect 67640 249772 67692 249824
rect 121460 249772 121512 249824
rect 221556 249772 221608 249824
rect 121644 249364 121696 249416
rect 122748 249364 122800 249416
rect 124220 249364 124272 249416
rect 56508 249092 56560 249144
rect 68284 249092 68336 249144
rect 43444 249024 43496 249076
rect 59084 249024 59136 249076
rect 65892 249024 65944 249076
rect 68100 249024 68152 249076
rect 173164 249024 173216 249076
rect 400864 249024 400916 249076
rect 64512 248480 64564 248532
rect 67640 248480 67692 248532
rect 59084 248412 59136 248464
rect 67732 248412 67784 248464
rect 121460 248412 121512 248464
rect 196716 248412 196768 248464
rect 159456 247732 159508 247784
rect 367100 247732 367152 247784
rect 122840 247664 122892 247716
rect 375380 247664 375432 247716
rect 63224 247120 63276 247172
rect 67732 247120 67784 247172
rect 61936 247052 61988 247104
rect 67640 247052 67692 247104
rect 121460 247052 121512 247104
rect 240140 247052 240192 247104
rect 121460 246304 121512 246356
rect 431960 246304 432012 246356
rect 121552 245692 121604 245744
rect 234804 245692 234856 245744
rect 121460 245624 121512 245676
rect 242900 245624 242952 245676
rect 121552 244332 121604 244384
rect 258724 244332 258776 244384
rect 64788 244264 64840 244316
rect 67640 244264 67692 244316
rect 126244 244264 126296 244316
rect 579620 244264 579672 244316
rect 579988 244264 580040 244316
rect 121460 244196 121512 244248
rect 142252 244196 142304 244248
rect 143448 244196 143500 244248
rect 143448 243516 143500 243568
rect 311164 243516 311216 243568
rect 66168 242972 66220 243024
rect 67732 242972 67784 243024
rect 121552 242972 121604 243024
rect 279516 242972 279568 243024
rect 48136 242836 48188 242888
rect 58624 242836 58676 242888
rect 67640 242904 67692 242956
rect 124864 242904 124916 242956
rect 413284 242904 413336 242956
rect 121552 242836 121604 242888
rect 128360 242836 128412 242888
rect 121460 242768 121512 242820
rect 126244 242768 126296 242820
rect 122104 242156 122156 242208
rect 433524 242156 433576 242208
rect 66076 241476 66128 241528
rect 68192 241476 68244 241528
rect 121644 240728 121696 240780
rect 182180 240728 182232 240780
rect 121460 240116 121512 240168
rect 241796 240116 241848 240168
rect 3148 240048 3200 240100
rect 37188 240048 37240 240100
rect 69848 240048 69900 240100
rect 133972 240048 134024 240100
rect 134524 240048 134576 240100
rect 117688 239912 117740 239964
rect 124864 239912 124916 239964
rect 75920 239776 75972 239828
rect 77104 239776 77156 239828
rect 77300 239776 77352 239828
rect 78392 239776 78444 239828
rect 80060 239776 80112 239828
rect 80968 239776 81020 239828
rect 86960 239776 87012 239828
rect 88052 239776 88104 239828
rect 89720 239776 89772 239828
rect 90628 239776 90680 239828
rect 95240 239776 95292 239828
rect 96424 239776 96476 239828
rect 96620 239776 96672 239828
rect 97712 239776 97764 239828
rect 104900 239776 104952 239828
rect 106084 239776 106136 239828
rect 114560 239776 114612 239828
rect 115744 239776 115796 239828
rect 64788 239436 64840 239488
rect 78312 239436 78364 239488
rect 37188 239368 37240 239420
rect 88248 239368 88300 239420
rect 231216 239368 231268 239420
rect 411260 239368 411312 239420
rect 74632 239300 74684 239352
rect 75828 239300 75880 239352
rect 93952 239300 94004 239352
rect 95148 239300 95200 239352
rect 60004 238756 60056 238808
rect 111892 238756 111944 238808
rect 112536 238756 112588 238808
rect 116032 238756 116084 238808
rect 117044 238756 117096 238808
rect 127072 238756 127124 238808
rect 3424 238688 3476 238740
rect 86776 238688 86828 238740
rect 88248 238688 88300 238740
rect 103520 238688 103572 238740
rect 114468 238688 114520 238740
rect 132592 238688 132644 238740
rect 133788 238688 133840 238740
rect 57796 238620 57848 238672
rect 86132 238620 86184 238672
rect 57704 238552 57756 238604
rect 72608 238552 72660 238604
rect 86776 238280 86828 238332
rect 98828 238280 98880 238332
rect 105452 238280 105504 238332
rect 178684 238280 178736 238332
rect 100300 238212 100352 238264
rect 233240 238212 233292 238264
rect 69940 238144 69992 238196
rect 288532 238144 288584 238196
rect 70676 238076 70728 238128
rect 313280 238076 313332 238128
rect 72608 238008 72660 238060
rect 86316 238008 86368 238060
rect 98828 238008 98880 238060
rect 99196 238008 99248 238060
rect 128544 238008 128596 238060
rect 133788 238008 133840 238060
rect 434720 238008 434772 238060
rect 103520 237464 103572 237516
rect 104164 237464 104216 237516
rect 85488 237396 85540 237448
rect 86224 237396 86276 237448
rect 102876 237396 102928 237448
rect 105544 237396 105596 237448
rect 69204 237328 69256 237380
rect 138020 237328 138072 237380
rect 52368 237260 52420 237312
rect 81624 237260 81676 237312
rect 99288 237260 99340 237312
rect 123576 237260 123628 237312
rect 66168 236716 66220 236768
rect 276756 236716 276808 236768
rect 138020 236648 138072 236700
rect 385040 236648 385092 236700
rect 81624 235968 81676 236020
rect 82084 235968 82136 236020
rect 110604 235900 110656 235952
rect 111064 235900 111116 235952
rect 136640 235900 136692 235952
rect 61936 235356 61988 235408
rect 245660 235356 245712 235408
rect 231124 235288 231176 235340
rect 446404 235288 446456 235340
rect 57612 235220 57664 235272
rect 290096 235220 290148 235272
rect 46848 234540 46900 234592
rect 118976 234540 119028 234592
rect 53656 234472 53708 234524
rect 91744 234472 91796 234524
rect 118976 234132 119028 234184
rect 119344 234132 119396 234184
rect 108028 233860 108080 233912
rect 284392 233860 284444 233912
rect 84200 233792 84252 233844
rect 84292 233588 84344 233640
rect 55128 233180 55180 233232
rect 109684 233180 109736 233232
rect 52184 232704 52236 232756
rect 157984 232704 158036 232756
rect 78312 232636 78364 232688
rect 222936 232636 222988 232688
rect 69112 232568 69164 232620
rect 281724 232568 281776 232620
rect 107384 232500 107436 232552
rect 411904 232500 411956 232552
rect 74448 231820 74500 231872
rect 75184 231820 75236 231872
rect 93768 231820 93820 231872
rect 94504 231820 94556 231872
rect 349068 231820 349120 231872
rect 580172 231820 580224 231872
rect 101496 231140 101548 231192
rect 229284 231140 229336 231192
rect 134524 231072 134576 231124
rect 443000 231072 443052 231124
rect 82912 230392 82964 230444
rect 83464 230392 83516 230444
rect 149060 230392 149112 230444
rect 89260 230324 89312 230376
rect 126980 230324 127032 230376
rect 127440 230324 127492 230376
rect 67456 229848 67508 229900
rect 230480 229848 230532 229900
rect 127440 229780 127492 229832
rect 173164 229780 173216 229832
rect 180064 229780 180116 229832
rect 382280 229780 382332 229832
rect 48228 229712 48280 229764
rect 276848 229712 276900 229764
rect 111892 228420 111944 228472
rect 378140 228420 378192 228472
rect 98644 228352 98696 228404
rect 418896 228352 418948 228404
rect 94044 226992 94096 227044
rect 236000 226992 236052 227044
rect 60556 225700 60608 225752
rect 164884 225700 164936 225752
rect 56324 225632 56376 225684
rect 252560 225632 252612 225684
rect 74724 225564 74776 225616
rect 303712 225564 303764 225616
rect 91744 224884 91796 224936
rect 438952 224884 439004 224936
rect 438952 224476 439004 224528
rect 439504 224476 439556 224528
rect 59176 224272 59228 224324
rect 187056 224272 187108 224324
rect 65984 224204 66036 224256
rect 230572 224204 230624 224256
rect 59084 222844 59136 222896
rect 417424 222844 417476 222896
rect 82912 222640 82964 222692
rect 83464 222640 83516 222692
rect 4804 222164 4856 222216
rect 82912 222164 82964 222216
rect 118240 222096 118292 222148
rect 146300 222096 146352 222148
rect 146760 222096 146812 222148
rect 282276 221552 282328 221604
rect 299480 221552 299532 221604
rect 146760 221484 146812 221536
rect 301504 221484 301556 221536
rect 86316 221416 86368 221468
rect 440240 221416 440292 221468
rect 233884 220124 233936 220176
rect 309140 220124 309192 220176
rect 48044 220056 48096 220108
rect 260196 220056 260248 220108
rect 89812 218764 89864 218816
rect 233424 218764 233476 218816
rect 61384 218696 61436 218748
rect 363604 218696 363656 218748
rect 446404 218696 446456 218748
rect 580172 218696 580224 218748
rect 74632 217404 74684 217456
rect 147680 217404 147732 217456
rect 41236 217336 41288 217388
rect 275284 217336 275336 217388
rect 104164 217268 104216 217320
rect 400220 217268 400272 217320
rect 54852 215908 54904 215960
rect 414020 215908 414072 215960
rect 81532 215228 81584 215280
rect 151820 215228 151872 215280
rect 153108 215228 153160 215280
rect 3332 214616 3384 214668
rect 7564 214616 7616 214668
rect 209044 214616 209096 214668
rect 153108 214548 153160 214600
rect 407120 214548 407172 214600
rect 69020 213188 69072 213240
rect 391940 213188 391992 213240
rect 58624 211760 58676 211812
rect 401600 211760 401652 211812
rect 45376 210400 45428 210452
rect 307760 210400 307812 210452
rect 109684 209788 109736 209840
rect 389180 209788 389232 209840
rect 113180 209108 113232 209160
rect 302240 209108 302292 209160
rect 50896 209040 50948 209092
rect 247040 209040 247092 209092
rect 111800 207680 111852 207732
rect 249892 207680 249944 207732
rect 56416 207612 56468 207664
rect 387800 207612 387852 207664
rect 100760 206320 100812 206372
rect 225696 206320 225748 206372
rect 78772 206252 78824 206304
rect 285680 206252 285732 206304
rect 450544 206252 450596 206304
rect 580172 206252 580224 206304
rect 82820 205572 82872 205624
rect 133880 205572 133932 205624
rect 135168 205572 135220 205624
rect 122104 205096 122156 205148
rect 310612 205096 310664 205148
rect 55036 205028 55088 205080
rect 248512 205028 248564 205080
rect 92572 204960 92624 205012
rect 288440 204960 288492 205012
rect 135168 204892 135220 204944
rect 429476 204892 429528 204944
rect 114468 203804 114520 203856
rect 166356 203804 166408 203856
rect 86960 203736 87012 203788
rect 251272 203736 251324 203788
rect 114560 203668 114612 203720
rect 283196 203668 283248 203720
rect 63132 203600 63184 203652
rect 299572 203600 299624 203652
rect 3332 203532 3384 203584
rect 120080 203532 120132 203584
rect 164884 203532 164936 203584
rect 439136 203532 439188 203584
rect 157984 202240 158036 202292
rect 296720 202240 296772 202292
rect 86224 202172 86276 202224
rect 242992 202172 243044 202224
rect 80152 202104 80204 202156
rect 278228 202104 278280 202156
rect 228456 201084 228508 201136
rect 298192 201084 298244 201136
rect 96712 201016 96764 201068
rect 241612 201016 241664 201068
rect 104900 200948 104952 201000
rect 272616 200948 272668 201000
rect 49516 200880 49568 200932
rect 237380 200880 237432 200932
rect 67364 200812 67416 200864
rect 307944 200812 307996 200864
rect 99196 200744 99248 200796
rect 443092 200744 443144 200796
rect 144184 199520 144236 199572
rect 223028 199520 223080 199572
rect 116032 199452 116084 199504
rect 428096 199452 428148 199504
rect 82084 199384 82136 199436
rect 432236 199384 432288 199436
rect 50804 198092 50856 198144
rect 217324 198092 217376 198144
rect 280896 198092 280948 198144
rect 301044 198092 301096 198144
rect 93952 198024 94004 198076
rect 305092 198024 305144 198076
rect 61844 197956 61896 198008
rect 302332 197956 302384 198008
rect 110420 196800 110472 196852
rect 233332 196800 233384 196852
rect 105544 196732 105596 196784
rect 240232 196732 240284 196784
rect 65892 196664 65944 196716
rect 295432 196664 295484 196716
rect 83464 196596 83516 196648
rect 369860 196596 369912 196648
rect 92480 195440 92532 195492
rect 211896 195440 211948 195492
rect 222844 195440 222896 195492
rect 294052 195440 294104 195492
rect 209136 195372 209188 195424
rect 437572 195372 437624 195424
rect 49424 195304 49476 195356
rect 306472 195304 306524 195356
rect 59268 195236 59320 195288
rect 436100 195236 436152 195288
rect 89720 194148 89772 194200
rect 252652 194148 252704 194200
rect 64604 194080 64656 194132
rect 230664 194080 230716 194132
rect 93860 194012 93912 194064
rect 309232 194012 309284 194064
rect 60648 193944 60700 193996
rect 278320 193944 278372 193996
rect 99288 193876 99340 193928
rect 329104 193876 329156 193928
rect 155224 193808 155276 193860
rect 447140 193808 447192 193860
rect 53564 192584 53616 192636
rect 221648 192584 221700 192636
rect 160744 192516 160796 192568
rect 434812 192516 434864 192568
rect 60464 192448 60516 192500
rect 451280 192448 451332 192500
rect 475384 192448 475436 192500
rect 579620 192448 579672 192500
rect 203524 191360 203576 191412
rect 244280 191360 244332 191412
rect 244924 191360 244976 191412
rect 337476 191360 337528 191412
rect 102140 191292 102192 191344
rect 292672 191292 292724 191344
rect 66076 191224 66128 191276
rect 256792 191224 256844 191276
rect 50988 191156 51040 191208
rect 245752 191156 245804 191208
rect 88340 191088 88392 191140
rect 285956 191088 286008 191140
rect 108948 190476 109000 190528
rect 214748 190476 214800 190528
rect 77300 189864 77352 189916
rect 229192 189864 229244 189916
rect 73252 189796 73304 189848
rect 285864 189796 285916 189848
rect 169024 189728 169076 189780
rect 436376 189728 436428 189780
rect 106188 189184 106240 189236
rect 169116 189184 169168 189236
rect 104808 189116 104860 189168
rect 173256 189116 173308 189168
rect 3516 189048 3568 189100
rect 4068 189048 4120 189100
rect 441712 189048 441764 189100
rect 3424 188980 3476 189032
rect 11704 188980 11756 189032
rect 279516 188640 279568 188692
rect 292764 188640 292816 188692
rect 278136 188572 278188 188624
rect 306564 188572 306616 188624
rect 99380 188504 99432 188556
rect 280344 188504 280396 188556
rect 118700 188436 118752 188488
rect 309324 188436 309376 188488
rect 71780 188368 71832 188420
rect 280160 188368 280212 188420
rect 54944 188300 54996 188352
rect 305184 188300 305236 188352
rect 103428 187756 103480 187808
rect 171784 187756 171836 187808
rect 131028 187688 131080 187740
rect 209136 187688 209188 187740
rect 146944 187076 146996 187128
rect 175924 187076 175976 187128
rect 95240 187008 95292 187060
rect 274088 187008 274140 187060
rect 73160 186940 73212 186992
rect 291292 186940 291344 186992
rect 348976 186940 349028 186992
rect 580908 186940 580960 186992
rect 153844 185852 153896 185904
rect 289912 185852 289964 185904
rect 84200 185784 84252 185836
rect 280252 185784 280304 185836
rect 52276 185716 52328 185768
rect 251364 185716 251416 185768
rect 264244 185716 264296 185768
rect 448612 185716 448664 185768
rect 80060 185648 80112 185700
rect 310704 185648 310756 185700
rect 39948 185580 40000 185632
rect 295524 185580 295576 185632
rect 350816 185580 350868 185632
rect 381544 185580 381596 185632
rect 395344 185580 395396 185632
rect 425796 185580 425848 185632
rect 100668 184900 100720 184952
rect 169208 184900 169260 184952
rect 151084 184424 151136 184476
rect 174544 184424 174596 184476
rect 210424 184424 210476 184476
rect 243084 184424 243136 184476
rect 103704 184356 103756 184408
rect 284484 184356 284536 184408
rect 63224 184288 63276 184340
rect 247132 184288 247184 184340
rect 271144 184288 271196 184340
rect 445852 184288 445904 184340
rect 75920 184220 75972 184272
rect 285772 184220 285824 184272
rect 44088 184152 44140 184204
rect 291200 184152 291252 184204
rect 358084 184152 358136 184204
rect 374644 184152 374696 184204
rect 129648 183540 129700 183592
rect 209320 183540 209372 183592
rect 187056 183064 187108 183116
rect 244372 183064 244424 183116
rect 255964 183064 256016 183116
rect 296904 183064 296956 183116
rect 142804 182996 142856 183048
rect 238760 182996 238812 183048
rect 265624 182996 265676 183048
rect 316868 182996 316920 183048
rect 411904 182996 411956 183048
rect 443184 182996 443236 183048
rect 115940 182928 115992 182980
rect 241704 182928 241756 182980
rect 262956 182928 263008 182980
rect 319444 182928 319496 182980
rect 400864 182928 400916 182980
rect 449900 182928 449952 182980
rect 64696 182860 64748 182912
rect 230756 182860 230808 182912
rect 269764 182860 269816 182912
rect 434904 182860 434956 182912
rect 107660 182792 107712 182844
rect 307852 182792 307904 182844
rect 360844 182792 360896 182844
rect 444472 182792 444524 182844
rect 119528 182180 119580 182232
rect 211804 182180 211856 182232
rect 220268 181772 220320 181824
rect 237472 181772 237524 181824
rect 269856 181772 269908 181824
rect 314108 181772 314160 181824
rect 162124 181704 162176 181756
rect 200764 181704 200816 181756
rect 200856 181704 200908 181756
rect 240324 181704 240376 181756
rect 251824 181704 251876 181756
rect 296812 181704 296864 181756
rect 199384 181636 199436 181688
rect 248604 181636 248656 181688
rect 249064 181636 249116 181688
rect 300216 181636 300268 181688
rect 167644 181568 167696 181620
rect 244464 181568 244516 181620
rect 264336 181568 264388 181620
rect 323676 181568 323728 181620
rect 96620 181500 96672 181552
rect 202236 181500 202288 181552
rect 214656 181500 214708 181552
rect 237564 181500 237616 181552
rect 245016 181500 245068 181552
rect 424416 181500 424468 181552
rect 53748 181432 53800 181484
rect 298284 181432 298336 181484
rect 361304 181432 361356 181484
rect 405740 181432 405792 181484
rect 132408 180956 132460 181008
rect 164884 180956 164936 181008
rect 122012 180888 122064 180940
rect 167828 180888 167880 180940
rect 116952 180820 117004 180872
rect 167736 180820 167788 180872
rect 223028 180412 223080 180464
rect 236184 180412 236236 180464
rect 272524 180412 272576 180464
rect 288624 180412 288676 180464
rect 222936 180344 222988 180396
rect 236092 180344 236144 180396
rect 273904 180344 273956 180396
rect 302424 180344 302476 180396
rect 225604 180276 225656 180328
rect 245844 180276 245896 180328
rect 273996 180276 274048 180328
rect 303804 180276 303856 180328
rect 414664 180276 414716 180328
rect 444380 180276 444432 180328
rect 220176 180208 220228 180260
rect 247224 180208 247276 180260
rect 258724 180208 258776 180260
rect 294144 180208 294196 180260
rect 363788 180208 363840 180260
rect 376760 180208 376812 180260
rect 407764 180208 407816 180260
rect 439044 180208 439096 180260
rect 159364 180140 159416 180192
rect 192484 180140 192536 180192
rect 198096 180140 198148 180192
rect 347320 180140 347372 180192
rect 359464 180140 359516 180192
rect 437480 180140 437532 180192
rect 173164 180072 173216 180124
rect 438860 180072 438912 180124
rect 133144 179664 133196 179716
rect 164424 179664 164476 179716
rect 121000 179596 121052 179648
rect 166540 179596 166592 179648
rect 115848 179528 115900 179580
rect 166448 179528 166500 179580
rect 97356 179460 97408 179512
rect 173348 179460 173400 179512
rect 112260 179392 112312 179444
rect 198188 179392 198240 179444
rect 276756 178984 276808 179036
rect 290004 178984 290056 179036
rect 217324 178916 217376 178968
rect 238944 178916 238996 178968
rect 272616 178916 272668 178968
rect 287244 178916 287296 178968
rect 178776 178848 178828 178900
rect 224960 178848 225012 178900
rect 257344 178848 257396 178900
rect 295340 178848 295392 178900
rect 418804 178848 418856 178900
rect 436192 178848 436244 178900
rect 214564 178780 214616 178832
rect 312544 178780 312596 178832
rect 399484 178780 399536 178832
rect 429384 178780 429436 178832
rect 64512 178712 64564 178764
rect 254032 178712 254084 178764
rect 271236 178712 271288 178764
rect 333336 178712 333388 178764
rect 358176 178712 358228 178764
rect 433432 178712 433484 178764
rect 220084 178644 220136 178696
rect 430580 178644 430632 178696
rect 148232 178304 148284 178356
rect 169024 178304 169076 178356
rect 114376 178236 114428 178288
rect 167920 178236 167972 178288
rect 109776 178168 109828 178220
rect 170496 178168 170548 178220
rect 127072 178100 127124 178152
rect 211988 178100 212040 178152
rect 118424 177964 118476 178016
rect 214656 178032 214708 178084
rect 468484 178032 468536 178084
rect 580172 178032 580224 178084
rect 278044 177624 278096 177676
rect 288716 177624 288768 177676
rect 221648 177556 221700 177608
rect 229560 177556 229612 177608
rect 275284 177556 275336 177608
rect 294236 177556 294288 177608
rect 417424 177556 417476 177608
rect 426900 177556 426952 177608
rect 227168 177488 227220 177540
rect 234896 177488 234948 177540
rect 250444 177488 250496 177540
rect 292580 177488 292632 177540
rect 413284 177488 413336 177540
rect 434996 177488 435048 177540
rect 211896 177420 211948 177472
rect 237656 177420 237708 177472
rect 268384 177420 268436 177472
rect 325148 177420 325200 177472
rect 352564 177420 352616 177472
rect 397460 177420 397512 177472
rect 418896 177420 418948 177472
rect 441620 177420 441672 177472
rect 206376 177352 206428 177404
rect 279424 177352 279476 177404
rect 363604 177352 363656 177404
rect 422300 177352 422352 177404
rect 166356 177284 166408 177336
rect 353300 177284 353352 177336
rect 370504 177284 370556 177336
rect 437664 177284 437716 177336
rect 134432 176944 134484 176996
rect 165252 176944 165304 176996
rect 125784 176876 125836 176928
rect 166632 176876 166684 176928
rect 111064 176808 111116 176860
rect 124496 176808 124548 176860
rect 170588 176808 170640 176860
rect 14464 176740 14516 176792
rect 109408 176740 109460 176792
rect 110696 176740 110748 176792
rect 214564 176740 214616 176792
rect 102048 176672 102100 176724
rect 213368 176672 213420 176724
rect 240784 176672 240836 176724
rect 241520 176672 241572 176724
rect 403624 176672 403676 176724
rect 404820 176672 404872 176724
rect 135720 176604 135772 176656
rect 213920 176604 213972 176656
rect 228364 176604 228416 176656
rect 229468 176604 229520 176656
rect 260196 176604 260248 176656
rect 279516 176604 279568 176656
rect 158904 176196 158956 176248
rect 167644 176196 167696 176248
rect 123116 176128 123168 176180
rect 166264 176128 166316 176180
rect 274088 176128 274140 176180
rect 281540 176128 281592 176180
rect 128176 176060 128228 176112
rect 214104 176060 214156 176112
rect 225696 176060 225748 176112
rect 232044 176060 232096 176112
rect 278228 176060 278280 176112
rect 287060 176060 287112 176112
rect 421564 176060 421616 176112
rect 430672 176060 430724 176112
rect 25504 175992 25556 176044
rect 109684 175992 109736 176044
rect 113180 175992 113232 176044
rect 209228 175992 209280 176044
rect 221464 175992 221516 176044
rect 229376 175992 229428 176044
rect 279608 175992 279660 176044
rect 289820 175992 289872 176044
rect 371884 175992 371936 176044
rect 440332 175992 440384 176044
rect 98368 175924 98420 175976
rect 206376 175924 206428 175976
rect 224224 175924 224276 175976
rect 240416 175924 240468 175976
rect 276848 175924 276900 175976
rect 291384 175924 291436 175976
rect 353944 175924 353996 175976
rect 436284 175924 436336 175976
rect 425796 175856 425848 175908
rect 429292 175856 429344 175908
rect 224960 175788 225012 175840
rect 227720 175788 227772 175840
rect 333244 175244 333296 175296
rect 165252 175176 165304 175228
rect 213920 175176 213972 175228
rect 427820 175176 427872 175228
rect 164424 175108 164476 175160
rect 214012 175108 214064 175160
rect 256056 174020 256108 174072
rect 265348 174020 265400 174072
rect 250444 173952 250496 174004
rect 265900 173952 265952 174004
rect 244924 173884 244976 173936
rect 265808 173884 265860 173936
rect 322296 173884 322348 173936
rect 347504 173884 347556 173936
rect 164884 173816 164936 173868
rect 213920 173816 213972 173868
rect 231400 173816 231452 173868
rect 238760 173816 238812 173868
rect 209136 173748 209188 173800
rect 214012 173748 214064 173800
rect 260104 172660 260156 172712
rect 265348 172660 265400 172712
rect 243820 172592 243872 172644
rect 265808 172592 265860 172644
rect 239404 172524 239456 172576
rect 265256 172524 265308 172576
rect 320916 172524 320968 172576
rect 347504 172524 347556 172576
rect 430580 172524 430632 172576
rect 433616 172524 433668 172576
rect 209320 172456 209372 172508
rect 213920 172456 213972 172508
rect 240140 172456 240192 172508
rect 241520 172456 241572 172508
rect 231676 172388 231728 172440
rect 240048 172388 240100 172440
rect 231768 172320 231820 172372
rect 240324 172320 240376 172372
rect 246396 171776 246448 171828
rect 265992 171776 266044 171828
rect 167092 171300 167144 171352
rect 169300 171300 169352 171352
rect 258724 171300 258776 171352
rect 265164 171300 265216 171352
rect 242256 171096 242308 171148
rect 265072 171096 265124 171148
rect 325056 171096 325108 171148
rect 347504 171096 347556 171148
rect 166632 171028 166684 171080
rect 213920 171028 213972 171080
rect 231768 171028 231820 171080
rect 245660 171028 245712 171080
rect 282736 171028 282788 171080
rect 291292 171028 291344 171080
rect 211988 170960 212040 171012
rect 214012 170960 214064 171012
rect 282828 170960 282880 171012
rect 289820 170960 289872 171012
rect 231676 170892 231728 170944
rect 237564 170892 237616 170944
rect 231768 170144 231820 170196
rect 237380 170144 237432 170196
rect 251916 169872 251968 169924
rect 265256 169872 265308 169924
rect 250536 169804 250588 169856
rect 265440 169804 265492 169856
rect 249708 169736 249760 169788
rect 265624 169736 265676 169788
rect 166264 169668 166316 169720
rect 214012 169668 214064 169720
rect 231676 169668 231728 169720
rect 241612 169668 241664 169720
rect 170588 169600 170640 169652
rect 213920 169600 213972 169652
rect 231400 169600 231452 169652
rect 240140 169600 240192 169652
rect 231768 169532 231820 169584
rect 240232 169532 240284 169584
rect 259000 169464 259052 169516
rect 265348 169464 265400 169516
rect 281908 168852 281960 168904
rect 287060 168852 287112 168904
rect 240968 168444 241020 168496
rect 240876 168376 240928 168428
rect 243084 168376 243136 168428
rect 246672 168444 246724 168496
rect 265348 168444 265400 168496
rect 265900 168376 265952 168428
rect 307024 168376 307076 168428
rect 347044 168376 347096 168428
rect 166540 168308 166592 168360
rect 214012 168308 214064 168360
rect 231768 168308 231820 168360
rect 238852 168308 238904 168360
rect 281908 168308 281960 168360
rect 295432 168308 295484 168360
rect 167828 168240 167880 168292
rect 213920 168240 213972 168292
rect 282368 168240 282420 168292
rect 290004 168240 290056 168292
rect 231216 167968 231268 168020
rect 237472 167968 237524 168020
rect 243728 167628 243780 167680
rect 265808 167628 265860 167680
rect 249064 167152 249116 167204
rect 265256 167152 265308 167204
rect 242164 167084 242216 167136
rect 249708 167084 249760 167136
rect 238024 167016 238076 167068
rect 265532 167016 265584 167068
rect 327816 167016 327868 167068
rect 347504 167016 347556 167068
rect 167736 166948 167788 167000
rect 213920 166948 213972 167000
rect 231768 166948 231820 167000
rect 241796 166948 241848 167000
rect 282092 166948 282144 167000
rect 295524 166948 295576 167000
rect 211804 166880 211856 166932
rect 214104 166880 214156 166932
rect 231492 166880 231544 166932
rect 238944 166880 238996 166932
rect 429108 166812 429160 166864
rect 433432 166812 433484 166864
rect 230572 166268 230624 166320
rect 230940 166268 230992 166320
rect 231584 166268 231636 166320
rect 237656 166268 237708 166320
rect 280804 166268 280856 166320
rect 281632 166268 281684 166320
rect 314016 166268 314068 166320
rect 346676 166268 346728 166320
rect 346860 166268 346912 166320
rect 263140 165724 263192 165776
rect 265808 165724 265860 165776
rect 253204 165656 253256 165708
rect 265624 165656 265676 165708
rect 238392 165588 238444 165640
rect 265900 165588 265952 165640
rect 166448 165520 166500 165572
rect 213920 165520 213972 165572
rect 231032 165520 231084 165572
rect 249800 165520 249852 165572
rect 282092 165520 282144 165572
rect 292672 165520 292724 165572
rect 167920 165452 167972 165504
rect 214012 165452 214064 165504
rect 231124 165452 231176 165504
rect 233424 165452 233476 165504
rect 247868 164840 247920 164892
rect 265440 164840 265492 164892
rect 327724 164840 327776 164892
rect 339500 164840 339552 164892
rect 467104 164840 467156 164892
rect 580172 164840 580224 164892
rect 282368 164228 282420 164280
rect 288532 164228 288584 164280
rect 339500 164228 339552 164280
rect 347504 164228 347556 164280
rect 198188 164160 198240 164212
rect 214012 164160 214064 164212
rect 231768 164160 231820 164212
rect 244464 164160 244516 164212
rect 282184 164160 282236 164212
rect 299572 164160 299624 164212
rect 430580 164160 430632 164212
rect 436376 164160 436428 164212
rect 436652 164160 436704 164212
rect 209228 164092 209280 164144
rect 213920 164092 213972 164144
rect 231676 164092 231728 164144
rect 244280 164092 244332 164144
rect 282828 164092 282880 164144
rect 291384 164092 291436 164144
rect 231492 164024 231544 164076
rect 239036 164024 239088 164076
rect 229928 163684 229980 163736
rect 234896 163684 234948 163736
rect 229744 163480 229796 163532
rect 242900 163480 242952 163532
rect 245016 163480 245068 163532
rect 265164 163480 265216 163532
rect 336188 163480 336240 163532
rect 345020 163480 345072 163532
rect 346676 163480 346728 163532
rect 436652 163480 436704 163532
rect 471244 163480 471296 163532
rect 240140 163140 240192 163192
rect 245752 163140 245804 163192
rect 260196 162936 260248 162988
rect 265624 162936 265676 162988
rect 234160 162868 234212 162920
rect 265532 162868 265584 162920
rect 170496 162800 170548 162852
rect 213920 162800 213972 162852
rect 282092 162800 282144 162852
rect 298100 162800 298152 162852
rect 430580 162800 430632 162852
rect 434996 162800 435048 162852
rect 436008 162800 436060 162852
rect 231768 162732 231820 162784
rect 244372 162732 244424 162784
rect 282828 162732 282880 162784
rect 292764 162732 292816 162784
rect 430580 162188 430632 162240
rect 439136 162188 439188 162240
rect 436008 162120 436060 162172
rect 464344 162120 464396 162172
rect 234068 161780 234120 161832
rect 240416 161780 240468 161832
rect 253296 161576 253348 161628
rect 264520 161576 264572 161628
rect 246304 161508 246356 161560
rect 265716 161508 265768 161560
rect 238116 161440 238168 161492
rect 265808 161440 265860 161492
rect 231768 161372 231820 161424
rect 241704 161372 241756 161424
rect 282736 161372 282788 161424
rect 293960 161372 294012 161424
rect 343640 161372 343692 161424
rect 347504 161372 347556 161424
rect 430580 161372 430632 161424
rect 444472 161372 444524 161424
rect 231308 161304 231360 161356
rect 238852 161304 238904 161356
rect 169300 160692 169352 160744
rect 214564 160692 214616 160744
rect 318156 160692 318208 160744
rect 343640 160692 343692 160744
rect 282828 160420 282880 160472
rect 288716 160420 288768 160472
rect 257344 160216 257396 160268
rect 265624 160216 265676 160268
rect 240784 160148 240836 160200
rect 265348 160148 265400 160200
rect 239496 160080 239548 160132
rect 265808 160080 265860 160132
rect 444472 160080 444524 160132
rect 447784 160080 447836 160132
rect 169116 160012 169168 160064
rect 213920 160012 213972 160064
rect 231768 160012 231820 160064
rect 245844 160012 245896 160064
rect 282092 160012 282144 160064
rect 313280 160012 313332 160064
rect 430580 160012 430632 160064
rect 454040 160012 454092 160064
rect 467104 160012 467156 160064
rect 173256 159944 173308 159996
rect 214012 159944 214064 159996
rect 231032 159944 231084 159996
rect 240140 159944 240192 159996
rect 231584 159876 231636 159928
rect 234068 159876 234120 159928
rect 250628 159332 250680 159384
rect 265992 159332 266044 159384
rect 316776 159332 316828 159384
rect 340880 159332 340932 159384
rect 347504 159332 347556 159384
rect 245200 158788 245252 158840
rect 265808 158788 265860 158840
rect 239680 158720 239732 158772
rect 265716 158720 265768 158772
rect 171784 158652 171836 158704
rect 213920 158652 213972 158704
rect 231768 158652 231820 158704
rect 252560 158652 252612 158704
rect 282736 158652 282788 158704
rect 302424 158652 302476 158704
rect 430580 158652 430632 158704
rect 450544 158652 450596 158704
rect 231216 158584 231268 158636
rect 240876 158584 240928 158636
rect 282828 158584 282880 158636
rect 300860 158584 300912 158636
rect 324964 157972 325016 158024
rect 342352 157972 342404 158024
rect 261576 157496 261628 157548
rect 265900 157496 265952 157548
rect 245292 157428 245344 157480
rect 265716 157428 265768 157480
rect 342352 157428 342404 157480
rect 347504 157428 347556 157480
rect 237380 157360 237432 157412
rect 265624 157360 265676 157412
rect 169208 157292 169260 157344
rect 213920 157292 213972 157344
rect 231768 157292 231820 157344
rect 256700 157292 256752 157344
rect 282092 157292 282144 157344
rect 303804 157292 303856 157344
rect 430580 157292 430632 157344
rect 475384 157292 475436 157344
rect 231124 157224 231176 157276
rect 248420 157224 248472 157276
rect 231584 156748 231636 156800
rect 234712 156748 234764 156800
rect 232688 156680 232740 156732
rect 251364 156680 251416 156732
rect 242440 156612 242492 156664
rect 265164 156612 265216 156664
rect 336096 156068 336148 156120
rect 343640 156068 343692 156120
rect 347044 156068 347096 156120
rect 252100 156000 252152 156052
rect 265532 156000 265584 156052
rect 240876 155932 240928 155984
rect 265900 155932 265952 155984
rect 281540 155932 281592 155984
rect 283104 155932 283156 155984
rect 173348 155864 173400 155916
rect 214012 155864 214064 155916
rect 231492 155864 231544 155916
rect 247224 155864 247276 155916
rect 282368 155864 282420 155916
rect 307944 155864 307996 155916
rect 430856 155864 430908 155916
rect 482284 155864 482336 155916
rect 206376 155796 206428 155848
rect 213920 155796 213972 155848
rect 231768 155796 231820 155848
rect 242992 155796 243044 155848
rect 282092 155796 282144 155848
rect 306564 155796 306616 155848
rect 430580 155796 430632 155848
rect 438952 155796 439004 155848
rect 256332 155252 256384 155304
rect 265348 155252 265400 155304
rect 238208 155184 238260 155236
rect 265992 155184 266044 155236
rect 241152 154572 241204 154624
rect 265808 154572 265860 154624
rect 231768 154504 231820 154556
rect 251272 154504 251324 154556
rect 282460 154504 282512 154556
rect 310704 154504 310756 154556
rect 430580 154504 430632 154556
rect 479524 154504 479576 154556
rect 231676 154436 231728 154488
rect 248512 154436 248564 154488
rect 281908 154164 281960 154216
rect 285956 154164 286008 154216
rect 252192 153824 252244 153876
rect 265992 153824 266044 153876
rect 309784 153824 309836 153876
rect 345020 153824 345072 153876
rect 346676 153824 346728 153876
rect 231124 153756 231176 153808
rect 238392 153756 238444 153808
rect 198096 153280 198148 153332
rect 214012 153280 214064 153332
rect 238300 153280 238352 153332
rect 265808 153280 265860 153332
rect 187056 153212 187108 153264
rect 213920 153212 213972 153264
rect 236736 153212 236788 153264
rect 265900 153212 265952 153264
rect 231768 153144 231820 153196
rect 260840 153144 260892 153196
rect 430580 153144 430632 153196
rect 457444 153144 457496 153196
rect 230480 152532 230532 152584
rect 233240 152532 233292 152584
rect 234160 152464 234212 152516
rect 265716 152464 265768 152516
rect 211804 152396 211856 152448
rect 213920 152396 213972 152448
rect 345112 152056 345164 152108
rect 346584 152056 346636 152108
rect 189724 151852 189776 151904
rect 214012 151852 214064 151904
rect 341616 151852 341668 151904
rect 345112 151852 345164 151904
rect 180248 151784 180300 151836
rect 213920 151784 213972 151836
rect 257528 151784 257580 151836
rect 265808 151784 265860 151836
rect 231676 151716 231728 151768
rect 252652 151716 252704 151768
rect 281908 151716 281960 151768
rect 284392 151716 284444 151768
rect 342260 151716 342312 151768
rect 346676 151716 346728 151768
rect 430580 151716 430632 151768
rect 465724 151716 465776 151768
rect 231768 151648 231820 151700
rect 249892 151648 249944 151700
rect 282276 151104 282328 151156
rect 285864 151104 285916 151156
rect 332048 151036 332100 151088
rect 342260 151036 342312 151088
rect 249156 150492 249208 150544
rect 265808 150492 265860 150544
rect 235448 150424 235500 150476
rect 265900 150424 265952 150476
rect 3424 150356 3476 150408
rect 22744 150356 22796 150408
rect 169024 150356 169076 150408
rect 213920 150356 213972 150408
rect 231676 150356 231728 150408
rect 259460 150356 259512 150408
rect 282736 150356 282788 150408
rect 310520 150356 310572 150408
rect 430580 150356 430632 150408
rect 437664 150356 437716 150408
rect 282828 150288 282880 150340
rect 294236 150288 294288 150340
rect 430856 150288 430908 150340
rect 436100 150288 436152 150340
rect 231768 149812 231820 149864
rect 236000 149812 236052 149864
rect 235264 149676 235316 149728
rect 265992 149676 266044 149728
rect 323584 149676 323636 149728
rect 342260 149676 342312 149728
rect 249248 149132 249300 149184
rect 265256 149132 265308 149184
rect 342260 149132 342312 149184
rect 347504 149132 347556 149184
rect 239588 149064 239640 149116
rect 265900 149064 265952 149116
rect 167644 148996 167696 149048
rect 213920 148996 213972 149048
rect 282828 148996 282880 149048
rect 296904 148996 296956 149048
rect 430580 148996 430632 149048
rect 434904 148996 434956 149048
rect 231308 148928 231360 148980
rect 234620 148928 234672 148980
rect 177488 148316 177540 148368
rect 214012 148316 214064 148368
rect 256240 148316 256292 148368
rect 265808 148316 265860 148368
rect 231216 147704 231268 147756
rect 238024 147704 238076 147756
rect 246488 147704 246540 147756
rect 265716 147704 265768 147756
rect 191196 147636 191248 147688
rect 213920 147636 213972 147688
rect 236920 147636 236972 147688
rect 265440 147636 265492 147688
rect 282828 147568 282880 147620
rect 289912 147568 289964 147620
rect 336004 146956 336056 147008
rect 338212 146956 338264 147008
rect 346676 146888 346728 146940
rect 167644 146276 167696 146328
rect 213920 146276 213972 146328
rect 235540 146276 235592 146328
rect 265716 146276 265768 146328
rect 282828 146208 282880 146260
rect 311900 146208 311952 146260
rect 430580 146208 430632 146260
rect 436284 146208 436336 146260
rect 231768 146140 231820 146192
rect 247040 146140 247092 146192
rect 282736 146140 282788 146192
rect 291200 146140 291252 146192
rect 231400 146072 231452 146124
rect 256792 146072 256844 146124
rect 230848 146004 230900 146056
rect 232688 146004 232740 146056
rect 232596 145528 232648 145580
rect 265532 145528 265584 145580
rect 313924 145528 313976 145580
rect 346676 145528 346728 145580
rect 232504 145052 232556 145104
rect 265808 145052 265860 145104
rect 196808 144984 196860 145036
rect 213920 144984 213972 145036
rect 242348 144984 242400 145036
rect 265900 144984 265952 145036
rect 171784 144916 171836 144968
rect 214012 144916 214064 144968
rect 282736 144848 282788 144900
rect 311992 144848 312044 144900
rect 430580 144848 430632 144900
rect 441712 144848 441764 144900
rect 282828 144780 282880 144832
rect 298284 144780 298336 144832
rect 430856 144780 430908 144832
rect 440424 144780 440476 144832
rect 300860 144168 300912 144220
rect 346308 144168 346360 144220
rect 231768 143964 231820 144016
rect 234804 143964 234856 144016
rect 264520 143692 264572 143744
rect 266084 143692 266136 143744
rect 210424 143624 210476 143676
rect 214012 143624 214064 143676
rect 253112 143624 253164 143676
rect 265532 143624 265584 143676
rect 176016 143556 176068 143608
rect 213920 143556 213972 143608
rect 235356 143556 235408 143608
rect 265808 143556 265860 143608
rect 344928 143556 344980 143608
rect 346676 143556 346728 143608
rect 231768 143488 231820 143540
rect 253940 143488 253992 143540
rect 282092 143488 282144 143540
rect 307760 143488 307812 143540
rect 233976 142876 234028 142928
rect 265716 142876 265768 142928
rect 169024 142808 169076 142860
rect 214104 142808 214156 142860
rect 230020 142808 230072 142860
rect 264428 142808 264480 142860
rect 322204 142808 322256 142860
rect 346584 142808 346636 142860
rect 282828 142468 282880 142520
rect 287336 142468 287388 142520
rect 254676 142196 254728 142248
rect 265532 142196 265584 142248
rect 195428 142128 195480 142180
rect 213920 142128 213972 142180
rect 253480 142128 253532 142180
rect 265624 142128 265676 142180
rect 430580 142128 430632 142180
rect 436100 142128 436152 142180
rect 231492 142060 231544 142112
rect 251180 142060 251232 142112
rect 282736 142060 282788 142112
rect 296812 142060 296864 142112
rect 231768 141992 231820 142044
rect 248604 141992 248656 142044
rect 300124 141380 300176 141432
rect 343824 141380 343876 141432
rect 346492 141380 346544 141432
rect 282828 141312 282880 141364
rect 287152 141312 287204 141364
rect 259184 140904 259236 140956
rect 264612 140904 264664 140956
rect 206376 140836 206428 140888
rect 213920 140836 213972 140888
rect 232688 140836 232740 140888
rect 264428 140836 264480 140888
rect 171876 140768 171928 140820
rect 214012 140768 214064 140820
rect 232780 140768 232832 140820
rect 265808 140768 265860 140820
rect 282828 140700 282880 140752
rect 309140 140700 309192 140752
rect 430580 140700 430632 140752
rect 445760 140700 445812 140752
rect 178868 140020 178920 140072
rect 214656 140020 214708 140072
rect 231400 140020 231452 140072
rect 240968 140020 241020 140072
rect 241060 140020 241112 140072
rect 265716 140020 265768 140072
rect 445760 140020 445812 140072
rect 493324 140020 493376 140072
rect 265716 139884 265768 139936
rect 266176 139884 266228 139936
rect 231308 139748 231360 139800
rect 236184 139748 236236 139800
rect 257436 139476 257488 139528
rect 265256 139476 265308 139528
rect 209136 139408 209188 139460
rect 213920 139408 213972 139460
rect 229928 139408 229980 139460
rect 265900 139408 265952 139460
rect 282736 139340 282788 139392
rect 305184 139340 305236 139392
rect 461676 139340 461728 139392
rect 580172 139340 580224 139392
rect 231308 139272 231360 139324
rect 233332 139272 233384 139324
rect 282828 139272 282880 139324
rect 299480 139272 299532 139324
rect 231768 139204 231820 139256
rect 247132 139204 247184 139256
rect 231584 138660 231636 138712
rect 242256 138660 242308 138712
rect 327724 138660 327776 138712
rect 346400 138660 346452 138712
rect 347136 138660 347188 138712
rect 436744 138660 436796 138712
rect 460940 138660 460992 138712
rect 461676 138660 461728 138712
rect 231492 138252 231544 138304
rect 236092 138252 236144 138304
rect 247776 138116 247828 138168
rect 264428 138116 264480 138168
rect 243636 138048 243688 138100
rect 265164 138048 265216 138100
rect 238024 137980 238076 138032
rect 265440 137980 265492 138032
rect 429752 137980 429804 138032
rect 436652 137980 436704 138032
rect 3240 137912 3292 137964
rect 17224 137912 17276 137964
rect 231400 137912 231452 137964
rect 258080 137912 258132 137964
rect 282828 137912 282880 137964
rect 305000 137912 305052 137964
rect 430856 137912 430908 137964
rect 436744 137912 436796 137964
rect 231768 137844 231820 137896
rect 254032 137844 254084 137896
rect 282276 137776 282328 137828
rect 285680 137776 285732 137828
rect 174636 137232 174688 137284
rect 213920 137232 213972 137284
rect 234252 137232 234304 137284
rect 265716 137232 265768 137284
rect 334716 137232 334768 137284
rect 343732 137232 343784 137284
rect 430580 137232 430632 137284
rect 436652 137232 436704 137284
rect 580264 137232 580316 137284
rect 436192 137164 436244 137216
rect 436744 137164 436796 137216
rect 343732 136688 343784 136740
rect 346676 136688 346728 136740
rect 229836 136620 229888 136672
rect 264428 136620 264480 136672
rect 231400 136552 231452 136604
rect 250444 136552 250496 136604
rect 282368 136552 282420 136604
rect 306380 136552 306432 136604
rect 331864 136552 331916 136604
rect 337384 136552 337436 136604
rect 430580 136552 430632 136604
rect 431132 136552 431184 136604
rect 468484 136552 468536 136604
rect 230756 136484 230808 136536
rect 246396 136484 246448 136536
rect 295984 135872 296036 135924
rect 340972 135872 341024 135924
rect 261668 135464 261720 135516
rect 265808 135464 265860 135516
rect 254768 135396 254820 135448
rect 264428 135396 264480 135448
rect 184296 135328 184348 135380
rect 213920 135328 213972 135380
rect 246580 135328 246632 135380
rect 261116 135328 261168 135380
rect 173256 135260 173308 135312
rect 214012 135260 214064 135312
rect 236644 135260 236696 135312
rect 260932 135260 260984 135312
rect 340972 135260 341024 135312
rect 347504 135260 347556 135312
rect 231768 135192 231820 135244
rect 256056 135192 256108 135244
rect 282736 135192 282788 135244
rect 300952 135192 301004 135244
rect 430580 135192 430632 135244
rect 446404 135192 446456 135244
rect 231676 135124 231728 135176
rect 244924 135124 244976 135176
rect 282828 135124 282880 135176
rect 298192 135124 298244 135176
rect 230572 135056 230624 135108
rect 239404 135056 239456 135108
rect 255964 134036 256016 134088
rect 265716 134036 265768 134088
rect 245108 133968 245160 134020
rect 265532 133968 265584 134020
rect 181444 133900 181496 133952
rect 213920 133900 213972 133952
rect 236828 133900 236880 133952
rect 265808 133900 265860 133952
rect 231768 133832 231820 133884
rect 260104 133832 260156 133884
rect 282000 133832 282052 133884
rect 310612 133832 310664 133884
rect 430580 133832 430632 133884
rect 485044 133832 485096 133884
rect 231676 133764 231728 133816
rect 243820 133764 243872 133816
rect 282184 133424 282236 133476
rect 284300 133424 284352 133476
rect 259092 133152 259144 133204
rect 265992 133152 266044 133204
rect 309784 133152 309836 133204
rect 346584 133152 346636 133204
rect 180156 132540 180208 132592
rect 214012 132540 214064 132592
rect 250444 132540 250496 132592
rect 265900 132540 265952 132592
rect 170588 132472 170640 132524
rect 213920 132472 213972 132524
rect 243544 132472 243596 132524
rect 265716 132472 265768 132524
rect 231676 132404 231728 132456
rect 259000 132404 259052 132456
rect 282828 132404 282880 132456
rect 314660 132404 314712 132456
rect 430580 132404 430632 132456
rect 452660 132404 452712 132456
rect 230664 132336 230716 132388
rect 258724 132336 258776 132388
rect 430856 132336 430908 132388
rect 440240 132336 440292 132388
rect 231768 132268 231820 132320
rect 250536 132268 250588 132320
rect 320824 131724 320876 131776
rect 345204 131724 345256 131776
rect 347412 131724 347464 131776
rect 282276 131316 282328 131368
rect 288624 131316 288676 131368
rect 258816 131248 258868 131300
rect 265716 131248 265768 131300
rect 258908 131180 258960 131232
rect 265440 131180 265492 131232
rect 193864 131112 193916 131164
rect 213920 131112 213972 131164
rect 253388 131112 253440 131164
rect 265900 131112 265952 131164
rect 231768 131044 231820 131096
rect 251916 131044 251968 131096
rect 231400 130976 231452 131028
rect 242164 130976 242216 131028
rect 231584 130364 231636 130416
rect 263140 130364 263192 130416
rect 281632 129820 281684 129872
rect 288440 129820 288492 129872
rect 251824 129752 251876 129804
rect 265256 129752 265308 129804
rect 231768 129684 231820 129736
rect 247868 129684 247920 129736
rect 282828 129684 282880 129736
rect 309324 129684 309376 129736
rect 430580 129684 430632 129736
rect 444380 129684 444432 129736
rect 231400 129616 231452 129668
rect 246672 129616 246724 129668
rect 207664 128392 207716 128444
rect 213920 128392 213972 128444
rect 247684 128392 247736 128444
rect 264428 128392 264480 128444
rect 173164 128324 173216 128376
rect 214012 128324 214064 128376
rect 246396 128324 246448 128376
rect 265716 128324 265768 128376
rect 231676 128256 231728 128308
rect 249064 128256 249116 128308
rect 281632 128256 281684 128308
rect 307852 128256 307904 128308
rect 312544 128256 312596 128308
rect 347964 128256 348016 128308
rect 231768 128188 231820 128240
rect 243728 128188 243780 128240
rect 231492 127576 231544 127628
rect 252100 127576 252152 127628
rect 287060 127576 287112 127628
rect 345112 127576 345164 127628
rect 282276 127440 282328 127492
rect 285772 127440 285824 127492
rect 252008 127032 252060 127084
rect 265900 127032 265952 127084
rect 250536 126964 250588 127016
rect 264428 126964 264480 127016
rect 231676 126896 231728 126948
rect 253204 126896 253256 126948
rect 282828 126896 282880 126948
rect 301044 126896 301096 126948
rect 323676 126896 323728 126948
rect 347688 126896 347740 126948
rect 447784 126896 447836 126948
rect 580172 126896 580224 126948
rect 231768 126828 231820 126880
rect 245016 126828 245068 126880
rect 305644 126216 305696 126268
rect 347688 126216 347740 126268
rect 180340 125672 180392 125724
rect 214012 125672 214064 125724
rect 59268 125604 59320 125656
rect 65156 125604 65208 125656
rect 176108 125604 176160 125656
rect 213920 125604 213972 125656
rect 254860 125604 254912 125656
rect 265900 125604 265952 125656
rect 231308 125536 231360 125588
rect 264244 125536 264296 125588
rect 282828 125536 282880 125588
rect 292580 125536 292632 125588
rect 430580 125536 430632 125588
rect 439044 125536 439096 125588
rect 231676 125468 231728 125520
rect 263048 125468 263100 125520
rect 311900 124856 311952 124908
rect 343824 124856 343876 124908
rect 170680 124244 170732 124296
rect 213920 124244 213972 124296
rect 264612 124244 264664 124296
rect 265624 124244 265676 124296
rect 169116 124176 169168 124228
rect 214012 124176 214064 124228
rect 242164 124176 242216 124228
rect 265900 124176 265952 124228
rect 231492 124108 231544 124160
rect 260196 124108 260248 124160
rect 338764 124108 338816 124160
rect 348976 124108 349028 124160
rect 430580 124108 430632 124160
rect 443184 124108 443236 124160
rect 231308 124040 231360 124092
rect 250628 124040 250680 124092
rect 231308 123428 231360 123480
rect 257344 123428 257396 123480
rect 325700 123428 325752 123480
rect 338304 123428 338356 123480
rect 261484 123088 261536 123140
rect 265900 123088 265952 123140
rect 177396 122884 177448 122936
rect 214012 122884 214064 122936
rect 260104 122884 260156 122936
rect 265900 122884 265952 122936
rect 167828 122816 167880 122868
rect 213920 122816 213972 122868
rect 256148 122816 256200 122868
rect 265992 122816 266044 122868
rect 231768 122748 231820 122800
rect 256332 122748 256384 122800
rect 430580 122748 430632 122800
rect 449900 122748 449952 122800
rect 231492 122680 231544 122732
rect 246304 122680 246356 122732
rect 282828 122680 282880 122732
rect 303712 122680 303764 122732
rect 231584 122612 231636 122664
rect 234068 122612 234120 122664
rect 257344 121592 257396 121644
rect 264244 121592 264296 121644
rect 172060 121524 172112 121576
rect 213920 121524 213972 121576
rect 249064 121524 249116 121576
rect 265992 121524 266044 121576
rect 170496 121456 170548 121508
rect 214012 121456 214064 121508
rect 233884 121456 233936 121508
rect 265900 121456 265952 121508
rect 231768 121388 231820 121440
rect 253296 121388 253348 121440
rect 281908 121388 281960 121440
rect 309232 121388 309284 121440
rect 430580 121388 430632 121440
rect 437572 121388 437624 121440
rect 231492 121320 231544 121372
rect 240784 121320 240836 121372
rect 281632 121320 281684 121372
rect 303620 121320 303672 121372
rect 231124 120912 231176 120964
rect 238116 120912 238168 120964
rect 430580 120844 430632 120896
rect 433340 120844 433392 120896
rect 170404 120708 170456 120760
rect 203524 120708 203576 120760
rect 260196 120232 260248 120284
rect 265532 120232 265584 120284
rect 178776 120164 178828 120216
rect 214012 120164 214064 120216
rect 253204 120164 253256 120216
rect 265716 120164 265768 120216
rect 173440 120096 173492 120148
rect 213920 120096 213972 120148
rect 239404 120096 239456 120148
rect 265624 120096 265676 120148
rect 231768 120028 231820 120080
rect 261576 120028 261628 120080
rect 282092 120028 282144 120080
rect 294144 120028 294196 120080
rect 315304 120028 315356 120080
rect 347044 120028 347096 120080
rect 231400 119960 231452 120012
rect 239496 119960 239548 120012
rect 430580 119892 430632 119944
rect 433524 119892 433576 119944
rect 231308 119348 231360 119400
rect 259184 119348 259236 119400
rect 210516 118804 210568 118856
rect 214104 118804 214156 118856
rect 185584 118736 185636 118788
rect 213920 118736 213972 118788
rect 258724 118736 258776 118788
rect 265716 118736 265768 118788
rect 178960 118668 179012 118720
rect 214012 118668 214064 118720
rect 246304 118668 246356 118720
rect 265624 118668 265676 118720
rect 231492 118600 231544 118652
rect 245292 118600 245344 118652
rect 282460 118600 282512 118652
rect 305092 118600 305144 118652
rect 231768 118532 231820 118584
rect 245200 118532 245252 118584
rect 231124 118464 231176 118516
rect 239680 118464 239732 118516
rect 430580 118396 430632 118448
rect 432236 118396 432288 118448
rect 282828 117988 282880 118040
rect 287244 117988 287296 118040
rect 318800 117920 318852 117972
rect 343732 117920 343784 117972
rect 244924 117444 244976 117496
rect 265992 117444 266044 117496
rect 177580 117376 177632 117428
rect 213920 117376 213972 117428
rect 245016 117376 245068 117428
rect 265716 117376 265768 117428
rect 166356 117308 166408 117360
rect 214012 117308 214064 117360
rect 239496 117308 239548 117360
rect 265348 117308 265400 117360
rect 231492 117240 231544 117292
rect 242440 117240 242492 117292
rect 282552 117240 282604 117292
rect 302240 117240 302292 117292
rect 430580 117240 430632 117292
rect 448612 117240 448664 117292
rect 231216 116764 231268 116816
rect 238300 116764 238352 116816
rect 231124 116560 231176 116612
rect 241152 116560 241204 116612
rect 323032 116560 323084 116612
rect 340972 116560 341024 116612
rect 256056 116084 256108 116136
rect 266084 116084 266136 116136
rect 176200 116016 176252 116068
rect 213920 116016 213972 116068
rect 242256 116016 242308 116068
rect 265992 116016 266044 116068
rect 173348 115948 173400 116000
rect 214012 115948 214064 116000
rect 240968 115948 241020 116000
rect 265716 115948 265768 116000
rect 282552 115880 282604 115932
rect 306472 115880 306524 115932
rect 330484 115880 330536 115932
rect 347504 115880 347556 115932
rect 430580 115880 430632 115932
rect 434812 115880 434864 115932
rect 282828 115812 282880 115864
rect 302332 115812 302384 115864
rect 230664 115744 230716 115796
rect 240876 115744 240928 115796
rect 231676 115472 231728 115524
rect 238208 115472 238260 115524
rect 230572 114792 230624 114844
rect 232596 114792 232648 114844
rect 247868 114656 247920 114708
rect 265992 114656 266044 114708
rect 209228 114588 209280 114640
rect 213920 114588 213972 114640
rect 240784 114588 240836 114640
rect 265716 114588 265768 114640
rect 169208 114520 169260 114572
rect 214012 114520 214064 114572
rect 238300 114520 238352 114572
rect 265256 114520 265308 114572
rect 231768 114452 231820 114504
rect 252192 114452 252244 114504
rect 430856 114452 430908 114504
rect 447140 114452 447192 114504
rect 230572 114384 230624 114436
rect 234160 114384 234212 114436
rect 430580 114384 430632 114436
rect 445852 114384 445904 114436
rect 230664 113772 230716 113824
rect 249156 113772 249208 113824
rect 252100 113296 252152 113348
rect 265716 113296 265768 113348
rect 198188 113228 198240 113280
rect 213920 113228 213972 113280
rect 251916 113228 251968 113280
rect 265256 113228 265308 113280
rect 167736 113160 167788 113212
rect 214012 113160 214064 113212
rect 229744 113160 229796 113212
rect 265716 113160 265768 113212
rect 282092 113092 282144 113144
rect 295340 113092 295392 113144
rect 231768 112820 231820 112872
rect 236736 112820 236788 112872
rect 230572 112480 230624 112532
rect 249248 112480 249300 112532
rect 231124 112412 231176 112464
rect 264336 112412 264388 112464
rect 188528 111868 188580 111920
rect 213920 111868 213972 111920
rect 181536 111800 181588 111852
rect 214012 111800 214064 111852
rect 249156 111800 249208 111852
rect 265716 111800 265768 111852
rect 3424 111732 3476 111784
rect 14464 111732 14516 111784
rect 167920 111732 167972 111784
rect 177488 111732 177540 111784
rect 231768 111732 231820 111784
rect 264520 111732 264572 111784
rect 282828 111732 282880 111784
rect 296720 111732 296772 111784
rect 430580 111732 430632 111784
rect 451280 111732 451332 111784
rect 231492 111664 231544 111716
rect 235264 111664 235316 111716
rect 316040 111052 316092 111104
rect 327724 111052 327776 111104
rect 329840 111052 329892 111104
rect 345204 111052 345256 111104
rect 238208 110576 238260 110628
rect 265992 110576 266044 110628
rect 207756 110508 207808 110560
rect 214012 110508 214064 110560
rect 166264 110440 166316 110492
rect 213920 110440 213972 110492
rect 260288 110440 260340 110492
rect 265716 110440 265768 110492
rect 168104 110372 168156 110424
rect 178868 110372 178920 110424
rect 231768 110372 231820 110424
rect 257528 110372 257580 110424
rect 282276 110372 282328 110424
rect 294052 110372 294104 110424
rect 344284 110372 344336 110424
rect 347044 110372 347096 110424
rect 231768 109964 231820 110016
rect 235448 109964 235500 110016
rect 257620 109148 257672 109200
rect 265716 109148 265768 109200
rect 206468 109080 206520 109132
rect 214012 109080 214064 109132
rect 235264 109080 235316 109132
rect 265164 109080 265216 109132
rect 171968 109012 172020 109064
rect 213920 109012 213972 109064
rect 234068 109012 234120 109064
rect 265532 109012 265584 109064
rect 167920 108944 167972 108996
rect 180248 108944 180300 108996
rect 231768 108944 231820 108996
rect 260380 108944 260432 108996
rect 301504 108944 301556 108996
rect 347504 108944 347556 108996
rect 430580 108944 430632 108996
rect 434720 108944 434772 108996
rect 231676 108876 231728 108928
rect 239588 108876 239640 108928
rect 231400 108264 231452 108316
rect 253480 108264 253532 108316
rect 240876 107856 240928 107908
rect 265716 107856 265768 107908
rect 281540 107856 281592 107908
rect 283196 107856 283248 107908
rect 261576 107788 261628 107840
rect 265992 107788 266044 107840
rect 178868 107720 178920 107772
rect 214012 107720 214064 107772
rect 253296 107720 253348 107772
rect 265716 107720 265768 107772
rect 174728 107652 174780 107704
rect 213920 107652 213972 107704
rect 263048 107652 263100 107704
rect 265164 107652 265216 107704
rect 231768 107584 231820 107636
rect 256240 107584 256292 107636
rect 333336 107584 333388 107636
rect 347504 107584 347556 107636
rect 430580 107584 430632 107636
rect 443000 107584 443052 107636
rect 231676 107516 231728 107568
rect 246488 107516 246540 107568
rect 231768 107040 231820 107092
rect 236920 107040 236972 107092
rect 177488 106360 177540 106412
rect 214012 106360 214064 106412
rect 249248 106360 249300 106412
rect 265532 106360 265584 106412
rect 170404 106292 170456 106344
rect 213920 106292 213972 106344
rect 245200 106292 245252 106344
rect 265716 106292 265768 106344
rect 231768 106224 231820 106276
rect 261852 106224 261904 106276
rect 262864 106224 262916 106276
rect 267188 106224 267240 106276
rect 430580 106224 430632 106276
rect 438860 106224 438912 106276
rect 231676 105340 231728 105392
rect 235540 105340 235592 105392
rect 192576 105000 192628 105052
rect 214012 105000 214064 105052
rect 261760 105000 261812 105052
rect 265532 105000 265584 105052
rect 205088 104932 205140 104984
rect 213920 104932 213972 104984
rect 256240 104932 256292 104984
rect 265992 104932 266044 104984
rect 239588 104864 239640 104916
rect 265716 104864 265768 104916
rect 231768 104796 231820 104848
rect 264612 104796 264664 104848
rect 282000 104796 282052 104848
rect 284484 104796 284536 104848
rect 311164 104796 311216 104848
rect 347044 104796 347096 104848
rect 430580 104796 430632 104848
rect 441620 104796 441672 104848
rect 231492 104728 231544 104780
rect 242348 104728 242400 104780
rect 231676 104660 231728 104712
rect 234252 104660 234304 104712
rect 262864 103708 262916 103760
rect 265992 103708 266044 103760
rect 242440 103640 242492 103692
rect 265716 103640 265768 103692
rect 202328 103572 202380 103624
rect 214012 103572 214064 103624
rect 199384 103504 199436 103556
rect 213920 103504 213972 103556
rect 430580 103436 430632 103488
rect 440332 103436 440384 103488
rect 430764 103368 430816 103420
rect 437480 103368 437532 103420
rect 230572 102960 230624 103012
rect 232504 102960 232556 103012
rect 175924 102756 175976 102808
rect 216220 102756 216272 102808
rect 293960 102756 294012 102808
rect 342260 102756 342312 102808
rect 253480 102348 253532 102400
rect 264612 102348 264664 102400
rect 233608 102280 233660 102332
rect 266084 102280 266136 102332
rect 232596 102212 232648 102264
rect 265716 102212 265768 102264
rect 200856 102144 200908 102196
rect 213920 102144 213972 102196
rect 231124 102144 231176 102196
rect 265164 102144 265216 102196
rect 231492 102076 231544 102128
rect 233976 102076 234028 102128
rect 282828 102076 282880 102128
rect 290096 102076 290148 102128
rect 336280 102076 336332 102128
rect 347228 102076 347280 102128
rect 430580 102076 430632 102128
rect 448520 102076 448572 102128
rect 231768 101940 231820 101992
rect 259092 101940 259144 101992
rect 231584 101464 231636 101516
rect 235356 101464 235408 101516
rect 231676 101396 231728 101448
rect 254676 101396 254728 101448
rect 280436 101396 280488 101448
rect 343640 101396 343692 101448
rect 259000 100852 259052 100904
rect 265716 100852 265768 100904
rect 257528 100784 257580 100836
rect 265348 100784 265400 100836
rect 203708 100716 203760 100768
rect 213920 100716 213972 100768
rect 246488 100716 246540 100768
rect 265532 100716 265584 100768
rect 231768 100648 231820 100700
rect 241060 100648 241112 100700
rect 319444 100648 319496 100700
rect 347504 100648 347556 100700
rect 436744 100648 436796 100700
rect 580172 100648 580224 100700
rect 284300 99968 284352 100020
rect 345020 99968 345072 100020
rect 230940 99560 230992 99612
rect 232780 99560 232832 99612
rect 254676 99492 254728 99544
rect 265532 99492 265584 99544
rect 169300 99424 169352 99476
rect 213920 99424 213972 99476
rect 238116 99424 238168 99476
rect 265716 99424 265768 99476
rect 164884 99356 164936 99408
rect 214012 99356 214064 99408
rect 236736 99356 236788 99408
rect 265992 99356 266044 99408
rect 230480 98200 230532 98252
rect 232688 98200 232740 98252
rect 248972 98132 249024 98184
rect 266084 98132 266136 98184
rect 167920 98064 167972 98116
rect 214012 98064 214064 98116
rect 232504 98064 232556 98116
rect 264612 98064 264664 98116
rect 166448 97996 166500 98048
rect 213920 97996 213972 98048
rect 231216 97996 231268 98048
rect 265624 97996 265676 98048
rect 316684 97928 316736 97980
rect 347504 97928 347556 97980
rect 430580 97928 430632 97980
rect 443092 97928 443144 97980
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 166540 97248 166592 97300
rect 214656 97248 214708 97300
rect 231768 96704 231820 96756
rect 239680 96704 239732 96756
rect 260380 96704 260432 96756
rect 264612 96704 264664 96756
rect 210608 96636 210660 96688
rect 213920 96636 213972 96688
rect 230480 96636 230532 96688
rect 233976 96636 234028 96688
rect 235356 96636 235408 96688
rect 261392 96636 261444 96688
rect 348884 96568 348936 96620
rect 580356 96568 580408 96620
rect 329104 96500 329156 96552
rect 428096 96500 428148 96552
rect 188436 96364 188488 96416
rect 281540 96364 281592 96416
rect 226984 95888 227036 95940
rect 248972 95888 249024 95940
rect 204996 95208 205048 95260
rect 213920 95208 213972 95260
rect 228364 95208 228416 95260
rect 265532 95208 265584 95260
rect 318064 95208 318116 95260
rect 389456 95208 389508 95260
rect 209044 95140 209096 95192
rect 427636 95140 427688 95192
rect 196716 95072 196768 95124
rect 280160 95072 280212 95124
rect 326344 95072 326396 95124
rect 428188 95072 428240 95124
rect 203616 95004 203668 95056
rect 280252 95004 280304 95056
rect 342904 95004 342956 95056
rect 400220 95004 400272 95056
rect 400864 95004 400916 95056
rect 340144 94936 340196 94988
rect 396172 94936 396224 94988
rect 397092 94936 397144 94988
rect 222844 94528 222896 94580
rect 233608 94528 233660 94580
rect 130384 94460 130436 94512
rect 214564 94460 214616 94512
rect 224224 94460 224276 94512
rect 267280 94460 267332 94512
rect 120632 94052 120684 94104
rect 167828 94052 167880 94104
rect 118240 93984 118292 94036
rect 172060 93984 172112 94036
rect 106648 93916 106700 93968
rect 170588 93916 170640 93968
rect 93860 93848 93912 93900
rect 174728 93848 174780 93900
rect 67640 93780 67692 93832
rect 199384 93780 199436 93832
rect 239680 93780 239732 93832
rect 270960 93780 271012 93832
rect 347688 93780 347740 93832
rect 582380 93780 582432 93832
rect 195336 93712 195388 93764
rect 281908 93712 281960 93764
rect 349804 93712 349856 93764
rect 360200 93712 360252 93764
rect 233976 93644 234028 93696
rect 276940 93644 276992 93696
rect 345664 93644 345716 93696
rect 356520 93644 356572 93696
rect 349896 93576 349948 93628
rect 358820 93576 358872 93628
rect 270960 93440 271012 93492
rect 351460 93440 351512 93492
rect 151728 93372 151780 93424
rect 187056 93372 187108 93424
rect 114376 93304 114428 93356
rect 173256 93304 173308 93356
rect 129464 93236 129516 93288
rect 176016 93236 176068 93288
rect 113824 93168 113876 93220
rect 185584 93168 185636 93220
rect 118700 93100 118752 93152
rect 214748 93100 214800 93152
rect 399484 93100 399536 93152
rect 406016 93100 406068 93152
rect 410524 93100 410576 93152
rect 427452 93100 427504 93152
rect 348424 92692 348476 92744
rect 353300 92692 353352 92744
rect 354036 92692 354088 92744
rect 356060 92488 356112 92540
rect 356520 92488 356572 92540
rect 395344 92488 395396 92540
rect 396080 92488 396132 92540
rect 396724 92488 396776 92540
rect 399576 92488 399628 92540
rect 406384 92488 406436 92540
rect 408500 92488 408552 92540
rect 88984 92420 89036 92472
rect 164884 92420 164936 92472
rect 192484 92420 192536 92472
rect 357440 92420 357492 92472
rect 202236 92352 202288 92404
rect 281632 92352 281684 92404
rect 337476 92352 337528 92404
rect 394700 92352 394752 92404
rect 98184 92284 98236 92336
rect 118700 92284 118752 92336
rect 133144 92284 133196 92336
rect 169024 92284 169076 92336
rect 178684 92284 178736 92336
rect 281724 92284 281776 92336
rect 298744 92284 298796 92336
rect 352012 92284 352064 92336
rect 125968 92216 126020 92268
rect 195428 92216 195480 92268
rect 216220 92216 216272 92268
rect 280344 92216 280396 92268
rect 115848 92148 115900 92200
rect 130384 92148 130436 92200
rect 136088 92148 136140 92200
rect 191196 92148 191248 92200
rect 152096 92080 152148 92132
rect 189724 92080 189776 92132
rect 84384 92012 84436 92064
rect 203708 92012 203760 92064
rect 352012 91740 352064 91792
rect 352748 91740 352800 91792
rect 74816 91060 74868 91112
rect 135904 91060 135956 91112
rect 105912 90992 105964 91044
rect 193864 90992 193916 91044
rect 316868 90992 316920 91044
rect 391940 90992 391992 91044
rect 111616 90924 111668 90976
rect 166356 90924 166408 90976
rect 126520 90856 126572 90908
rect 180340 90856 180392 90908
rect 122840 90788 122892 90840
rect 170680 90788 170732 90840
rect 124588 90720 124640 90772
rect 171876 90720 171928 90772
rect 151544 90652 151596 90704
rect 198096 90652 198148 90704
rect 298100 90312 298152 90364
rect 366640 90312 366692 90364
rect 65984 89632 66036 89684
rect 210608 89632 210660 89684
rect 100576 89564 100628 89616
rect 207756 89564 207808 89616
rect 102876 89496 102928 89548
rect 198188 89496 198240 89548
rect 115848 89428 115900 89480
rect 178960 89428 179012 89480
rect 132408 89360 132460 89412
rect 171784 89360 171836 89412
rect 291844 89020 291896 89072
rect 327080 89020 327132 89072
rect 355324 89020 355376 89072
rect 198096 88952 198148 89004
rect 265900 88952 265952 89004
rect 300216 88952 300268 89004
rect 351920 88952 351972 89004
rect 388168 88952 388220 89004
rect 411260 88952 411312 89004
rect 412272 88952 412324 89004
rect 101864 88272 101916 88324
rect 181536 88272 181588 88324
rect 230572 88272 230624 88324
rect 233976 88272 234028 88324
rect 85856 88204 85908 88256
rect 166448 88204 166500 88256
rect 107200 88136 107252 88188
rect 169208 88136 169260 88188
rect 117136 88068 117188 88120
rect 178776 88068 178828 88120
rect 151636 88000 151688 88052
rect 211804 88000 211856 88052
rect 135076 87932 135128 87984
rect 167644 87932 167696 87984
rect 198004 87592 198056 87644
rect 302240 87592 302292 87644
rect 365720 87592 365772 87644
rect 67732 86912 67784 86964
rect 214932 86912 214984 86964
rect 439504 86912 439556 86964
rect 580172 86912 580224 86964
rect 100668 86844 100720 86896
rect 188528 86844 188580 86896
rect 128176 86776 128228 86828
rect 210424 86776 210476 86828
rect 88064 86708 88116 86760
rect 169300 86708 169352 86760
rect 110144 86640 110196 86692
rect 177580 86640 177632 86692
rect 115756 86572 115808 86624
rect 173440 86572 173492 86624
rect 276020 86232 276072 86284
rect 342352 86232 342404 86284
rect 345020 86232 345072 86284
rect 428004 86232 428056 86284
rect 3148 85484 3200 85536
rect 46940 85484 46992 85536
rect 67548 85484 67600 85536
rect 200856 85484 200908 85536
rect 304264 85484 304316 85536
rect 305000 85484 305052 85536
rect 90640 85416 90692 85468
rect 213460 85416 213512 85468
rect 118240 85348 118292 85400
rect 213368 85348 213420 85400
rect 92296 85280 92348 85332
rect 170404 85280 170456 85332
rect 125416 85212 125468 85264
rect 176108 85212 176160 85264
rect 305000 84804 305052 84856
rect 404360 84804 404412 84856
rect 67456 84124 67508 84176
rect 214840 84124 214892 84176
rect 122656 84056 122708 84108
rect 209136 84056 209188 84108
rect 108856 83988 108908 84040
rect 180156 83988 180208 84040
rect 99196 83920 99248 83972
rect 166264 83920 166316 83972
rect 104716 83852 104768 83904
rect 167736 83852 167788 83904
rect 119988 83784 120040 83836
rect 170496 83784 170548 83836
rect 291200 83512 291252 83564
rect 332048 83512 332100 83564
rect 325148 83444 325200 83496
rect 331220 83444 331272 83496
rect 397460 83444 397512 83496
rect 106096 82764 106148 82816
rect 209228 82764 209280 82816
rect 124036 82696 124088 82748
rect 206376 82696 206428 82748
rect 96528 82628 96580 82680
rect 171968 82628 172020 82680
rect 122748 82560 122800 82612
rect 177396 82560 177448 82612
rect 324320 82084 324372 82136
rect 396080 82084 396132 82136
rect 112996 81336 113048 81388
rect 210516 81336 210568 81388
rect 93768 81268 93820 81320
rect 177488 81268 177540 81320
rect 131028 81200 131080 81252
rect 196808 81200 196860 81252
rect 273260 80656 273312 80708
rect 340880 80656 340932 80708
rect 342260 80656 342312 80708
rect 390560 80656 390612 80708
rect 97908 79976 97960 80028
rect 206468 79976 206520 80028
rect 338120 79976 338172 80028
rect 393320 79976 393372 80028
rect 126888 79908 126940 79960
rect 213276 79908 213328 79960
rect 102048 79840 102100 79892
rect 173164 79840 173216 79892
rect 108948 79772 109000 79824
rect 176200 79772 176252 79824
rect 124128 79704 124180 79756
rect 169116 79704 169168 79756
rect 335360 79568 335412 79620
rect 338120 79568 338172 79620
rect 99288 78616 99340 78668
rect 207664 78616 207716 78668
rect 95148 78548 95200 78600
rect 178868 78548 178920 78600
rect 86868 78480 86920 78532
rect 167920 78480 167972 78532
rect 113088 78412 113140 78464
rect 184296 78412 184348 78464
rect 135904 78344 135956 78396
rect 204996 78344 205048 78396
rect 278044 77936 278096 77988
rect 372620 77936 372672 77988
rect 110236 77188 110288 77240
rect 181444 77188 181496 77240
rect 110328 77120 110380 77172
rect 173348 77120 173400 77172
rect 122840 76576 122892 76628
rect 254860 76576 254912 76628
rect 37280 76508 37332 76560
rect 240968 76508 241020 76560
rect 314108 76508 314160 76560
rect 328460 76508 328512 76560
rect 395344 76508 395396 76560
rect 59268 75828 59320 75880
rect 202328 75828 202380 75880
rect 317420 75828 317472 75880
rect 322940 75828 322992 75880
rect 396724 75828 396776 75880
rect 104900 75216 104952 75268
rect 256148 75216 256200 75268
rect 11060 75148 11112 75200
rect 260380 75148 260432 75200
rect 269120 75148 269172 75200
rect 318156 75148 318208 75200
rect 75920 73788 75972 73840
rect 249248 73788 249300 73840
rect 314660 73788 314712 73840
rect 400220 73788 400272 73840
rect 349988 73108 350040 73160
rect 579988 73108 580040 73160
rect 64420 72428 64472 72480
rect 311808 72428 311860 72480
rect 3424 71680 3476 71732
rect 57888 71680 57940 71732
rect 436100 71680 436152 71732
rect 60740 71000 60792 71052
rect 253388 71000 253440 71052
rect 110420 69708 110472 69760
rect 247776 69708 247828 69760
rect 98000 69640 98052 69692
rect 263140 69640 263192 69692
rect 311164 69640 311216 69692
rect 311808 69640 311860 69692
rect 401600 69640 401652 69692
rect 74540 68280 74592 68332
rect 245108 68280 245160 68332
rect 322204 68280 322256 68332
rect 402980 68280 403032 68332
rect 81440 66920 81492 66972
rect 236828 66920 236880 66972
rect 6920 66852 6972 66904
rect 226984 66852 227036 66904
rect 299664 66852 299716 66904
rect 399484 66852 399536 66904
rect 296720 66172 296772 66224
rect 297364 66172 297416 66224
rect 407120 66172 407172 66224
rect 46940 65560 46992 65612
rect 222844 65560 222896 65612
rect 85580 65492 85632 65544
rect 261668 65492 261720 65544
rect 215944 64268 215996 64320
rect 295340 64268 295392 64320
rect 87604 64200 87656 64252
rect 265808 64200 265860 64252
rect 51172 64132 51224 64184
rect 242440 64132 242492 64184
rect 409880 64132 409932 64184
rect 88340 62840 88392 62892
rect 254768 62840 254820 62892
rect 57980 62772 58032 62824
rect 264520 62772 264572 62824
rect 286324 62772 286376 62824
rect 411352 62772 411404 62824
rect 92480 61412 92532 61464
rect 246580 61412 246632 61464
rect 64880 61344 64932 61396
rect 239588 61344 239640 61396
rect 267096 61344 267148 61396
rect 280252 61344 280304 61396
rect 412640 61344 412692 61396
rect 113180 60120 113232 60172
rect 243636 60120 243688 60172
rect 69020 60052 69072 60104
rect 261760 60052 261812 60104
rect 4252 59984 4304 60036
rect 228364 59984 228416 60036
rect 276664 59984 276716 60036
rect 414020 59984 414072 60036
rect 3056 59304 3108 59356
rect 51080 59304 51132 59356
rect 111800 58692 111852 58744
rect 264428 58692 264480 58744
rect 71780 58624 71832 58676
rect 245200 58624 245252 58676
rect 267188 58624 267240 58676
rect 271880 58624 271932 58676
rect 415400 58624 415452 58676
rect 85672 57264 85724 57316
rect 240876 57264 240928 57316
rect 13820 57196 13872 57248
rect 252008 57196 252060 57248
rect 268384 57196 268436 57248
rect 416780 57196 416832 57248
rect 124220 55972 124272 56024
rect 257436 55972 257488 56024
rect 52460 55904 52512 55956
rect 258908 55904 258960 55956
rect 2780 55836 2832 55888
rect 229928 55836 229980 55888
rect 264428 55836 264480 55888
rect 419540 55836 419592 55888
rect 60832 54544 60884 54596
rect 256240 54544 256292 54596
rect 15200 54476 15252 54528
rect 235356 54476 235408 54528
rect 254584 54476 254636 54528
rect 422300 54476 422352 54528
rect 177304 53184 177356 53236
rect 251180 53184 251232 53236
rect 107660 53116 107712 53168
rect 260288 53116 260340 53168
rect 30380 53048 30432 53100
rect 247868 53048 247920 53100
rect 423680 53048 423732 53100
rect 118700 51756 118752 51808
rect 249156 51756 249208 51808
rect 17960 51688 18012 51740
rect 248512 51688 248564 51740
rect 425060 51756 425112 51808
rect 252100 51620 252152 51672
rect 313280 50396 313332 50448
rect 360200 50396 360252 50448
rect 19340 50328 19392 50380
rect 250536 50328 250588 50380
rect 259460 50328 259512 50380
rect 314016 50328 314068 50380
rect 347780 50328 347832 50380
rect 432052 50328 432104 50380
rect 96620 49036 96672 49088
rect 234068 49036 234120 49088
rect 309232 49036 309284 49088
rect 361580 49036 361632 49088
rect 56600 48968 56652 49020
rect 258816 48968 258868 49020
rect 340144 48968 340196 49020
rect 394700 48968 394752 49020
rect 93860 47608 93912 47660
rect 263048 47608 263100 47660
rect 44180 47540 44232 47592
rect 242256 47540 242308 47592
rect 302884 47540 302936 47592
rect 364340 47540 364392 47592
rect 464344 46860 464396 46912
rect 580172 46860 580224 46912
rect 117320 46316 117372 46368
rect 238024 46316 238076 46368
rect 106280 46248 106332 46300
rect 229836 46248 229888 46300
rect 244280 46248 244332 46300
rect 426532 46248 426584 46300
rect 40040 46180 40092 46232
rect 253480 46180 253532 46232
rect 3424 45500 3476 45552
rect 25504 45500 25556 45552
rect 48320 44888 48372 44940
rect 256056 44888 256108 44940
rect 31760 44820 31812 44872
rect 247684 44820 247736 44872
rect 269764 44820 269816 44872
rect 386420 44820 386472 44872
rect 240416 43528 240468 43580
rect 410524 43528 410576 43580
rect 52552 43460 52604 43512
rect 245016 43460 245068 43512
rect 27620 43392 27672 43444
rect 246396 43392 246448 43444
rect 338120 42168 338172 42220
rect 352012 42168 352064 42220
rect 262220 42100 262272 42152
rect 339500 42100 339552 42152
rect 53840 42032 53892 42084
rect 262864 42032 262916 42084
rect 349252 42032 349304 42084
rect 430672 42032 430724 42084
rect 340880 41352 340932 41404
rect 341524 41352 341576 41404
rect 427912 41352 427964 41404
rect 100760 40740 100812 40792
rect 235264 40740 235316 40792
rect 41420 40672 41472 40724
rect 265716 40672 265768 40724
rect 298100 40672 298152 40724
rect 338212 40672 338264 40724
rect 333980 39992 334032 40044
rect 334624 39992 334676 40044
rect 429292 39992 429344 40044
rect 110512 39380 110564 39432
rect 264336 39380 264388 39432
rect 27712 39312 27764 39364
rect 240784 39312 240836 39364
rect 255320 39312 255372 39364
rect 327816 39312 327868 39364
rect 35900 37952 35952 38004
rect 232596 37952 232648 38004
rect 324412 37952 324464 38004
rect 356060 37952 356112 38004
rect 24860 37884 24912 37936
rect 231216 37884 231268 37936
rect 248512 37884 248564 37936
rect 325056 37884 325108 37936
rect 356704 37884 356756 37936
rect 389180 37884 389232 37936
rect 337384 37204 337436 37256
rect 429200 37204 429252 37256
rect 336740 36864 336792 36916
rect 337384 36864 337436 36916
rect 266360 36524 266412 36576
rect 336188 36524 336240 36576
rect 103520 35232 103572 35284
rect 257620 35232 257672 35284
rect 320180 35232 320232 35284
rect 357440 35232 357492 35284
rect 34520 35164 34572 35216
rect 238300 35164 238352 35216
rect 241888 35164 241940 35216
rect 322296 35164 322348 35216
rect 340972 35164 341024 35216
rect 433616 35164 433668 35216
rect 22008 34416 22060 34468
rect 429384 34416 429436 34468
rect 3240 33736 3292 33788
rect 22008 33736 22060 33788
rect 45560 33736 45612 33788
rect 251824 33736 251876 33788
rect 349160 33056 349212 33108
rect 580172 33056 580224 33108
rect 174544 32444 174596 32496
rect 244280 32444 244332 32496
rect 55220 32376 55272 32428
rect 239496 32376 239548 32428
rect 316132 32444 316184 32496
rect 358820 32444 358872 32496
rect 320916 32376 320968 32428
rect 95240 31152 95292 31204
rect 236644 31152 236696 31204
rect 121460 31084 121512 31136
rect 264244 31084 264296 31136
rect 22100 31016 22152 31068
rect 251916 31016 251968 31068
rect 294144 31016 294196 31068
rect 367100 31016 367152 31068
rect 204904 29792 204956 29844
rect 283564 29792 283616 29844
rect 200764 29724 200816 29776
rect 114560 29656 114612 29708
rect 238208 29656 238260 29708
rect 59360 29588 59412 29640
rect 244924 29588 244976 29640
rect 288440 29588 288492 29640
rect 368480 29588 368532 29640
rect 196624 28908 196676 28960
rect 276112 28908 276164 28960
rect 276664 28908 276716 28960
rect 73160 28296 73212 28348
rect 253204 28296 253256 28348
rect 44272 28228 44324 28280
rect 231124 28228 231176 28280
rect 287704 28228 287756 28280
rect 369860 28228 369912 28280
rect 206284 26936 206336 26988
rect 29000 26868 29052 26920
rect 259000 26868 259052 26920
rect 259552 26868 259604 26920
rect 379520 26868 379572 26920
rect 33140 25508 33192 25560
rect 257528 25508 257580 25560
rect 289084 25508 289136 25560
rect 374000 25508 374052 25560
rect 252928 24216 252980 24268
rect 380992 24216 381044 24268
rect 36544 24148 36596 24200
rect 263600 24148 263652 24200
rect 11152 24080 11204 24132
rect 254676 24080 254728 24132
rect 115940 22788 115992 22840
rect 224224 22788 224276 22840
rect 26240 22720 26292 22772
rect 246488 22720 246540 22772
rect 245752 22652 245804 22704
rect 383660 22720 383712 22772
rect 203524 21496 203576 21548
rect 89720 21428 89772 21480
rect 261576 21428 261628 21480
rect 67640 21360 67692 21412
rect 243544 21360 243596 21412
rect 270500 21360 270552 21412
rect 375380 21360 375432 21412
rect 3424 20612 3476 20664
rect 29644 20612 29696 20664
rect 191104 20612 191156 20664
rect 267740 20612 267792 20664
rect 268384 20612 268436 20664
rect 493324 20612 493376 20664
rect 579988 20612 580040 20664
rect 84200 20000 84252 20052
rect 233884 20000 233936 20052
rect 77300 19932 77352 19984
rect 260196 19932 260248 19984
rect 273352 19932 273404 19984
rect 376760 19932 376812 19984
rect 263600 19252 263652 19304
rect 378140 19252 378192 19304
rect 195244 19184 195296 19236
rect 273352 19184 273404 19236
rect 82820 18640 82872 18692
rect 253296 18640 253348 18692
rect 70400 18572 70452 18624
rect 250444 18572 250496 18624
rect 180064 17212 180116 17264
rect 249800 17212 249852 17264
rect 382280 17212 382332 17264
rect 102140 15920 102192 15972
rect 262956 15920 263008 15972
rect 21824 15852 21876 15904
rect 238116 15852 238168 15904
rect 243544 15852 243596 15904
rect 385040 15852 385092 15904
rect 87512 14492 87564 14544
rect 257344 14492 257396 14544
rect 339500 14492 339552 14544
rect 391940 14492 391992 14544
rect 164424 14424 164476 14476
rect 350632 14424 350684 14476
rect 293224 13744 293276 13796
rect 406384 13744 406436 13796
rect 188344 13200 188396 13252
rect 261760 13200 261812 13252
rect 264428 13200 264480 13252
rect 80888 13132 80940 13184
rect 239404 13132 239456 13184
rect 94688 13064 94740 13116
rect 260104 13064 260156 13116
rect 283104 12384 283156 12436
rect 283564 12384 283616 12436
rect 411260 12384 411312 12436
rect 20168 11772 20220 11824
rect 232504 11772 232556 11824
rect 63408 11704 63460 11756
rect 281908 11704 281960 11756
rect 33140 10956 33192 11008
rect 34336 10956 34388 11008
rect 230480 10956 230532 11008
rect 258448 10888 258500 10940
rect 259368 10888 259420 10940
rect 5448 10276 5500 10328
rect 33140 10276 33192 10328
rect 78128 10276 78180 10328
rect 255964 10276 256016 10328
rect 259368 10276 259420 10328
rect 420920 10276 420972 10328
rect 186964 9596 187016 9648
rect 278044 9596 278096 9648
rect 278320 9596 278372 9648
rect 102232 8984 102284 9036
rect 261484 8984 261536 9036
rect 13544 8916 13596 8968
rect 229744 8916 229796 8968
rect 264980 8916 265032 8968
rect 418160 8916 418212 8968
rect 251272 8168 251324 8220
rect 252376 8168 252428 8220
rect 202144 7692 202196 7744
rect 256700 7692 256752 7744
rect 70308 7624 70360 7676
rect 246304 7624 246356 7676
rect 17040 7556 17092 7608
rect 236736 7556 236788 7608
rect 252376 7556 252428 7608
rect 307024 7624 307076 7676
rect 306748 7556 306800 7608
rect 362960 7556 363012 7608
rect 3424 6808 3476 6860
rect 15844 6808 15896 6860
rect 281908 6808 281960 6860
rect 371240 6808 371292 6860
rect 471244 6808 471296 6860
rect 580172 6808 580224 6860
rect 38568 6264 38620 6316
rect 136456 6264 136508 6316
rect 34428 6196 34480 6248
rect 132960 6196 133012 6248
rect 15200 6128 15252 6180
rect 265624 6128 265676 6180
rect 256700 5448 256752 5500
rect 257068 5448 257120 5500
rect 380900 5448 380952 5500
rect 184204 4904 184256 4956
rect 239128 4904 239180 4956
rect 91560 4836 91612 4888
rect 249064 4836 249116 4888
rect 63224 4768 63276 4820
rect 258724 4768 258776 4820
rect 349160 4224 349212 4276
rect 353300 4224 353352 4276
rect 239128 4088 239180 4140
rect 239312 4088 239364 4140
rect 269764 4088 269816 4140
rect 308404 4088 308456 4140
rect 322204 4088 322256 4140
rect 216036 4020 216088 4072
rect 242900 4020 242952 4072
rect 243544 4020 243596 4072
rect 125876 3612 125928 3664
rect 173900 3612 173952 3664
rect 35808 3544 35860 3596
rect 129372 3544 129424 3596
rect 244096 3544 244148 3596
rect 245108 3544 245160 3596
rect 276020 3544 276072 3596
rect 276756 3544 276808 3596
rect 292580 3544 292632 3596
rect 294052 3544 294104 3596
rect 316132 3544 316184 3596
rect 317328 3544 317380 3596
rect 322112 3544 322164 3596
rect 331220 3544 331272 3596
rect 346952 3544 347004 3596
rect 356704 3544 356756 3596
rect 27620 3476 27672 3528
rect 28540 3476 28592 3528
rect 44180 3476 44232 3528
rect 45100 3476 45152 3528
rect 52460 3476 52512 3528
rect 53380 3476 53432 3528
rect 64328 3476 64380 3528
rect 87604 3476 87656 3528
rect 102140 3476 102192 3528
rect 103336 3476 103388 3528
rect 103428 3476 103480 3528
rect 198096 3476 198148 3528
rect 267004 3476 267056 3528
rect 274824 3476 274876 3528
rect 289084 3476 289136 3528
rect 290188 3476 290240 3528
rect 295340 3476 295392 3528
rect 304356 3476 304408 3528
rect 305000 3476 305052 3528
rect 309048 3476 309100 3528
rect 309784 3476 309836 3528
rect 324320 3476 324372 3528
rect 325608 3476 325660 3528
rect 332600 3476 332652 3528
rect 333888 3476 333940 3528
rect 6460 3408 6512 3460
rect 15200 3408 15252 3460
rect 35992 3408 36044 3460
rect 214564 3408 214616 3460
rect 216128 3408 216180 3460
rect 285404 3408 285456 3460
rect 287704 3408 287756 3460
rect 332692 3408 332744 3460
rect 340144 3476 340196 3528
rect 340880 3476 340932 3528
rect 342168 3476 342220 3528
rect 350448 3476 350500 3528
rect 351920 3476 351972 3528
rect 99840 3340 99892 3392
rect 103428 3340 103480 3392
rect 331588 3340 331640 3392
rect 349160 3408 349212 3460
rect 351644 3408 351696 3460
rect 388444 3408 388496 3460
rect 267740 3272 267792 3324
rect 273352 3272 273404 3324
rect 1676 3204 1728 3256
rect 5448 3204 5500 3256
rect 299664 3136 299716 3188
rect 302240 3136 302292 3188
rect 233976 3000 234028 3052
rect 235816 3000 235868 3052
rect 279516 2932 279568 2984
rect 280252 2932 280304 2984
rect 109316 2048 109368 2100
rect 242164 2048 242216 2100
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 2832 632088 2834 632097
rect 2778 632023 2834 632032
rect 3436 595474 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 4804 632120 4856 632126
rect 4804 632062 4856 632068
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3424 595468 3476 595474
rect 3424 595410 3476 595416
rect 3424 582480 3476 582486
rect 3424 582422 3476 582428
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3436 553897 3464 582422
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 4816 538898 4844 632062
rect 6932 598262 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 698970 24348 703520
rect 24308 698964 24360 698970
rect 24308 698906 24360 698912
rect 11704 656940 11756 656946
rect 11704 656882 11756 656888
rect 6920 598256 6972 598262
rect 6920 598198 6972 598204
rect 11716 588606 11744 656882
rect 35164 605872 35216 605878
rect 35164 605814 35216 605820
rect 11704 588600 11756 588606
rect 11704 588542 11756 588548
rect 34244 568608 34296 568614
rect 34244 568550 34296 568556
rect 25504 565888 25556 565894
rect 25504 565830 25556 565836
rect 25516 544406 25544 565830
rect 25504 544400 25556 544406
rect 25504 544342 25556 544348
rect 4804 538892 4856 538898
rect 4804 538834 4856 538840
rect 3148 528556 3200 528562
rect 3148 528498 3200 528504
rect 3160 527921 3188 528498
rect 3146 527912 3202 527921
rect 3146 527847 3202 527856
rect 34152 525836 34204 525842
rect 34152 525778 34204 525784
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 7564 514820 7616 514826
rect 3424 514762 3476 514768
rect 7564 514762 7616 514768
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 3436 495446 3464 501735
rect 7576 500274 7604 514762
rect 7564 500268 7616 500274
rect 7564 500210 7616 500216
rect 3424 495440 3476 495446
rect 3424 495382 3476 495388
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 25504 474768 25556 474774
rect 25504 474710 25556 474716
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 4804 462596 4856 462602
rect 2780 462538 2832 462544
rect 4804 462538 4856 462544
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 3436 438598 3464 449511
rect 3424 438592 3476 438598
rect 3424 438534 3476 438540
rect 4816 438190 4844 462538
rect 25516 438938 25544 474710
rect 32954 458824 33010 458833
rect 32954 458759 33010 458768
rect 30288 455456 30340 455462
rect 30288 455398 30340 455404
rect 25504 438932 25556 438938
rect 25504 438874 25556 438880
rect 4804 438184 4856 438190
rect 4804 438126 4856 438132
rect 3424 429888 3476 429894
rect 3424 429830 3476 429836
rect 3436 410553 3464 429830
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3436 392630 3464 397423
rect 3424 392624 3476 392630
rect 3424 392566 3476 392572
rect 4804 388476 4856 388482
rect 4804 388418 4856 388424
rect 3240 372564 3292 372570
rect 3240 372506 3292 372512
rect 3252 371385 3280 372506
rect 3238 371376 3294 371385
rect 3238 371311 3294 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 4816 346322 4844 388418
rect 18604 380180 18656 380186
rect 18604 380122 18656 380128
rect 7564 352572 7616 352578
rect 7564 352514 7616 352520
rect 2780 346316 2832 346322
rect 2780 346258 2832 346264
rect 4804 346316 4856 346322
rect 4804 346258 4856 346264
rect 2792 345409 2820 346258
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 4804 328500 4856 328506
rect 4804 328442 4856 328448
rect 3240 319524 3292 319530
rect 3240 319466 3292 319472
rect 3252 319297 3280 319466
rect 3238 319288 3294 319297
rect 3238 319223 3294 319232
rect 3424 306264 3476 306270
rect 3422 306232 3424 306241
rect 3476 306232 3478 306241
rect 3422 306167 3478 306176
rect 4816 293214 4844 328442
rect 7576 306270 7604 352514
rect 18616 319530 18644 380122
rect 30300 358086 30328 455398
rect 32968 361554 32996 458759
rect 34164 442950 34192 525778
rect 34256 469198 34284 568550
rect 34336 547936 34388 547942
rect 34336 547878 34388 547884
rect 34244 469192 34296 469198
rect 34244 469134 34296 469140
rect 34348 447030 34376 547878
rect 35176 539578 35204 605814
rect 40052 590714 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 77944 703248 77996 703254
rect 77944 703190 77996 703196
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 76564 703044 76616 703050
rect 76564 702986 76616 702992
rect 68928 702500 68980 702506
rect 68928 702442 68980 702448
rect 62028 700324 62080 700330
rect 62028 700266 62080 700272
rect 54484 670744 54536 670750
rect 54484 670686 54536 670692
rect 52368 598256 52420 598262
rect 52368 598198 52420 598204
rect 52380 597582 52408 598198
rect 52368 597576 52420 597582
rect 52368 597518 52420 597524
rect 42800 595468 42852 595474
rect 42800 595410 42852 595416
rect 42812 594862 42840 595410
rect 42800 594856 42852 594862
rect 42800 594798 42852 594804
rect 44088 594856 44140 594862
rect 44088 594798 44140 594804
rect 40040 590708 40092 590714
rect 40040 590650 40092 590656
rect 39764 586628 39816 586634
rect 39764 586570 39816 586576
rect 37096 581324 37148 581330
rect 37096 581266 37148 581272
rect 35808 581120 35860 581126
rect 35808 581062 35860 581068
rect 35716 550656 35768 550662
rect 35716 550598 35768 550604
rect 35164 539572 35216 539578
rect 35164 539514 35216 539520
rect 35532 490612 35584 490618
rect 35532 490554 35584 490560
rect 34428 476128 34480 476134
rect 34428 476070 34480 476076
rect 34336 447024 34388 447030
rect 34336 446966 34388 446972
rect 34336 443692 34388 443698
rect 34336 443634 34388 443640
rect 33048 442944 33100 442950
rect 33048 442886 33100 442892
rect 34152 442944 34204 442950
rect 34152 442886 34204 442892
rect 32956 361548 33008 361554
rect 32956 361490 33008 361496
rect 30288 358080 30340 358086
rect 30288 358022 30340 358028
rect 33060 340814 33088 442886
rect 34244 383716 34296 383722
rect 34244 383658 34296 383664
rect 33048 340808 33100 340814
rect 33048 340750 33100 340756
rect 18604 319524 18656 319530
rect 18604 319466 18656 319472
rect 7564 306264 7616 306270
rect 7564 306206 7616 306212
rect 29642 298344 29698 298353
rect 29642 298279 29698 298288
rect 2780 293208 2832 293214
rect 2778 293176 2780 293185
rect 4804 293208 4856 293214
rect 2832 293176 2834 293185
rect 4804 293150 4856 293156
rect 2778 293111 2834 293120
rect 11704 292596 11756 292602
rect 11704 292538 11756 292544
rect 4068 291848 4120 291854
rect 4068 291790 4120 291796
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3146 241088 3202 241097
rect 3146 241023 3202 241032
rect 3160 240106 3188 241023
rect 3148 240100 3200 240106
rect 3148 240042 3200 240048
rect 3436 238746 3464 267135
rect 3424 238740 3476 238746
rect 3424 238682 3476 238688
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 214674 3372 214911
rect 3332 214668 3384 214674
rect 3332 214610 3384 214616
rect 3332 203584 3384 203590
rect 3332 203526 3384 203532
rect 3344 201929 3372 203526
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 4080 189106 4108 291790
rect 7564 264240 7616 264246
rect 7564 264182 7616 264188
rect 4804 222216 4856 222222
rect 4804 222158 4856 222164
rect 3516 189100 3568 189106
rect 3516 189042 3568 189048
rect 4068 189100 4120 189106
rect 4068 189042 4120 189048
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3528 180794 3556 189042
rect 3436 180766 3556 180794
rect 3436 162897 3464 180766
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 4816 97782 4844 222158
rect 7576 214674 7604 264182
rect 7564 214668 7616 214674
rect 7564 214610 7616 214616
rect 11716 189038 11744 292538
rect 22744 290488 22796 290494
rect 22744 290430 22796 290436
rect 15844 279472 15896 279478
rect 15844 279414 15896 279420
rect 11704 189032 11756 189038
rect 11704 188974 11756 188980
rect 14464 176792 14516 176798
rect 14464 176734 14516 176740
rect 14476 111790 14504 176734
rect 14464 111784 14516 111790
rect 14464 111726 14516 111732
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 11060 75200 11112 75206
rect 11060 75142 11112 75148
rect 9678 73808 9734 73817
rect 9678 73743 9734 73752
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 18 69592 74 69601
rect 18 69527 74 69536
rect 32 16574 60 69527
rect 6920 66904 6972 66910
rect 6920 66846 6972 66852
rect 4252 60036 4304 60042
rect 4252 59978 4304 59984
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 2780 55888 2832 55894
rect 2780 55830 2832 55836
rect 32 16546 152 16574
rect 124 354 152 16546
rect 2792 6914 2820 55830
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3240 33788 3292 33794
rect 3240 33730 3292 33736
rect 3252 32473 3280 33730
rect 3238 32464 3294 32473
rect 3238 32399 3294 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 2870 17232 2926 17241
rect 2870 17167 2926 17176
rect 2884 16574 2912 17167
rect 4264 16574 4292 59978
rect 6932 16574 6960 66846
rect 8298 36544 8354 36553
rect 8298 36479 8354 36488
rect 8312 16574 8340 36479
rect 2884 16546 3648 16574
rect 4264 16546 5304 16574
rect 6932 16546 7696 16574
rect 8312 16546 8800 16574
rect 2792 6886 2912 6914
rect 1676 3256 1728 3262
rect 1676 3198 1728 3204
rect 1688 480 1716 3198
rect 2884 480 2912 6886
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5276 480 5304 16546
rect 5448 10328 5500 10334
rect 5448 10270 5500 10276
rect 5460 3262 5488 10270
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 5448 3256 5500 3262
rect 5448 3198 5500 3204
rect 6472 480 6500 3402
rect 7668 480 7696 16546
rect 8772 480 8800 16546
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 73743
rect 11072 6914 11100 75142
rect 13820 57248 13872 57254
rect 13820 57190 13872 57196
rect 11152 24132 11204 24138
rect 11152 24074 11204 24080
rect 11164 16574 11192 24074
rect 13832 16574 13860 57190
rect 15200 54528 15252 54534
rect 15200 54470 15252 54476
rect 15212 16574 15240 54470
rect 11164 16546 11928 16574
rect 13832 16546 14320 16574
rect 15212 16546 15792 16574
rect 11072 6886 11192 6914
rect 11164 480 11192 6886
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13556 480 13584 8910
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15212 3466 15240 6122
rect 15764 3482 15792 16546
rect 15856 6866 15884 279414
rect 22008 268388 22060 268394
rect 22008 268330 22060 268336
rect 17224 257372 17276 257378
rect 17224 257314 17276 257320
rect 17236 137970 17264 257314
rect 17224 137964 17276 137970
rect 17224 137906 17276 137912
rect 17960 51740 18012 51746
rect 17960 51682 18012 51688
rect 17040 7608 17092 7614
rect 17040 7550 17092 7556
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15200 3460 15252 3466
rect 15764 3454 15976 3482
rect 15200 3402 15252 3408
rect 15948 480 15976 3454
rect 17052 480 17080 7550
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 51682
rect 19340 50380 19392 50386
rect 19340 50322 19392 50328
rect 19352 16574 19380 50322
rect 22020 34474 22048 268330
rect 22756 150414 22784 290430
rect 25504 176044 25556 176050
rect 25504 175986 25556 175992
rect 22744 150408 22796 150414
rect 22744 150350 22796 150356
rect 25516 45558 25544 175986
rect 25504 45552 25556 45558
rect 25504 45494 25556 45500
rect 27620 43444 27672 43450
rect 27620 43386 27672 43392
rect 23478 42120 23534 42129
rect 23478 42055 23534 42064
rect 22008 34468 22060 34474
rect 22008 34410 22060 34416
rect 22020 33794 22048 34410
rect 22008 33788 22060 33794
rect 22008 33730 22060 33736
rect 22100 31068 22152 31074
rect 22100 31010 22152 31016
rect 22112 16574 22140 31010
rect 23492 16574 23520 42055
rect 24860 37936 24912 37942
rect 24860 37878 24912 37884
rect 24872 16574 24900 37878
rect 26240 22772 26292 22778
rect 26240 22714 26292 22720
rect 19352 16546 19472 16574
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 19444 480 19472 16546
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20180 354 20208 11766
rect 21836 480 21864 15846
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 22714
rect 27632 3534 27660 43386
rect 27712 39364 27764 39370
rect 27712 39306 27764 39312
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27724 480 27752 39306
rect 29000 26920 29052 26926
rect 29000 26862 29052 26868
rect 29012 16574 29040 26862
rect 29656 20670 29684 298279
rect 33324 255264 33376 255270
rect 33324 255206 33376 255212
rect 33336 254590 33364 255206
rect 34256 254590 34284 383658
rect 34348 342922 34376 443634
rect 34336 342916 34388 342922
rect 34336 342858 34388 342864
rect 34336 294024 34388 294030
rect 34336 293966 34388 293972
rect 33324 254584 33376 254590
rect 33324 254526 33376 254532
rect 34244 254584 34296 254590
rect 34244 254526 34296 254532
rect 30380 53100 30432 53106
rect 30380 53042 30432 53048
rect 29644 20664 29696 20670
rect 29644 20606 29696 20612
rect 30392 16574 30420 53042
rect 31760 44872 31812 44878
rect 31760 44814 31812 44820
rect 31772 16574 31800 44814
rect 33140 25560 33192 25566
rect 33140 25502 33192 25508
rect 33152 16574 33180 25502
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3470
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33140 11008 33192 11014
rect 33140 10950 33192 10956
rect 33152 10334 33180 10950
rect 33140 10328 33192 10334
rect 33140 10270 33192 10276
rect 33612 480 33640 16546
rect 34348 11014 34376 293966
rect 34336 11008 34388 11014
rect 34336 10950 34388 10956
rect 34440 6254 34468 476070
rect 35544 387938 35572 490554
rect 35624 475380 35676 475386
rect 35624 475322 35676 475328
rect 35532 387932 35584 387938
rect 35532 387874 35584 387880
rect 35636 380254 35664 475322
rect 35728 451217 35756 550598
rect 35820 487150 35848 581062
rect 36544 554804 36596 554810
rect 36544 554746 36596 554752
rect 35808 487144 35860 487150
rect 35808 487086 35860 487092
rect 36556 455394 36584 554746
rect 37108 490618 37136 581266
rect 38568 575544 38620 575550
rect 38568 575486 38620 575492
rect 37188 536104 37240 536110
rect 37188 536046 37240 536052
rect 37096 490612 37148 490618
rect 37096 490554 37148 490560
rect 37096 483064 37148 483070
rect 37096 483006 37148 483012
rect 36544 455388 36596 455394
rect 36544 455330 36596 455336
rect 35714 451208 35770 451217
rect 35714 451143 35770 451152
rect 37004 445052 37056 445058
rect 37004 444994 37056 445000
rect 36636 389156 36688 389162
rect 36636 389098 36688 389104
rect 36648 388482 36676 389098
rect 36636 388476 36688 388482
rect 36636 388418 36688 388424
rect 35716 387932 35768 387938
rect 35716 387874 35768 387880
rect 35624 380248 35676 380254
rect 35624 380190 35676 380196
rect 35728 257378 35756 387874
rect 35808 382288 35860 382294
rect 35808 382230 35860 382236
rect 35716 257372 35768 257378
rect 35716 257314 35768 257320
rect 34520 35216 34572 35222
rect 34520 35158 34572 35164
rect 34428 6248 34480 6254
rect 34428 6190 34480 6196
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 35158
rect 35820 3602 35848 382230
rect 36544 361616 36596 361622
rect 36544 361558 36596 361564
rect 35900 38004 35952 38010
rect 35900 37946 35952 37952
rect 35912 16574 35940 37946
rect 36556 24206 36584 361558
rect 37016 358766 37044 444994
rect 37108 389162 37136 483006
rect 37200 437306 37228 536046
rect 38476 492040 38528 492046
rect 38476 491982 38528 491988
rect 37188 437300 37240 437306
rect 37188 437242 37240 437248
rect 38488 395350 38516 491982
rect 38476 395344 38528 395350
rect 38476 395286 38528 395292
rect 37096 389156 37148 389162
rect 37096 389098 37148 389104
rect 37188 365696 37240 365702
rect 37188 365638 37240 365644
rect 37004 358760 37056 358766
rect 37004 358702 37056 358708
rect 37200 240106 37228 365638
rect 37188 240100 37240 240106
rect 37188 240042 37240 240048
rect 37200 239426 37228 240042
rect 37188 239420 37240 239426
rect 37188 239362 37240 239368
rect 37280 76560 37332 76566
rect 37280 76502 37332 76508
rect 36544 24200 36596 24206
rect 36544 24142 36596 24148
rect 37292 16574 37320 76502
rect 35912 16546 36768 16574
rect 37292 16546 38424 16574
rect 35808 3596 35860 3602
rect 35808 3538 35860 3544
rect 35992 3460 36044 3466
rect 35992 3402 36044 3408
rect 36004 480 36032 3402
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 38580 6322 38608 575486
rect 39672 526448 39724 526454
rect 39672 526390 39724 526396
rect 39684 431934 39712 526390
rect 39776 495582 39804 586570
rect 42616 586560 42668 586566
rect 42616 586502 42668 586508
rect 41144 585200 41196 585206
rect 41144 585142 41196 585148
rect 39948 580304 40000 580310
rect 39948 580246 40000 580252
rect 39856 534744 39908 534750
rect 39856 534686 39908 534692
rect 39764 495576 39816 495582
rect 39764 495518 39816 495524
rect 39672 431928 39724 431934
rect 39672 431870 39724 431876
rect 39684 336666 39712 431870
rect 39776 399498 39804 495518
rect 39868 437374 39896 534686
rect 39960 480962 39988 580246
rect 41052 529304 41104 529310
rect 41052 529246 41104 529252
rect 39948 480956 40000 480962
rect 39948 480898 40000 480904
rect 39856 437368 39908 437374
rect 39856 437310 39908 437316
rect 39764 399492 39816 399498
rect 39764 399434 39816 399440
rect 39856 396840 39908 396846
rect 39856 396782 39908 396788
rect 39764 393440 39816 393446
rect 39764 393382 39816 393388
rect 39672 336660 39724 336666
rect 39672 336602 39724 336608
rect 39776 271674 39804 393382
rect 39868 273465 39896 396782
rect 39960 389094 39988 480898
rect 40960 459604 41012 459610
rect 40960 459546 41012 459552
rect 39948 389088 40000 389094
rect 39948 389030 40000 389036
rect 40972 365702 41000 459546
rect 41064 434722 41092 529246
rect 41156 495514 41184 585142
rect 41328 583772 41380 583778
rect 41328 583714 41380 583720
rect 41236 558952 41288 558958
rect 41236 558894 41288 558900
rect 41144 495508 41196 495514
rect 41144 495450 41196 495456
rect 41052 434716 41104 434722
rect 41052 434658 41104 434664
rect 41156 399566 41184 495450
rect 41248 460222 41276 558894
rect 41340 491434 41368 583714
rect 42524 529236 42576 529242
rect 42524 529178 42576 529184
rect 41328 491428 41380 491434
rect 41328 491370 41380 491376
rect 41236 460216 41288 460222
rect 41236 460158 41288 460164
rect 41248 459610 41276 460158
rect 41236 459604 41288 459610
rect 41236 459546 41288 459552
rect 41236 434716 41288 434722
rect 41236 434658 41288 434664
rect 41144 399560 41196 399566
rect 41144 399502 41196 399508
rect 40960 365696 41012 365702
rect 40960 365638 41012 365644
rect 41144 342916 41196 342922
rect 41144 342858 41196 342864
rect 39854 273456 39910 273465
rect 39854 273391 39910 273400
rect 39776 271646 39896 271674
rect 39868 269074 39896 271646
rect 39948 269136 40000 269142
rect 39948 269078 40000 269084
rect 39856 269068 39908 269074
rect 39856 269010 39908 269016
rect 39868 268394 39896 269010
rect 39856 268388 39908 268394
rect 39856 268330 39908 268336
rect 39960 185638 39988 269078
rect 41156 267034 41184 342858
rect 41248 333985 41276 434658
rect 41340 392601 41368 491370
rect 42536 434722 42564 529178
rect 42628 495650 42656 586502
rect 43996 582616 44048 582622
rect 43996 582558 44048 582564
rect 42708 556232 42760 556238
rect 42708 556174 42760 556180
rect 42616 495644 42668 495650
rect 42616 495586 42668 495592
rect 42524 434716 42576 434722
rect 42524 434658 42576 434664
rect 41326 392592 41382 392601
rect 41326 392527 41382 392536
rect 41328 385688 41380 385694
rect 41328 385630 41380 385636
rect 41234 333976 41290 333985
rect 41234 333911 41290 333920
rect 41236 274712 41288 274718
rect 41236 274654 41288 274660
rect 41144 267028 41196 267034
rect 41144 266970 41196 266976
rect 41248 217394 41276 274654
rect 41340 263022 41368 385630
rect 42536 339454 42564 434658
rect 42628 396778 42656 495586
rect 42720 456754 42748 556174
rect 43812 537600 43864 537606
rect 43812 537542 43864 537548
rect 43720 493332 43772 493338
rect 43720 493274 43772 493280
rect 42708 456748 42760 456754
rect 42708 456690 42760 456696
rect 42706 454744 42762 454753
rect 42706 454679 42762 454688
rect 42616 396772 42668 396778
rect 42616 396714 42668 396720
rect 42720 356726 42748 454679
rect 43732 395418 43760 493274
rect 43824 440910 43852 537542
rect 44008 492046 44036 582558
rect 43996 492040 44048 492046
rect 43996 491982 44048 491988
rect 43904 491972 43956 491978
rect 43904 491914 43956 491920
rect 43812 440904 43864 440910
rect 43812 440846 43864 440852
rect 43916 395486 43944 491914
rect 44100 484362 44128 594798
rect 48228 590708 48280 590714
rect 48228 590650 48280 590656
rect 45376 583840 45428 583846
rect 45376 583782 45428 583788
rect 45388 491978 45416 583782
rect 46664 582548 46716 582554
rect 46664 582490 46716 582496
rect 45468 536172 45520 536178
rect 45468 536114 45520 536120
rect 45376 491972 45428 491978
rect 45376 491914 45428 491920
rect 45376 490680 45428 490686
rect 45376 490622 45428 490628
rect 44088 484356 44140 484362
rect 44088 484298 44140 484304
rect 44088 474020 44140 474026
rect 44088 473962 44140 473968
rect 43996 398132 44048 398138
rect 43996 398074 44048 398080
rect 43904 395480 43956 395486
rect 43904 395422 43956 395428
rect 43720 395412 43772 395418
rect 43720 395354 43772 395360
rect 42984 389224 43036 389230
rect 42984 389166 43036 389172
rect 43444 389224 43496 389230
rect 43444 389166 43496 389172
rect 42996 389094 43024 389166
rect 42984 389088 43036 389094
rect 42984 389030 43036 389036
rect 42800 380860 42852 380866
rect 42800 380802 42852 380808
rect 42812 380186 42840 380802
rect 42800 380180 42852 380186
rect 42800 380122 42852 380128
rect 42708 356720 42760 356726
rect 42708 356662 42760 356668
rect 42524 339448 42576 339454
rect 42524 339390 42576 339396
rect 42720 279478 42748 356662
rect 42708 279472 42760 279478
rect 42708 279414 42760 279420
rect 41328 263016 41380 263022
rect 41328 262958 41380 262964
rect 41328 262880 41380 262886
rect 41328 262822 41380 262828
rect 41236 217388 41288 217394
rect 41236 217330 41288 217336
rect 39948 185632 40000 185638
rect 39948 185574 40000 185580
rect 41340 181393 41368 262822
rect 43456 249082 43484 389166
rect 43902 383208 43958 383217
rect 43902 383143 43958 383152
rect 43536 358760 43588 358766
rect 43536 358702 43588 358708
rect 43548 345710 43576 358702
rect 43536 345704 43588 345710
rect 43536 345646 43588 345652
rect 43916 339522 43944 383143
rect 43904 339516 43956 339522
rect 43904 339458 43956 339464
rect 44008 338094 44036 398074
rect 44100 380866 44128 473962
rect 44824 456748 44876 456754
rect 44824 456690 44876 456696
rect 44088 380860 44140 380866
rect 44088 380802 44140 380808
rect 44836 360874 44864 456690
rect 45284 434036 45336 434042
rect 45284 433978 45336 433984
rect 44824 360868 44876 360874
rect 44824 360810 44876 360816
rect 45296 339697 45324 433978
rect 45388 394058 45416 490622
rect 45480 437170 45508 536114
rect 46676 490686 46704 582490
rect 48044 564528 48096 564534
rect 48044 564470 48096 564476
rect 46754 537432 46810 537441
rect 46754 537367 46810 537376
rect 46664 490680 46716 490686
rect 46664 490622 46716 490628
rect 46664 469872 46716 469878
rect 46664 469814 46716 469820
rect 45468 437164 45520 437170
rect 45468 437106 45520 437112
rect 45376 394052 45428 394058
rect 45376 393994 45428 394000
rect 46572 393984 46624 393990
rect 46572 393926 46624 393932
rect 45468 360868 45520 360874
rect 45468 360810 45520 360816
rect 45282 339688 45338 339697
rect 45282 339623 45338 339632
rect 43996 338088 44048 338094
rect 43996 338030 44048 338036
rect 45376 280220 45428 280226
rect 45376 280162 45428 280168
rect 44088 255332 44140 255338
rect 44088 255274 44140 255280
rect 43444 249076 43496 249082
rect 43444 249018 43496 249024
rect 44100 184210 44128 255274
rect 45388 210458 45416 280162
rect 45480 253910 45508 360810
rect 46584 335306 46612 393926
rect 46676 375358 46704 469814
rect 46768 439006 46796 537367
rect 46848 534812 46900 534818
rect 46848 534754 46900 534760
rect 46756 439000 46808 439006
rect 46756 438942 46808 438948
rect 46664 375352 46716 375358
rect 46664 375294 46716 375300
rect 46768 339386 46796 438942
rect 46860 436014 46888 534754
rect 47952 532024 48004 532030
rect 47952 531966 48004 531972
rect 47964 437442 47992 531966
rect 48056 465050 48084 564470
rect 48136 556300 48188 556306
rect 48136 556242 48188 556248
rect 48044 465044 48096 465050
rect 48044 464986 48096 464992
rect 48044 458244 48096 458250
rect 48044 458186 48096 458192
rect 47952 437436 48004 437442
rect 47952 437378 48004 437384
rect 46848 436008 46900 436014
rect 46848 435950 46900 435956
rect 47952 387320 48004 387326
rect 47952 387262 48004 387268
rect 46848 349104 46900 349110
rect 46848 349046 46900 349052
rect 46756 339380 46808 339386
rect 46756 339322 46808 339328
rect 46572 335300 46624 335306
rect 46572 335242 46624 335248
rect 45468 253904 45520 253910
rect 45468 253846 45520 253852
rect 46860 234598 46888 349046
rect 47964 336462 47992 387262
rect 48056 363662 48084 458186
rect 48148 456754 48176 556242
rect 48240 487898 48268 590650
rect 52276 585336 52328 585342
rect 52276 585278 52328 585284
rect 50894 583944 50950 583953
rect 50894 583879 50950 583888
rect 50344 581256 50396 581262
rect 50344 581198 50396 581204
rect 49516 572008 49568 572014
rect 49516 571950 49568 571956
rect 49332 532160 49384 532166
rect 49332 532102 49384 532108
rect 48228 487892 48280 487898
rect 48228 487834 48280 487840
rect 48228 462324 48280 462330
rect 48228 462266 48280 462272
rect 48136 456748 48188 456754
rect 48136 456690 48188 456696
rect 48134 446448 48190 446457
rect 48134 446383 48190 446392
rect 48044 363656 48096 363662
rect 48044 363598 48096 363604
rect 48056 363118 48084 363598
rect 48044 363112 48096 363118
rect 48044 363054 48096 363060
rect 48148 349110 48176 446383
rect 48240 367062 48268 462266
rect 49344 434586 49372 532102
rect 49528 473346 49556 571950
rect 49608 542428 49660 542434
rect 49608 542370 49660 542376
rect 49516 473340 49568 473346
rect 49516 473282 49568 473288
rect 49422 449984 49478 449993
rect 49422 449919 49478 449928
rect 49332 434580 49384 434586
rect 49332 434522 49384 434528
rect 48228 367056 48280 367062
rect 48228 366998 48280 367004
rect 48228 363112 48280 363118
rect 48228 363054 48280 363060
rect 48136 349104 48188 349110
rect 48136 349046 48188 349052
rect 48148 348430 48176 349046
rect 48136 348424 48188 348430
rect 48136 348366 48188 348372
rect 47952 336456 48004 336462
rect 47952 336398 48004 336404
rect 48136 329112 48188 329118
rect 48136 329054 48188 329060
rect 48148 328506 48176 329054
rect 48136 328500 48188 328506
rect 48136 328442 48188 328448
rect 48044 277432 48096 277438
rect 48044 277374 48096 277380
rect 47308 253904 47360 253910
rect 47308 253846 47360 253852
rect 47320 252618 47348 253846
rect 46940 252612 46992 252618
rect 46940 252554 46992 252560
rect 47308 252612 47360 252618
rect 47308 252554 47360 252560
rect 46848 234592 46900 234598
rect 46848 234534 46900 234540
rect 45376 210452 45428 210458
rect 45376 210394 45428 210400
rect 44088 184204 44140 184210
rect 44088 184146 44140 184152
rect 41326 181384 41382 181393
rect 41326 181319 41382 181328
rect 46952 85542 46980 252554
rect 48056 220114 48084 277374
rect 48148 242894 48176 328442
rect 48240 264926 48268 363054
rect 49436 350606 49464 449919
rect 49620 442882 49648 542370
rect 50356 483070 50384 581198
rect 50712 496120 50764 496126
rect 50712 496062 50764 496068
rect 50344 483064 50396 483070
rect 50344 483006 50396 483012
rect 50344 465044 50396 465050
rect 50344 464986 50396 464992
rect 49608 442876 49660 442882
rect 49608 442818 49660 442824
rect 49516 438184 49568 438190
rect 49516 438126 49568 438132
rect 49424 350600 49476 350606
rect 49424 350542 49476 350548
rect 49528 333946 49556 438126
rect 49608 434580 49660 434586
rect 49608 434522 49660 434528
rect 49620 434042 49648 434522
rect 49608 434036 49660 434042
rect 49608 433978 49660 433984
rect 49608 390720 49660 390726
rect 49608 390662 49660 390668
rect 49516 333940 49568 333946
rect 49516 333882 49568 333888
rect 49424 284368 49476 284374
rect 49424 284310 49476 284316
rect 48228 264920 48280 264926
rect 48228 264862 48280 264868
rect 48240 264246 48268 264862
rect 48228 264240 48280 264246
rect 48228 264182 48280 264188
rect 48228 260908 48280 260914
rect 48228 260850 48280 260856
rect 48136 242888 48188 242894
rect 48136 242830 48188 242836
rect 48240 229770 48268 260850
rect 48228 229764 48280 229770
rect 48228 229706 48280 229712
rect 48044 220108 48096 220114
rect 48044 220050 48096 220056
rect 49436 195362 49464 284310
rect 49620 284306 49648 390662
rect 50356 370598 50384 464986
rect 50724 439550 50752 496062
rect 50908 489914 50936 583879
rect 52184 574116 52236 574122
rect 52184 574058 52236 574064
rect 50988 537532 51040 537538
rect 50988 537474 51040 537480
rect 50816 489886 50936 489914
rect 50816 487830 50844 489886
rect 50804 487824 50856 487830
rect 50804 487766 50856 487772
rect 50712 439544 50764 439550
rect 50712 439486 50764 439492
rect 50816 389298 50844 487766
rect 51000 441614 51028 537474
rect 52000 532092 52052 532098
rect 52000 532034 52052 532040
rect 51908 492856 51960 492862
rect 51908 492798 51960 492804
rect 51080 475448 51132 475454
rect 51080 475390 51132 475396
rect 51092 474026 51120 475390
rect 51080 474020 51132 474026
rect 51080 473962 51132 473968
rect 50908 441586 51028 441614
rect 50908 438802 50936 441586
rect 50896 438796 50948 438802
rect 50896 438738 50948 438744
rect 50804 389292 50856 389298
rect 50804 389234 50856 389240
rect 50344 370592 50396 370598
rect 50344 370534 50396 370540
rect 50804 370524 50856 370530
rect 50804 370466 50856 370472
rect 50712 339380 50764 339386
rect 50712 339322 50764 339328
rect 50724 338162 50752 339322
rect 50712 338156 50764 338162
rect 50712 338098 50764 338104
rect 49608 284300 49660 284306
rect 49608 284242 49660 284248
rect 49516 274780 49568 274786
rect 49516 274722 49568 274728
rect 49528 200938 49556 274722
rect 50724 246945 50752 338098
rect 50816 335238 50844 370466
rect 50908 337414 50936 438738
rect 50988 395480 51040 395486
rect 50988 395422 51040 395428
rect 51000 394738 51028 395422
rect 50988 394732 51040 394738
rect 50988 394674 51040 394680
rect 50896 337408 50948 337414
rect 50896 337350 50948 337356
rect 50804 335232 50856 335238
rect 50804 335174 50856 335180
rect 51000 292618 51028 394674
rect 51920 387161 51948 492798
rect 52012 438734 52040 532034
rect 52196 475454 52224 574058
rect 52288 492862 52316 585278
rect 52276 492856 52328 492862
rect 52276 492798 52328 492804
rect 52380 491434 52408 597518
rect 53472 585268 53524 585274
rect 53472 585210 53524 585216
rect 53104 579692 53156 579698
rect 53104 579634 53156 579640
rect 53116 538218 53144 579634
rect 53104 538212 53156 538218
rect 53104 538154 53156 538160
rect 53484 493338 53512 585210
rect 53748 583976 53800 583982
rect 53748 583918 53800 583924
rect 53564 560992 53616 560998
rect 53564 560934 53616 560940
rect 53472 493332 53524 493338
rect 53472 493274 53524 493280
rect 52368 491428 52420 491434
rect 52368 491370 52420 491376
rect 52380 489914 52408 491370
rect 52288 489886 52408 489914
rect 52184 475448 52236 475454
rect 52184 475390 52236 475396
rect 52092 451988 52144 451994
rect 52092 451930 52144 451936
rect 52000 438728 52052 438734
rect 52000 438670 52052 438676
rect 52012 438190 52040 438670
rect 52000 438184 52052 438190
rect 52000 438126 52052 438132
rect 51906 387152 51962 387161
rect 51906 387087 51962 387096
rect 52104 355366 52132 451930
rect 52184 389836 52236 389842
rect 52184 389778 52236 389784
rect 52092 355360 52144 355366
rect 52092 355302 52144 355308
rect 51184 292670 51212 292701
rect 51172 292664 51224 292670
rect 51000 292612 51172 292618
rect 51000 292606 51224 292612
rect 51000 292590 51212 292606
rect 51080 292528 51132 292534
rect 51080 292470 51132 292476
rect 51092 291854 51120 292470
rect 51080 291848 51132 291854
rect 51080 291790 51132 291796
rect 50988 288448 51040 288454
rect 50988 288390 51040 288396
rect 50804 262268 50856 262274
rect 50804 262210 50856 262216
rect 50710 246936 50766 246945
rect 50710 246871 50766 246880
rect 49516 200932 49568 200938
rect 49516 200874 49568 200880
rect 50816 198150 50844 262210
rect 50896 249824 50948 249830
rect 50896 249766 50948 249772
rect 50908 209098 50936 249766
rect 50896 209092 50948 209098
rect 50896 209034 50948 209040
rect 50804 198144 50856 198150
rect 50804 198086 50856 198092
rect 49424 195356 49476 195362
rect 49424 195298 49476 195304
rect 51000 191214 51028 288390
rect 51184 277394 51212 292590
rect 52196 292534 52224 389778
rect 52288 388006 52316 489886
rect 53288 484424 53340 484430
rect 53288 484366 53340 484372
rect 52460 463004 52512 463010
rect 52460 462946 52512 462952
rect 52472 462330 52500 462946
rect 52460 462324 52512 462330
rect 52460 462266 52512 462272
rect 52460 456884 52512 456890
rect 52460 456826 52512 456832
rect 53196 456884 53248 456890
rect 53196 456826 53248 456832
rect 52472 456754 52500 456826
rect 52460 456748 52512 456754
rect 52460 456690 52512 456696
rect 52460 438184 52512 438190
rect 52460 438126 52512 438132
rect 52472 437306 52500 438126
rect 52460 437300 52512 437306
rect 52460 437242 52512 437248
rect 53104 437300 53156 437306
rect 53104 437242 53156 437248
rect 52276 388000 52328 388006
rect 52276 387942 52328 387948
rect 52184 292528 52236 292534
rect 52184 292470 52236 292476
rect 51092 277366 51212 277394
rect 50988 191208 51040 191214
rect 50988 191150 51040 191156
rect 46940 85536 46992 85542
rect 46940 85478 46992 85484
rect 49698 72448 49754 72457
rect 49698 72383 49754 72392
rect 46940 65612 46992 65618
rect 46940 65554 46992 65560
rect 44180 47592 44232 47598
rect 44180 47534 44232 47540
rect 40040 46232 40092 46238
rect 40040 46174 40092 46180
rect 38658 32464 38714 32473
rect 38658 32399 38714 32408
rect 38672 16574 38700 32399
rect 40052 16574 40080 46174
rect 41420 40724 41472 40730
rect 41420 40666 41472 40672
rect 41432 16574 41460 40666
rect 42798 26888 42854 26897
rect 42798 26823 42854 26832
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 38568 6316 38620 6322
rect 38568 6258 38620 6264
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 26823
rect 44192 3534 44220 47534
rect 45560 33788 45612 33794
rect 45560 33730 45612 33736
rect 44272 28280 44324 28286
rect 44272 28222 44324 28228
rect 44180 3528 44232 3534
rect 44180 3470 44232 3476
rect 44284 480 44312 28222
rect 45572 16574 45600 33730
rect 46952 16574 46980 65554
rect 48320 44940 48372 44946
rect 48320 44882 48372 44888
rect 48332 16574 48360 44882
rect 49712 16574 49740 72383
rect 51092 59362 51120 277366
rect 52288 266354 52316 387942
rect 52368 387252 52420 387258
rect 52368 387194 52420 387200
rect 52380 387161 52408 387194
rect 52366 387152 52422 387161
rect 52366 387087 52422 387096
rect 52368 385076 52420 385082
rect 52368 385018 52420 385024
rect 52276 266348 52328 266354
rect 52276 266290 52328 266296
rect 52184 264988 52236 264994
rect 52184 264930 52236 264936
rect 52196 232762 52224 264930
rect 52276 258120 52328 258126
rect 52276 258062 52328 258068
rect 52184 232756 52236 232762
rect 52184 232698 52236 232704
rect 52288 185774 52316 258062
rect 52380 237318 52408 385018
rect 53116 338065 53144 437242
rect 53208 359514 53236 456826
rect 53300 391270 53328 484366
rect 53576 463010 53604 560934
rect 53656 534880 53708 534886
rect 53656 534822 53708 534828
rect 53564 463004 53616 463010
rect 53564 462946 53616 462952
rect 53668 437306 53696 534822
rect 53760 482905 53788 583918
rect 54496 538966 54524 670686
rect 56416 587920 56468 587926
rect 56416 587862 56468 587868
rect 55036 572076 55088 572082
rect 55036 572018 55088 572024
rect 54944 552084 54996 552090
rect 54944 552026 54996 552032
rect 54484 538960 54536 538966
rect 54484 538902 54536 538908
rect 54852 529372 54904 529378
rect 54852 529314 54904 529320
rect 53746 482896 53802 482905
rect 53746 482831 53802 482840
rect 54208 460284 54260 460290
rect 54208 460226 54260 460232
rect 54220 458250 54248 460226
rect 54208 458244 54260 458250
rect 54208 458186 54260 458192
rect 53656 437300 53708 437306
rect 53656 437242 53708 437248
rect 54864 437238 54892 529314
rect 54956 453354 54984 552026
rect 55048 472666 55076 572018
rect 55128 560312 55180 560318
rect 55128 560254 55180 560260
rect 55036 472660 55088 472666
rect 55036 472602 55088 472608
rect 54944 453348 54996 453354
rect 54944 453290 54996 453296
rect 54956 451994 54984 453290
rect 54944 451988 54996 451994
rect 54944 451930 54996 451936
rect 54852 437232 54904 437238
rect 54852 437174 54904 437180
rect 53288 391264 53340 391270
rect 53288 391206 53340 391212
rect 53748 389292 53800 389298
rect 53748 389234 53800 389240
rect 53564 385756 53616 385762
rect 53564 385698 53616 385704
rect 53196 359508 53248 359514
rect 53196 359450 53248 359456
rect 53102 338056 53158 338065
rect 53102 337991 53158 338000
rect 53576 336530 53604 385698
rect 53656 359508 53708 359514
rect 53656 359450 53708 359456
rect 53564 336524 53616 336530
rect 53564 336466 53616 336472
rect 53564 276072 53616 276078
rect 53564 276014 53616 276020
rect 52460 257372 52512 257378
rect 52460 257314 52512 257320
rect 52472 256766 52500 257314
rect 52460 256760 52512 256766
rect 52460 256702 52512 256708
rect 53472 256760 53524 256766
rect 53472 256702 53524 256708
rect 52368 237312 52420 237318
rect 52368 237254 52420 237260
rect 53484 191049 53512 256702
rect 53576 192642 53604 276014
rect 53668 234530 53696 359450
rect 53760 255270 53788 389234
rect 54942 386608 54998 386617
rect 54942 386543 54998 386552
rect 54956 386510 54984 386543
rect 54944 386504 54996 386510
rect 54944 386446 54996 386452
rect 53840 350600 53892 350606
rect 53840 350542 53892 350548
rect 53852 349858 53880 350542
rect 53840 349852 53892 349858
rect 53840 349794 53892 349800
rect 54956 294778 54984 386446
rect 55048 376718 55076 472602
rect 55140 460290 55168 560254
rect 56324 535492 56376 535498
rect 56324 535434 56376 535440
rect 56232 490748 56284 490754
rect 56232 490690 56284 490696
rect 55128 460284 55180 460290
rect 55128 460226 55180 460232
rect 55128 453416 55180 453422
rect 55128 453358 55180 453364
rect 55036 376712 55088 376718
rect 55036 376654 55088 376660
rect 55036 376032 55088 376038
rect 55036 375974 55088 375980
rect 55048 336598 55076 375974
rect 55140 356046 55168 453358
rect 56244 440978 56272 490690
rect 56336 455326 56364 535434
rect 56428 492726 56456 587862
rect 59176 586696 59228 586702
rect 59176 586638 59228 586644
rect 57796 584044 57848 584050
rect 57796 583986 57848 583992
rect 57702 583808 57758 583817
rect 57702 583743 57758 583752
rect 56508 563100 56560 563106
rect 56508 563042 56560 563048
rect 56416 492720 56468 492726
rect 56416 492662 56468 492668
rect 56324 455320 56376 455326
rect 56324 455262 56376 455268
rect 56232 440972 56284 440978
rect 56232 440914 56284 440920
rect 56324 438252 56376 438258
rect 56324 438194 56376 438200
rect 56336 437170 56364 438194
rect 55864 437164 55916 437170
rect 55864 437106 55916 437112
rect 56324 437164 56376 437170
rect 56324 437106 56376 437112
rect 55128 356040 55180 356046
rect 55128 355982 55180 355988
rect 55128 349852 55180 349858
rect 55128 349794 55180 349800
rect 55036 336592 55088 336598
rect 55036 336534 55088 336540
rect 54944 294772 54996 294778
rect 54944 294714 54996 294720
rect 55036 269204 55088 269210
rect 55036 269146 55088 269152
rect 53840 263016 53892 263022
rect 53840 262958 53892 262964
rect 53852 262342 53880 262958
rect 53840 262336 53892 262342
rect 53840 262278 53892 262284
rect 54852 262336 54904 262342
rect 54852 262278 54904 262284
rect 53748 255264 53800 255270
rect 53748 255206 53800 255212
rect 53748 249892 53800 249898
rect 53748 249834 53800 249840
rect 53656 234524 53708 234530
rect 53656 234466 53708 234472
rect 53564 192636 53616 192642
rect 53564 192578 53616 192584
rect 53470 191040 53526 191049
rect 53470 190975 53526 190984
rect 52276 185768 52328 185774
rect 52276 185710 52328 185716
rect 53760 181490 53788 249834
rect 54864 215966 54892 262278
rect 54944 251252 54996 251258
rect 54944 251194 54996 251200
rect 54852 215960 54904 215966
rect 54852 215902 54904 215908
rect 54956 188358 54984 251194
rect 55048 205086 55076 269146
rect 55140 233238 55168 349794
rect 55876 337890 55904 437106
rect 56428 396914 56456 492662
rect 56520 463690 56548 563042
rect 57612 554872 57664 554878
rect 57612 554814 57664 554820
rect 57624 536246 57652 554814
rect 57612 536240 57664 536246
rect 57612 536182 57664 536188
rect 57624 535498 57652 536182
rect 57612 535492 57664 535498
rect 57612 535434 57664 535440
rect 57716 493406 57744 583743
rect 57704 493400 57756 493406
rect 57702 493368 57704 493377
rect 57756 493368 57758 493377
rect 57702 493303 57758 493312
rect 57244 487892 57296 487898
rect 57244 487834 57296 487840
rect 57256 487218 57284 487834
rect 56600 487212 56652 487218
rect 56600 487154 56652 487160
rect 57244 487212 57296 487218
rect 57244 487154 57296 487160
rect 56508 463684 56560 463690
rect 56508 463626 56560 463632
rect 56508 455320 56560 455326
rect 56508 455262 56560 455268
rect 56520 454714 56548 455262
rect 56508 454708 56560 454714
rect 56508 454650 56560 454656
rect 56416 396908 56468 396914
rect 56416 396850 56468 396856
rect 56416 392692 56468 392698
rect 56416 392634 56468 392640
rect 56324 345092 56376 345098
rect 56324 345034 56376 345040
rect 55864 337884 55916 337890
rect 55864 337826 55916 337832
rect 56336 300121 56364 345034
rect 56428 337958 56456 392634
rect 56520 358766 56548 454650
rect 56612 387841 56640 487154
rect 57808 485790 57836 583986
rect 59084 583024 59136 583030
rect 59084 582966 59136 582972
rect 57888 581188 57940 581194
rect 57888 581130 57940 581136
rect 57900 537810 57928 581130
rect 58992 560380 59044 560386
rect 58992 560322 59044 560328
rect 58624 553444 58676 553450
rect 58624 553386 58676 553392
rect 57888 537804 57940 537810
rect 57888 537746 57940 537752
rect 57888 537668 57940 537674
rect 57888 537610 57940 537616
rect 57796 485784 57848 485790
rect 57796 485726 57848 485732
rect 57244 463684 57296 463690
rect 57244 463626 57296 463632
rect 56598 387832 56654 387841
rect 56598 387767 56654 387776
rect 57256 369170 57284 463626
rect 57702 453928 57758 453937
rect 57702 453863 57758 453872
rect 57716 453422 57744 453863
rect 57704 453416 57756 453422
rect 57704 453358 57756 453364
rect 57900 438161 57928 537610
rect 58636 492697 58664 553386
rect 58900 492788 58952 492794
rect 58900 492730 58952 492736
rect 58622 492688 58678 492697
rect 58622 492623 58678 492632
rect 58636 491298 58664 492623
rect 58624 491292 58676 491298
rect 58624 491234 58676 491240
rect 57886 438152 57942 438161
rect 57886 438087 57942 438096
rect 57612 394052 57664 394058
rect 57612 393994 57664 394000
rect 57624 393514 57652 393994
rect 57612 393508 57664 393514
rect 57612 393450 57664 393456
rect 57336 389904 57388 389910
rect 57336 389846 57388 389852
rect 57348 372570 57376 389846
rect 57336 372564 57388 372570
rect 57336 372506 57388 372512
rect 57244 369164 57296 369170
rect 57244 369106 57296 369112
rect 57256 364334 57284 369106
rect 57256 364306 57560 364334
rect 56508 358760 56560 358766
rect 56508 358702 56560 358708
rect 56416 337952 56468 337958
rect 56416 337894 56468 337900
rect 56508 334620 56560 334626
rect 56508 334562 56560 334568
rect 56322 300112 56378 300121
rect 56322 300047 56378 300056
rect 56416 279472 56468 279478
rect 56416 279414 56468 279420
rect 56428 278798 56456 279414
rect 56416 278792 56468 278798
rect 56416 278734 56468 278740
rect 56324 255400 56376 255406
rect 56324 255342 56376 255348
rect 55128 233232 55180 233238
rect 55128 233174 55180 233180
rect 56336 225690 56364 255342
rect 56324 225684 56376 225690
rect 56324 225626 56376 225632
rect 56428 207670 56456 278734
rect 56520 260846 56548 334562
rect 57532 304298 57560 364306
rect 57624 314022 57652 393450
rect 57900 338026 57928 438087
rect 58912 390114 58940 492730
rect 59004 462330 59032 560322
rect 59096 536790 59124 582966
rect 59188 558210 59216 586638
rect 60648 583908 60700 583914
rect 60648 583850 60700 583856
rect 59268 578332 59320 578338
rect 59268 578274 59320 578280
rect 59176 558204 59228 558210
rect 59176 558146 59228 558152
rect 59084 536784 59136 536790
rect 59084 536726 59136 536732
rect 59096 536178 59124 536726
rect 59084 536172 59136 536178
rect 59084 536114 59136 536120
rect 59280 512038 59308 578274
rect 60464 567248 60516 567254
rect 60464 567190 60516 567196
rect 60280 542496 60332 542502
rect 60280 542438 60332 542444
rect 59268 512032 59320 512038
rect 59268 511974 59320 511980
rect 59084 490816 59136 490822
rect 59084 490758 59136 490764
rect 58992 462324 59044 462330
rect 58992 462266 59044 462272
rect 59096 436082 59124 490758
rect 59280 480865 59308 511974
rect 59266 480856 59322 480865
rect 59266 480791 59322 480800
rect 59280 480282 59308 480791
rect 59268 480276 59320 480282
rect 59268 480218 59320 480224
rect 59176 465044 59228 465050
rect 59176 464986 59228 464992
rect 59084 436076 59136 436082
rect 59084 436018 59136 436024
rect 58990 407008 59046 407017
rect 58990 406943 59046 406952
rect 59004 405793 59032 406943
rect 58990 405784 59046 405793
rect 58990 405719 59046 405728
rect 58900 390108 58952 390114
rect 58900 390050 58952 390056
rect 58912 389842 58940 390050
rect 58900 389836 58952 389842
rect 58900 389778 58952 389784
rect 58530 388376 58586 388385
rect 58530 388311 58586 388320
rect 58544 387870 58572 388311
rect 58532 387864 58584 387870
rect 58532 387806 58584 387812
rect 59004 373998 59032 405719
rect 59084 387184 59136 387190
rect 59084 387126 59136 387132
rect 58992 373992 59044 373998
rect 58992 373934 59044 373940
rect 58992 367804 59044 367810
rect 58992 367746 59044 367752
rect 57888 338020 57940 338026
rect 57888 337962 57940 337968
rect 57900 335354 57928 337962
rect 57808 335326 57928 335354
rect 57704 333328 57756 333334
rect 57704 333270 57756 333276
rect 57612 314016 57664 314022
rect 57612 313958 57664 313964
rect 57520 304292 57572 304298
rect 57520 304234 57572 304240
rect 57612 270564 57664 270570
rect 57612 270506 57664 270512
rect 56508 260840 56560 260846
rect 56508 260782 56560 260788
rect 56508 249144 56560 249150
rect 56508 249086 56560 249092
rect 56416 207664 56468 207670
rect 56416 207606 56468 207612
rect 55036 205080 55088 205086
rect 55036 205022 55088 205028
rect 56520 195265 56548 249086
rect 57624 235278 57652 270506
rect 57716 238610 57744 333270
rect 57808 238678 57836 335326
rect 59004 335102 59032 367746
rect 59096 336734 59124 387126
rect 59188 367878 59216 464986
rect 60292 442814 60320 542438
rect 60372 474700 60424 474706
rect 60372 474642 60424 474648
rect 60280 442808 60332 442814
rect 60280 442750 60332 442756
rect 59268 395480 59320 395486
rect 59268 395422 59320 395428
rect 59176 367872 59228 367878
rect 59176 367814 59228 367820
rect 59176 355360 59228 355366
rect 59176 355302 59228 355308
rect 59188 354754 59216 355302
rect 59176 354748 59228 354754
rect 59176 354690 59228 354696
rect 59084 336728 59136 336734
rect 59084 336670 59136 336676
rect 58992 335096 59044 335102
rect 58992 335038 59044 335044
rect 59188 298790 59216 354690
rect 59280 331226 59308 395422
rect 60384 380798 60412 474642
rect 60476 469169 60504 567190
rect 60556 546508 60608 546514
rect 60556 546450 60608 546456
rect 60462 469160 60518 469169
rect 60462 469095 60518 469104
rect 60476 467945 60504 469095
rect 60462 467936 60518 467945
rect 60462 467871 60518 467880
rect 60568 460934 60596 546450
rect 60660 541686 60688 583850
rect 61936 572756 61988 572762
rect 61936 572698 61988 572704
rect 60740 562352 60792 562358
rect 60740 562294 60792 562300
rect 60752 560998 60780 562294
rect 61752 561740 61804 561746
rect 61752 561682 61804 561688
rect 60740 560992 60792 560998
rect 60740 560934 60792 560940
rect 60648 541680 60700 541686
rect 60648 541622 60700 541628
rect 61764 462398 61792 561682
rect 61844 549296 61896 549302
rect 61844 549238 61896 549244
rect 61752 462392 61804 462398
rect 61752 462334 61804 462340
rect 60568 460906 60688 460934
rect 60660 445754 60688 460906
rect 61856 449954 61884 549238
rect 61948 474706 61976 572698
rect 62040 562358 62068 700266
rect 68744 596828 68796 596834
rect 68744 596770 68796 596776
rect 68756 596174 68784 596770
rect 68572 596146 68784 596174
rect 68468 583976 68520 583982
rect 68468 583918 68520 583924
rect 66168 581868 66220 581874
rect 66168 581810 66220 581816
rect 66076 577448 66128 577454
rect 66076 577390 66128 577396
rect 65984 572824 66036 572830
rect 65984 572766 66036 572772
rect 63224 569968 63276 569974
rect 63224 569910 63276 569916
rect 63132 563168 63184 563174
rect 63132 563110 63184 563116
rect 62028 562352 62080 562358
rect 62028 562294 62080 562300
rect 62028 539640 62080 539646
rect 62028 539582 62080 539588
rect 61936 474700 61988 474706
rect 61936 474642 61988 474648
rect 61936 471980 61988 471986
rect 61936 471922 61988 471928
rect 61844 449948 61896 449954
rect 61844 449890 61896 449896
rect 61384 447160 61436 447166
rect 61384 447102 61436 447108
rect 60740 445800 60792 445806
rect 60660 445748 60740 445754
rect 60660 445742 60792 445748
rect 60660 445726 60780 445742
rect 60648 387116 60700 387122
rect 60648 387058 60700 387064
rect 60372 380792 60424 380798
rect 60372 380734 60424 380740
rect 60188 380248 60240 380254
rect 60188 380190 60240 380196
rect 60200 379574 60228 380190
rect 60188 379568 60240 379574
rect 60188 379510 60240 379516
rect 60464 379568 60516 379574
rect 60464 379510 60516 379516
rect 60188 367056 60240 367062
rect 60188 366998 60240 367004
rect 60200 366382 60228 366998
rect 60188 366376 60240 366382
rect 60188 366318 60240 366324
rect 60200 365945 60228 366318
rect 60186 365936 60242 365945
rect 60186 365871 60242 365880
rect 59360 358760 59412 358766
rect 59360 358702 59412 358708
rect 59372 357474 59400 358702
rect 59360 357468 59412 357474
rect 59360 357410 59412 357416
rect 59268 331220 59320 331226
rect 59268 331162 59320 331168
rect 59176 298784 59228 298790
rect 59176 298726 59228 298732
rect 57888 296880 57940 296886
rect 57888 296822 57940 296828
rect 57796 238672 57848 238678
rect 57796 238614 57848 238620
rect 57704 238604 57756 238610
rect 57704 238546 57756 238552
rect 57612 235272 57664 235278
rect 57612 235214 57664 235220
rect 56506 195256 56562 195265
rect 56506 195191 56562 195200
rect 54944 188352 54996 188358
rect 54944 188294 54996 188300
rect 53748 181484 53800 181490
rect 53748 181426 53800 181432
rect 57900 71738 57928 296822
rect 59176 280288 59228 280294
rect 59176 280230 59228 280236
rect 59084 249076 59136 249082
rect 59084 249018 59136 249024
rect 59096 248470 59124 249018
rect 59084 248464 59136 248470
rect 59084 248406 59136 248412
rect 58624 242888 58676 242894
rect 58624 242830 58676 242836
rect 58636 211818 58664 242830
rect 59096 222902 59124 248406
rect 59188 224330 59216 280230
rect 59372 272082 59400 357410
rect 60476 330546 60504 379510
rect 60556 365764 60608 365770
rect 60556 365706 60608 365712
rect 60568 364342 60596 365706
rect 60556 364336 60608 364342
rect 60556 364278 60608 364284
rect 60556 337408 60608 337414
rect 60556 337350 60608 337356
rect 60464 330540 60516 330546
rect 60464 330482 60516 330488
rect 59280 272054 59400 272082
rect 59280 271182 59308 272054
rect 59268 271176 59320 271182
rect 59268 271118 59320 271124
rect 59176 224324 59228 224330
rect 59176 224266 59228 224272
rect 59084 222896 59136 222902
rect 59084 222838 59136 222844
rect 58624 211812 58676 211818
rect 58624 211754 58676 211760
rect 59280 195294 59308 271118
rect 60188 267028 60240 267034
rect 60188 266970 60240 266976
rect 60200 266422 60228 266970
rect 60188 266416 60240 266422
rect 60188 266358 60240 266364
rect 60464 266416 60516 266422
rect 60464 266358 60516 266364
rect 60004 254584 60056 254590
rect 60004 254526 60056 254532
rect 60016 238814 60044 254526
rect 60004 238808 60056 238814
rect 60004 238750 60056 238756
rect 59268 195288 59320 195294
rect 59268 195230 59320 195236
rect 60476 192506 60504 266358
rect 60568 254590 60596 337350
rect 60660 335170 60688 387058
rect 61396 349178 61424 447102
rect 61752 445800 61804 445806
rect 61750 445768 61752 445777
rect 61804 445768 61806 445777
rect 61750 445703 61806 445712
rect 61844 442808 61896 442814
rect 61844 442750 61896 442756
rect 61476 356040 61528 356046
rect 61476 355982 61528 355988
rect 61384 349172 61436 349178
rect 61384 349114 61436 349120
rect 60648 335164 60700 335170
rect 60648 335106 60700 335112
rect 60660 334121 60688 335106
rect 60646 334112 60702 334121
rect 60646 334047 60702 334056
rect 61488 301481 61516 355982
rect 61856 342310 61884 442750
rect 61948 397526 61976 471922
rect 62040 441590 62068 539582
rect 63144 465050 63172 563110
rect 63236 471986 63264 569910
rect 64604 567316 64656 567322
rect 64604 567258 64656 567264
rect 63316 549364 63368 549370
rect 63316 549306 63368 549312
rect 63224 471980 63276 471986
rect 63224 471922 63276 471928
rect 63132 465044 63184 465050
rect 63132 464986 63184 464992
rect 63132 462324 63184 462330
rect 63132 462266 63184 462272
rect 63144 460970 63172 462266
rect 63132 460964 63184 460970
rect 63132 460906 63184 460912
rect 62028 441584 62080 441590
rect 62028 441526 62080 441532
rect 61936 397520 61988 397526
rect 61936 397462 61988 397468
rect 61948 376650 61976 397462
rect 61936 376644 61988 376650
rect 61936 376586 61988 376592
rect 63144 365022 63172 460906
rect 63328 448594 63356 549306
rect 64144 541068 64196 541074
rect 64144 541010 64196 541016
rect 63408 541000 63460 541006
rect 63408 540942 63460 540948
rect 63316 448588 63368 448594
rect 63316 448530 63368 448536
rect 63222 447400 63278 447409
rect 63222 447335 63278 447344
rect 63132 365016 63184 365022
rect 63132 364958 63184 364964
rect 63236 348498 63264 447335
rect 63420 441590 63448 540942
rect 64156 525842 64184 541010
rect 64144 525836 64196 525842
rect 64144 525778 64196 525784
rect 63498 491328 63554 491337
rect 63498 491263 63500 491272
rect 63552 491263 63554 491272
rect 63500 491234 63552 491240
rect 64512 484560 64564 484566
rect 64512 484502 64564 484508
rect 64420 449948 64472 449954
rect 64420 449890 64472 449896
rect 64432 442338 64460 449890
rect 64420 442332 64472 442338
rect 64420 442274 64472 442280
rect 63316 441584 63368 441590
rect 63316 441526 63368 441532
rect 63408 441584 63460 441590
rect 63408 441526 63460 441532
rect 63328 441046 63356 441526
rect 63316 441040 63368 441046
rect 63316 440982 63368 440988
rect 63224 348492 63276 348498
rect 63224 348434 63276 348440
rect 61936 345704 61988 345710
rect 61936 345646 61988 345652
rect 61948 345166 61976 345646
rect 61936 345160 61988 345166
rect 61936 345102 61988 345108
rect 61844 342304 61896 342310
rect 61844 342246 61896 342252
rect 61948 331974 61976 345102
rect 62120 343664 62172 343670
rect 62120 343606 62172 343612
rect 62132 342922 62160 343606
rect 62120 342916 62172 342922
rect 62120 342858 62172 342864
rect 61936 331968 61988 331974
rect 61936 331910 61988 331916
rect 63236 325106 63264 348434
rect 63328 340882 63356 440982
rect 64418 437608 64474 437617
rect 64418 437543 64474 437552
rect 64432 432041 64460 437543
rect 64524 436762 64552 484502
rect 64616 467906 64644 567258
rect 64696 565888 64748 565894
rect 64696 565830 64748 565836
rect 64604 467900 64656 467906
rect 64604 467842 64656 467848
rect 64708 466478 64736 565830
rect 64788 558272 64840 558278
rect 64788 558214 64840 558220
rect 64696 466472 64748 466478
rect 64696 466414 64748 466420
rect 64604 462392 64656 462398
rect 64604 462334 64656 462340
rect 64512 436756 64564 436762
rect 64512 436698 64564 436704
rect 64418 432032 64474 432041
rect 64418 431967 64474 431976
rect 64510 431896 64566 431905
rect 64510 431831 64566 431840
rect 64524 422385 64552 431831
rect 64510 422376 64566 422385
rect 64510 422311 64566 422320
rect 64510 412584 64566 412593
rect 64510 412519 64566 412528
rect 64524 403073 64552 412519
rect 64510 403064 64566 403073
rect 64510 402999 64566 403008
rect 64510 400344 64566 400353
rect 64510 400279 64566 400288
rect 63408 374672 63460 374678
rect 63408 374614 63460 374620
rect 63316 340876 63368 340882
rect 63316 340818 63368 340824
rect 63224 325100 63276 325106
rect 63224 325042 63276 325048
rect 61474 301472 61530 301481
rect 61474 301407 61530 301416
rect 60648 276140 60700 276146
rect 60648 276082 60700 276088
rect 60556 254584 60608 254590
rect 60556 254526 60608 254532
rect 60568 225758 60596 254526
rect 60556 225752 60608 225758
rect 60556 225694 60608 225700
rect 60660 194002 60688 276082
rect 60740 266552 60792 266558
rect 60740 266494 60792 266500
rect 61384 266552 61436 266558
rect 61384 266494 61436 266500
rect 60752 266354 60780 266494
rect 60740 266348 60792 266354
rect 60740 266290 60792 266296
rect 61396 218754 61424 266494
rect 62026 265704 62082 265713
rect 62026 265639 62028 265648
rect 62080 265639 62082 265648
rect 62028 265610 62080 265616
rect 63132 259480 63184 259486
rect 63132 259422 63184 259428
rect 61844 256828 61896 256834
rect 61844 256770 61896 256776
rect 61384 218748 61436 218754
rect 61384 218690 61436 218696
rect 61856 198014 61884 256770
rect 61936 247104 61988 247110
rect 61936 247046 61988 247052
rect 61948 235414 61976 247046
rect 61936 235408 61988 235414
rect 61936 235350 61988 235356
rect 63144 203658 63172 259422
rect 63316 258188 63368 258194
rect 63316 258130 63368 258136
rect 63224 247172 63276 247178
rect 63224 247114 63276 247120
rect 63132 203652 63184 203658
rect 63132 203594 63184 203600
rect 61844 198008 61896 198014
rect 61844 197950 61896 197956
rect 60648 193996 60700 194002
rect 60648 193938 60700 193944
rect 60464 192500 60516 192506
rect 60464 192442 60516 192448
rect 63236 184346 63264 247114
rect 63224 184340 63276 184346
rect 63224 184282 63276 184288
rect 63328 180033 63356 258130
rect 63314 180024 63370 180033
rect 63314 179959 63370 179968
rect 59268 125656 59320 125662
rect 59268 125598 59320 125604
rect 59280 75886 59308 125598
rect 59268 75880 59320 75886
rect 59268 75822 59320 75828
rect 57888 71732 57940 71738
rect 57888 71674 57940 71680
rect 60740 71052 60792 71058
rect 60740 70994 60792 71000
rect 51172 64184 51224 64190
rect 51172 64126 51224 64132
rect 51080 59356 51132 59362
rect 51080 59298 51132 59304
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 45100 3528 45152 3534
rect 45100 3470 45152 3476
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45112 354 45140 3470
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51184 354 51212 64126
rect 57980 62824 58032 62830
rect 57980 62766 58032 62772
rect 52460 55956 52512 55962
rect 52460 55898 52512 55904
rect 52472 3534 52500 55898
rect 56600 49020 56652 49026
rect 56600 48962 56652 48968
rect 52552 43512 52604 43518
rect 52552 43454 52604 43460
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 52564 480 52592 43454
rect 53840 42084 53892 42090
rect 53840 42026 53892 42032
rect 53852 16574 53880 42026
rect 55220 32428 55272 32434
rect 55220 32370 55272 32376
rect 55232 16574 55260 32370
rect 56612 16574 56640 48962
rect 57992 16574 58020 62766
rect 59360 29640 59412 29646
rect 59360 29582 59412 29588
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 53380 3528 53432 3534
rect 53380 3470 53432 3476
rect 51326 354 51438 480
rect 51184 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53392 354 53420 3470
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 29582
rect 60752 6914 60780 70994
rect 60832 54596 60884 54602
rect 60832 54538 60884 54544
rect 60844 16574 60872 54538
rect 60844 16546 61608 16574
rect 60752 6886 60872 6914
rect 60844 480 60872 6886
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63420 11762 63448 374614
rect 64524 370666 64552 400279
rect 64512 370660 64564 370666
rect 64512 370602 64564 370608
rect 64616 366450 64644 462334
rect 64694 460864 64750 460873
rect 64694 460799 64750 460808
rect 64708 451489 64736 460799
rect 64800 458250 64828 558214
rect 65892 536240 65944 536246
rect 65892 536182 65944 536188
rect 65904 535430 65932 536182
rect 65892 535424 65944 535430
rect 65892 535366 65944 535372
rect 65524 485852 65576 485858
rect 65524 485794 65576 485800
rect 64788 458244 64840 458250
rect 64788 458186 64840 458192
rect 64694 451480 64750 451489
rect 64694 451415 64750 451424
rect 64786 451208 64842 451217
rect 64786 451143 64842 451152
rect 64696 448588 64748 448594
rect 64696 448530 64748 448536
rect 64604 366444 64656 366450
rect 64604 366386 64656 366392
rect 64708 351218 64736 448530
rect 64800 447137 64828 451143
rect 64786 447128 64842 447137
rect 64786 447063 64842 447072
rect 64788 442332 64840 442338
rect 64788 442274 64840 442280
rect 64800 352646 64828 442274
rect 65536 435402 65564 485794
rect 65996 475386 66024 572766
rect 66088 479738 66116 577390
rect 66180 571334 66208 581810
rect 67638 581360 67694 581369
rect 67638 581295 67694 581304
rect 67652 581262 67680 581295
rect 67640 581256 67692 581262
rect 67640 581198 67692 581204
rect 67822 580680 67878 580689
rect 67822 580615 67878 580624
rect 67836 580310 67864 580615
rect 67824 580304 67876 580310
rect 67824 580246 67876 580252
rect 67362 579184 67418 579193
rect 67362 579119 67418 579128
rect 66168 571328 66220 571334
rect 66168 571270 66220 571276
rect 66168 568676 66220 568682
rect 66168 568618 66220 568624
rect 66076 479732 66128 479738
rect 66076 479674 66128 479680
rect 65984 475380 66036 475386
rect 65984 475322 66036 475328
rect 65616 473408 65668 473414
rect 65616 473350 65668 473356
rect 65628 466177 65656 473350
rect 65984 467900 66036 467906
rect 65984 467842 66036 467848
rect 65614 466168 65670 466177
rect 65614 466103 65670 466112
rect 65524 435396 65576 435402
rect 65524 435338 65576 435344
rect 65996 398886 66024 467842
rect 65984 398880 66036 398886
rect 65984 398822 66036 398828
rect 65154 379536 65210 379545
rect 65154 379471 65210 379480
rect 65168 378826 65196 379471
rect 65156 378820 65208 378826
rect 65156 378762 65208 378768
rect 65524 376780 65576 376786
rect 65524 376722 65576 376728
rect 64788 352640 64840 352646
rect 64788 352582 64840 352588
rect 64696 351212 64748 351218
rect 64696 351154 64748 351160
rect 64420 349172 64472 349178
rect 64420 349114 64472 349120
rect 63500 348424 63552 348430
rect 63500 348366 63552 348372
rect 63512 347750 63540 348366
rect 63500 347744 63552 347750
rect 63500 347686 63552 347692
rect 64144 340944 64196 340950
rect 64144 340886 64196 340892
rect 64156 331906 64184 340886
rect 64144 331900 64196 331906
rect 64144 331842 64196 331848
rect 64432 72486 64460 349114
rect 64800 338774 64828 352582
rect 64788 338768 64840 338774
rect 64788 338710 64840 338716
rect 65536 311914 65564 376722
rect 65996 373182 66024 398822
rect 66088 386306 66116 479674
rect 66180 469946 66208 568618
rect 67270 564496 67326 564505
rect 67270 564431 67326 564440
rect 66902 477456 66958 477465
rect 66902 477391 66958 477400
rect 66916 476513 66944 477391
rect 66902 476504 66958 476513
rect 66902 476439 66958 476448
rect 66168 469940 66220 469946
rect 66168 469882 66220 469888
rect 66258 443048 66314 443057
rect 66258 442983 66314 442992
rect 66272 442882 66300 442983
rect 66260 442876 66312 442882
rect 66260 442818 66312 442824
rect 66168 441584 66220 441590
rect 66168 441526 66220 441532
rect 66180 441182 66208 441526
rect 66168 441176 66220 441182
rect 66168 441118 66220 441124
rect 66076 386300 66128 386306
rect 66076 386242 66128 386248
rect 65984 373176 66036 373182
rect 65984 373118 66036 373124
rect 65984 358080 66036 358086
rect 65984 358022 66036 358028
rect 65524 311908 65576 311914
rect 65524 311850 65576 311856
rect 65996 296041 66024 358022
rect 66076 342304 66128 342310
rect 66076 342246 66128 342252
rect 66088 327826 66116 342246
rect 66180 341630 66208 441118
rect 66916 382129 66944 476439
rect 66996 469192 67048 469198
rect 66996 469134 67048 469140
rect 66902 382120 66958 382129
rect 66902 382055 66958 382064
rect 67008 375902 67036 469134
rect 67284 466449 67312 564431
rect 67376 480593 67404 579119
rect 67638 578504 67694 578513
rect 67638 578439 67694 578448
rect 67652 578338 67680 578439
rect 67640 578332 67692 578338
rect 67640 578274 67692 578280
rect 68190 577824 68246 577833
rect 68190 577759 68246 577768
rect 68204 577454 68232 577759
rect 68192 577448 68244 577454
rect 68192 577390 68244 577396
rect 67546 577144 67602 577153
rect 67546 577079 67602 577088
rect 67456 512032 67508 512038
rect 67456 511974 67508 511980
rect 67468 511290 67496 511974
rect 67456 511284 67508 511290
rect 67456 511226 67508 511232
rect 67560 485774 67588 577079
rect 67638 575784 67694 575793
rect 67638 575719 67694 575728
rect 67652 575550 67680 575719
rect 67640 575544 67692 575550
rect 67640 575486 67692 575492
rect 67638 574424 67694 574433
rect 67638 574359 67694 574368
rect 67652 574122 67680 574359
rect 67640 574116 67692 574122
rect 67640 574058 67692 574064
rect 67730 573472 67786 573481
rect 67730 573407 67786 573416
rect 67638 573064 67694 573073
rect 67638 572999 67694 573008
rect 67652 572762 67680 572999
rect 67744 572830 67772 573407
rect 67732 572824 67784 572830
rect 67732 572766 67784 572772
rect 67640 572756 67692 572762
rect 67640 572698 67692 572704
rect 67824 572076 67876 572082
rect 67824 572018 67876 572024
rect 67836 571713 67864 572018
rect 67916 572008 67968 572014
rect 67916 571950 67968 571956
rect 67928 571849 67956 571950
rect 67914 571840 67970 571849
rect 67914 571775 67970 571784
rect 68480 571713 68508 583918
rect 68572 580689 68600 596146
rect 68940 586514 68968 702442
rect 69664 700392 69716 700398
rect 69664 700334 69716 700340
rect 69020 594108 69072 594114
rect 69020 594050 69072 594056
rect 68664 586486 68968 586514
rect 68558 580680 68614 580689
rect 68558 580615 68614 580624
rect 68664 571849 68692 586486
rect 68836 585812 68888 585818
rect 68836 585754 68888 585760
rect 68744 581732 68796 581738
rect 68744 581674 68796 581680
rect 68756 581126 68784 581674
rect 68744 581120 68796 581126
rect 68744 581062 68796 581068
rect 68742 576464 68798 576473
rect 68742 576399 68798 576408
rect 68650 571840 68706 571849
rect 68650 571775 68706 571784
rect 67822 571704 67878 571713
rect 67822 571639 67878 571648
rect 68466 571704 68522 571713
rect 68466 571639 68522 571648
rect 68284 571328 68336 571334
rect 68284 571270 68336 571276
rect 67638 570072 67694 570081
rect 67638 570007 67694 570016
rect 67652 569974 67680 570007
rect 67640 569968 67692 569974
rect 67640 569910 67692 569916
rect 67638 568984 67694 568993
rect 67638 568919 67694 568928
rect 67652 568614 67680 568919
rect 67730 568712 67786 568721
rect 67730 568647 67732 568656
rect 67784 568647 67786 568656
rect 67732 568618 67784 568624
rect 67640 568608 67692 568614
rect 67640 568550 67692 568556
rect 67730 567624 67786 567633
rect 67730 567559 67786 567568
rect 67640 567316 67692 567322
rect 67640 567258 67692 567264
rect 67652 567225 67680 567258
rect 67744 567254 67772 567559
rect 67732 567248 67784 567254
rect 67638 567216 67694 567225
rect 67732 567190 67784 567196
rect 67638 567151 67694 567160
rect 67640 565888 67692 565894
rect 67638 565856 67640 565865
rect 67692 565856 67694 565865
rect 67638 565791 67694 565800
rect 67638 564904 67694 564913
rect 67638 564839 67694 564848
rect 67652 564534 67680 564839
rect 67640 564528 67692 564534
rect 67640 564470 67692 564476
rect 67730 563544 67786 563553
rect 67730 563479 67786 563488
rect 67640 563168 67692 563174
rect 67638 563136 67640 563145
rect 67692 563136 67694 563145
rect 67744 563106 67772 563479
rect 67638 563071 67694 563080
rect 67732 563100 67784 563106
rect 67732 563042 67784 563048
rect 67640 562352 67692 562358
rect 67638 562320 67640 562329
rect 67692 562320 67694 562329
rect 67638 562255 67694 562264
rect 67638 562184 67694 562193
rect 67638 562119 67694 562128
rect 67652 561746 67680 562119
rect 67640 561740 67692 561746
rect 67640 561682 67692 561688
rect 67730 560824 67786 560833
rect 67730 560759 67786 560768
rect 67638 560416 67694 560425
rect 67744 560386 67772 560759
rect 67638 560351 67694 560360
rect 67732 560380 67784 560386
rect 67652 560318 67680 560351
rect 67732 560322 67784 560328
rect 67640 560312 67692 560318
rect 67640 560254 67692 560260
rect 67638 559464 67694 559473
rect 67638 559399 67694 559408
rect 67652 558958 67680 559399
rect 67640 558952 67692 558958
rect 67640 558894 67692 558900
rect 68296 557433 68324 571270
rect 68282 557424 68338 557433
rect 68282 557359 68338 557368
rect 67730 556744 67786 556753
rect 67730 556679 67786 556688
rect 67640 556300 67692 556306
rect 67640 556242 67692 556248
rect 67652 556209 67680 556242
rect 67744 556238 67772 556679
rect 67732 556232 67784 556238
rect 67638 556200 67694 556209
rect 67732 556174 67784 556180
rect 67638 556135 67694 556144
rect 67730 555384 67786 555393
rect 67730 555319 67786 555328
rect 67640 554872 67692 554878
rect 67638 554840 67640 554849
rect 67692 554840 67694 554849
rect 67744 554810 67772 555319
rect 67638 554775 67694 554784
rect 67732 554804 67784 554810
rect 67732 554746 67784 554752
rect 67638 553480 67694 553489
rect 67638 553415 67640 553424
rect 67692 553415 67694 553424
rect 67640 553386 67692 553392
rect 67638 552120 67694 552129
rect 67638 552055 67640 552064
rect 67692 552055 67694 552064
rect 67640 552026 67692 552032
rect 67638 551304 67694 551313
rect 67638 551239 67694 551248
rect 67652 550662 67680 551239
rect 67640 550656 67692 550662
rect 67640 550598 67692 550604
rect 67730 549944 67786 549953
rect 67730 549879 67786 549888
rect 67638 549400 67694 549409
rect 67638 549335 67640 549344
rect 67692 549335 67694 549344
rect 67640 549306 67692 549312
rect 67744 549302 67772 549879
rect 67732 549296 67784 549302
rect 67732 549238 67784 549244
rect 67638 548040 67694 548049
rect 67638 547975 67694 547984
rect 67652 547942 67680 547975
rect 67640 547936 67692 547942
rect 67640 547878 67692 547884
rect 67638 546544 67694 546553
rect 67638 546479 67640 546488
rect 67692 546479 67694 546488
rect 67640 546450 67692 546456
rect 67732 544400 67784 544406
rect 67732 544342 67784 544348
rect 67744 543969 67772 544342
rect 67730 543960 67786 543969
rect 67730 543895 67786 543904
rect 68282 543960 68338 543969
rect 68282 543895 68338 543904
rect 68006 543280 68062 543289
rect 68006 543215 68062 543224
rect 67638 542600 67694 542609
rect 67638 542535 67694 542544
rect 67652 542502 67680 542535
rect 67640 542496 67692 542502
rect 67640 542438 67692 542444
rect 68020 542434 68048 543215
rect 68008 542428 68060 542434
rect 68008 542370 68060 542376
rect 67730 541784 67786 541793
rect 67730 541719 67786 541728
rect 67638 541240 67694 541249
rect 67638 541175 67694 541184
rect 67652 541006 67680 541175
rect 67744 541074 67772 541719
rect 67732 541068 67784 541074
rect 67732 541010 67784 541016
rect 67640 541000 67692 541006
rect 67640 540942 67692 540948
rect 67638 540152 67694 540161
rect 67638 540087 67694 540096
rect 67652 539646 67680 540087
rect 67640 539640 67692 539646
rect 67640 539582 67692 539588
rect 67638 487928 67694 487937
rect 67638 487863 67694 487872
rect 67652 487830 67680 487863
rect 67640 487824 67692 487830
rect 67640 487766 67692 487772
rect 67638 487248 67694 487257
rect 67638 487183 67640 487192
rect 67692 487183 67694 487192
rect 67640 487154 67692 487160
rect 68100 487144 68152 487150
rect 68100 487086 68152 487092
rect 67638 486568 67694 486577
rect 67638 486503 67694 486512
rect 67652 485858 67680 486503
rect 68112 486033 68140 487086
rect 68098 486024 68154 486033
rect 68098 485959 68154 485968
rect 67640 485852 67692 485858
rect 67640 485794 67692 485800
rect 67468 485746 67588 485774
rect 67362 480584 67418 480593
rect 67362 480519 67418 480528
rect 67468 478553 67496 485746
rect 67638 485208 67694 485217
rect 67638 485143 67694 485152
rect 67652 484430 67680 485143
rect 67640 484424 67692 484430
rect 67640 484366 67692 484372
rect 67640 482996 67692 483002
rect 67640 482938 67692 482944
rect 67652 482633 67680 482938
rect 67638 482624 67694 482633
rect 67638 482559 67694 482568
rect 67638 481128 67694 481137
rect 67638 481063 67694 481072
rect 67652 480962 67680 481063
rect 67640 480956 67692 480962
rect 67640 480898 67692 480904
rect 67548 480276 67600 480282
rect 67548 480218 67600 480224
rect 67560 479913 67588 480218
rect 67546 479904 67602 479913
rect 67546 479839 67602 479848
rect 67454 478544 67510 478553
rect 67454 478479 67510 478488
rect 67638 477048 67694 477057
rect 67638 476983 67694 476992
rect 67652 476134 67680 476983
rect 67640 476128 67692 476134
rect 67640 476070 67692 476076
rect 67638 475688 67694 475697
rect 67638 475623 67694 475632
rect 67652 475454 67680 475623
rect 67640 475448 67692 475454
rect 67640 475390 67692 475396
rect 67732 475380 67784 475386
rect 67732 475322 67784 475328
rect 67744 475153 67772 475322
rect 67730 475144 67786 475153
rect 67730 475079 67786 475088
rect 67640 474700 67692 474706
rect 67640 474642 67692 474648
rect 67652 474337 67680 474642
rect 67638 474328 67694 474337
rect 67638 474263 67694 474272
rect 67638 473648 67694 473657
rect 67638 473583 67694 473592
rect 67652 473414 67680 473583
rect 67640 473408 67692 473414
rect 67640 473350 67692 473356
rect 67640 472660 67692 472666
rect 67640 472602 67692 472608
rect 67652 472569 67680 472602
rect 67638 472560 67694 472569
rect 67638 472495 67694 472504
rect 67640 471980 67692 471986
rect 67640 471922 67692 471928
rect 67652 471073 67680 471922
rect 67638 471064 67694 471073
rect 67638 470999 67694 471008
rect 67546 470248 67602 470257
rect 67546 470183 67602 470192
rect 67560 469198 67588 470183
rect 67640 469940 67692 469946
rect 67640 469882 67692 469888
rect 67652 469713 67680 469882
rect 67638 469704 67694 469713
rect 67638 469639 67694 469648
rect 67548 469192 67600 469198
rect 67548 469134 67600 469140
rect 67638 468208 67694 468217
rect 67638 468143 67694 468152
rect 67652 467906 67680 468143
rect 67640 467900 67692 467906
rect 67640 467842 67692 467848
rect 67638 466848 67694 466857
rect 67638 466783 67694 466792
rect 67652 466478 67680 466783
rect 67640 466472 67692 466478
rect 67270 466440 67326 466449
rect 67270 466375 67326 466384
rect 67454 466440 67510 466449
rect 67454 466375 67510 466384
rect 67560 466432 67640 466460
rect 67468 465633 67496 466375
rect 67454 465624 67510 465633
rect 67454 465559 67510 465568
rect 67560 460934 67588 466432
rect 67640 466414 67692 466420
rect 67638 466168 67694 466177
rect 67638 466103 67694 466112
rect 67652 465118 67680 466103
rect 67640 465112 67692 465118
rect 67640 465054 67692 465060
rect 67732 465044 67784 465050
rect 67732 464986 67784 464992
rect 67638 464808 67694 464817
rect 67638 464743 67694 464752
rect 67652 463758 67680 464743
rect 67744 464273 67772 464986
rect 67730 464264 67786 464273
rect 67730 464199 67786 464208
rect 67640 463752 67692 463758
rect 67640 463694 67692 463700
rect 67640 463004 67692 463010
rect 67640 462946 67692 462952
rect 67652 462913 67680 462946
rect 67638 462904 67694 462913
rect 67638 462839 67694 462848
rect 67638 462768 67694 462777
rect 67638 462703 67694 462712
rect 67652 462398 67680 462703
rect 67640 462392 67692 462398
rect 67640 462334 67692 462340
rect 67638 461408 67694 461417
rect 67638 461343 67694 461352
rect 67652 460970 67680 461343
rect 67468 460906 67588 460934
rect 67640 460964 67692 460970
rect 67640 460906 67692 460912
rect 67468 392018 67496 460906
rect 67638 460728 67694 460737
rect 67638 460663 67694 460672
rect 67652 460290 67680 460663
rect 67640 460284 67692 460290
rect 67640 460226 67692 460232
rect 67732 460216 67784 460222
rect 67730 460184 67732 460193
rect 67784 460184 67786 460193
rect 67730 460119 67786 460128
rect 67638 459368 67694 459377
rect 67638 459303 67694 459312
rect 67652 458250 67680 459303
rect 67640 458244 67692 458250
rect 67560 458204 67640 458232
rect 67456 392012 67508 392018
rect 67456 391954 67508 391960
rect 66996 375896 67048 375902
rect 66996 375838 67048 375844
rect 67468 371793 67496 391954
rect 67454 371784 67510 371793
rect 67454 371719 67510 371728
rect 67272 370592 67324 370598
rect 67272 370534 67324 370540
rect 67086 345944 67142 345953
rect 67086 345879 67142 345888
rect 67100 345098 67128 345879
rect 67088 345092 67140 345098
rect 67088 345034 67140 345040
rect 66168 341624 66220 341630
rect 66168 341566 66220 341572
rect 66076 327820 66128 327826
rect 66076 327762 66128 327768
rect 67284 312633 67312 370534
rect 67560 362386 67588 458204
rect 67640 458186 67692 458192
rect 67730 457328 67786 457337
rect 67730 457263 67786 457272
rect 67638 456920 67694 456929
rect 67638 456855 67640 456864
rect 67692 456855 67694 456864
rect 67640 456826 67692 456832
rect 67744 456822 67772 457263
rect 67732 456816 67784 456822
rect 67732 456758 67784 456764
rect 67638 455968 67694 455977
rect 67638 455903 67694 455912
rect 67652 455462 67680 455903
rect 67640 455456 67692 455462
rect 67640 455398 67692 455404
rect 67638 454744 67694 454753
rect 67638 454679 67640 454688
rect 67692 454679 67694 454688
rect 67640 454650 67692 454656
rect 67640 453416 67692 453422
rect 67638 453384 67640 453393
rect 67692 453384 67694 453393
rect 67638 453319 67694 453328
rect 67732 453348 67784 453354
rect 67732 453290 67784 453296
rect 67744 453257 67772 453290
rect 67730 453248 67786 453257
rect 67730 453183 67786 453192
rect 67638 449984 67694 449993
rect 67638 449919 67640 449928
rect 67692 449919 67694 449928
rect 67640 449890 67692 449896
rect 67638 449168 67694 449177
rect 67638 449103 67694 449112
rect 67652 448594 67680 449103
rect 67640 448588 67692 448594
rect 67640 448530 67692 448536
rect 67638 447808 67694 447817
rect 67638 447743 67694 447752
rect 67652 447166 67680 447743
rect 67640 447160 67692 447166
rect 67640 447102 67692 447108
rect 67638 446584 67694 446593
rect 67638 446519 67694 446528
rect 67652 445806 67680 446519
rect 67640 445800 67692 445806
rect 67640 445742 67692 445748
rect 67638 445088 67694 445097
rect 67638 445023 67640 445032
rect 67692 445023 67694 445032
rect 67640 444994 67692 445000
rect 68296 443873 68324 543895
rect 68756 489914 68784 576399
rect 68848 558929 68876 585754
rect 68834 558920 68890 558929
rect 68834 558855 68890 558864
rect 68848 558278 68876 558855
rect 68836 558272 68888 558278
rect 68836 558214 68888 558220
rect 68926 550760 68982 550769
rect 68926 550695 68982 550704
rect 68834 544504 68890 544513
rect 68834 544439 68890 544448
rect 68664 489886 68784 489914
rect 68374 484664 68430 484673
rect 68374 484599 68430 484608
rect 68388 484566 68416 484599
rect 68376 484560 68428 484566
rect 68376 484502 68428 484508
rect 68374 479768 68430 479777
rect 68374 479703 68376 479712
rect 68428 479703 68430 479712
rect 68376 479674 68428 479680
rect 68664 477193 68692 489886
rect 68650 477184 68706 477193
rect 68650 477119 68706 477128
rect 68664 476114 68692 477119
rect 68388 476086 68692 476114
rect 67638 443864 67694 443873
rect 67638 443799 67694 443808
rect 68282 443864 68338 443873
rect 68282 443799 68338 443808
rect 67652 443698 67680 443799
rect 67640 443692 67692 443698
rect 67640 443634 67692 443640
rect 67640 442944 67692 442950
rect 67640 442886 67692 442892
rect 67652 441833 67680 442886
rect 67732 442808 67784 442814
rect 67730 442776 67732 442785
rect 67784 442776 67786 442785
rect 67730 442711 67786 442720
rect 67638 441824 67694 441833
rect 67638 441759 67694 441768
rect 67640 441176 67692 441182
rect 67638 441144 67640 441153
rect 67692 441144 67694 441153
rect 67638 441079 67694 441088
rect 67640 441040 67692 441046
rect 67638 441008 67640 441017
rect 67692 441008 67694 441017
rect 67638 440943 67694 440952
rect 68388 402974 68416 476086
rect 68848 451274 68876 544439
rect 68940 451897 68968 550695
rect 69032 543289 69060 594050
rect 69676 583982 69704 700334
rect 70400 584044 70452 584050
rect 70400 583986 70452 583992
rect 69664 583976 69716 583982
rect 69664 583918 69716 583924
rect 69204 582412 69256 582418
rect 69204 582354 69256 582360
rect 69112 579080 69164 579086
rect 69112 579022 69164 579028
rect 69018 543280 69074 543289
rect 69018 543215 69074 543224
rect 69124 482905 69152 579022
rect 69216 545193 69244 582354
rect 70412 581890 70440 583986
rect 71792 583030 71820 702986
rect 75184 702840 75236 702846
rect 75184 702782 75236 702788
rect 71872 594856 71924 594862
rect 71872 594798 71924 594804
rect 71780 583024 71832 583030
rect 71780 582966 71832 582972
rect 71884 582162 71912 594798
rect 74632 590708 74684 590714
rect 74632 590650 74684 590656
rect 73344 584112 73396 584118
rect 73344 584054 73396 584060
rect 71792 582134 71912 582162
rect 70412 581862 70702 581890
rect 70964 581874 71300 581890
rect 70952 581868 71300 581874
rect 71004 581862 71300 581868
rect 70952 581810 71004 581816
rect 71792 581754 71820 582134
rect 73356 581890 73384 584054
rect 74644 581890 74672 590650
rect 75196 586514 75224 702782
rect 75104 586486 75224 586514
rect 75104 583953 75132 586486
rect 76576 585342 76604 702986
rect 77956 596174 77984 703190
rect 79324 702636 79376 702642
rect 79324 702578 79376 702584
rect 79336 596174 79364 702578
rect 89180 702434 89208 703520
rect 95148 703180 95200 703186
rect 95148 703122 95200 703128
rect 88352 702406 89208 702434
rect 86960 618316 87012 618322
rect 86960 618258 87012 618264
rect 85580 597576 85632 597582
rect 85580 597518 85632 597524
rect 77956 596146 78076 596174
rect 76564 585336 76616 585342
rect 76564 585278 76616 585284
rect 75090 583944 75146 583953
rect 73278 581862 73384 581890
rect 74566 581862 74672 581890
rect 75012 583902 75090 583930
rect 75012 581754 75040 583902
rect 75090 583879 75146 583888
rect 76576 581890 76604 585278
rect 78048 585274 78076 596146
rect 79244 596146 79364 596174
rect 85592 596174 85620 597518
rect 85592 596146 85712 596174
rect 78036 585268 78088 585274
rect 78036 585210 78088 585216
rect 77852 584044 77904 584050
rect 77852 583986 77904 583992
rect 77864 583778 77892 583986
rect 77852 583772 77904 583778
rect 77852 583714 77904 583720
rect 76748 582616 76800 582622
rect 76748 582558 76800 582564
rect 76498 581862 76604 581890
rect 76760 581890 76788 582558
rect 77864 581890 77892 583714
rect 76760 581862 77096 581890
rect 77786 581862 77892 581890
rect 78048 581890 78076 585210
rect 79244 584050 79272 596146
rect 81808 591320 81860 591326
rect 81808 591262 81860 591268
rect 79324 586628 79376 586634
rect 79324 586570 79376 586576
rect 79232 584044 79284 584050
rect 79232 583986 79284 583992
rect 78680 583840 78732 583846
rect 78680 583782 78732 583788
rect 78692 581890 78720 583782
rect 79336 581890 79364 586570
rect 80612 585200 80664 585206
rect 80612 585142 80664 585148
rect 80624 581890 80652 585142
rect 81820 583817 81848 591262
rect 83188 586696 83240 586702
rect 83188 586638 83240 586644
rect 83004 586560 83056 586566
rect 83004 586502 83056 586508
rect 81900 583908 81952 583914
rect 81900 583850 81952 583856
rect 81438 583808 81494 583817
rect 81438 583743 81494 583752
rect 81806 583808 81862 583817
rect 81806 583743 81862 583752
rect 81452 581890 81480 583743
rect 81912 581890 81940 583850
rect 83016 581890 83044 586502
rect 78048 581862 78384 581890
rect 78692 581862 79028 581890
rect 79336 581862 79672 581890
rect 80624 581862 80960 581890
rect 81452 581862 81604 581890
rect 81912 581862 82248 581890
rect 82938 581862 83044 581890
rect 83200 581890 83228 586638
rect 85304 586560 85356 586566
rect 85304 586502 85356 586508
rect 84476 582548 84528 582554
rect 84476 582490 84528 582496
rect 84488 581890 84516 582490
rect 83200 581862 83536 581890
rect 84488 581862 84824 581890
rect 75460 581800 75512 581806
rect 71792 581726 71944 581754
rect 72252 581738 72588 581754
rect 72240 581732 72588 581738
rect 72292 581726 72588 581732
rect 75012 581726 75164 581754
rect 85316 581754 85344 586502
rect 85684 581890 85712 596146
rect 86972 589014 87000 618258
rect 86960 589008 87012 589014
rect 86960 588950 87012 588956
rect 88248 589008 88300 589014
rect 88248 588950 88300 588956
rect 86972 587926 87000 588950
rect 87696 588600 87748 588606
rect 87696 588542 87748 588548
rect 86960 587920 87012 587926
rect 86960 587862 87012 587868
rect 87708 586634 87736 588542
rect 87696 586628 87748 586634
rect 87696 586570 87748 586576
rect 87708 581890 87736 586570
rect 88260 585138 88288 588950
rect 88352 588606 88380 702406
rect 90364 670744 90416 670750
rect 90364 670686 90416 670692
rect 90376 591326 90404 670686
rect 90364 591320 90416 591326
rect 90364 591262 90416 591268
rect 91468 589348 91520 589354
rect 91468 589290 91520 589296
rect 88340 588600 88392 588606
rect 88340 588542 88392 588548
rect 89628 585200 89680 585206
rect 89628 585142 89680 585148
rect 88248 585132 88300 585138
rect 88248 585074 88300 585080
rect 88246 584080 88302 584089
rect 88246 584015 88302 584024
rect 88260 581890 88288 584015
rect 88982 583944 89038 583953
rect 88982 583879 89038 583888
rect 88996 581890 89024 583879
rect 89640 581890 89668 585142
rect 91374 583808 91430 583817
rect 91374 583743 91430 583752
rect 90272 582616 90324 582622
rect 90272 582558 90324 582564
rect 90284 581890 90312 582558
rect 91008 582548 91060 582554
rect 91008 582490 91060 582496
rect 91020 581890 91048 582490
rect 91388 581890 91416 583743
rect 85684 581862 86112 581890
rect 87446 581862 87736 581890
rect 88090 581862 88288 581890
rect 88734 581862 89024 581890
rect 89378 581862 89668 581890
rect 90022 581862 90312 581890
rect 90666 581862 91048 581890
rect 91310 581862 91416 581890
rect 91480 581890 91508 589290
rect 94872 586696 94924 586702
rect 94872 586638 94924 586644
rect 94136 585268 94188 585274
rect 94136 585210 94188 585216
rect 92848 582684 92900 582690
rect 92848 582626 92900 582632
rect 92860 581890 92888 582626
rect 94148 581890 94176 585210
rect 94884 581890 94912 586638
rect 95160 585342 95188 703122
rect 104808 702976 104860 702982
rect 104808 702918 104860 702924
rect 104820 585478 104848 702918
rect 105464 702434 105492 703520
rect 110328 703112 110380 703118
rect 110328 703054 110380 703060
rect 108948 702568 109000 702574
rect 108948 702510 109000 702516
rect 105464 702406 105584 702434
rect 105556 596174 105584 702406
rect 106280 698964 106332 698970
rect 106280 698906 106332 698912
rect 105556 596146 105676 596174
rect 103520 585472 103572 585478
rect 103520 585414 103572 585420
rect 104808 585472 104860 585478
rect 104808 585414 104860 585420
rect 102416 585404 102468 585410
rect 102416 585346 102468 585352
rect 95148 585336 95200 585342
rect 95148 585278 95200 585284
rect 95160 582162 95188 585278
rect 95424 585132 95476 585138
rect 95424 585074 95476 585080
rect 91480 581862 91908 581890
rect 92598 581862 92888 581890
rect 93886 581862 94176 581890
rect 94530 581862 94912 581890
rect 94976 582134 95188 582162
rect 94976 581754 95004 582134
rect 95436 581890 95464 585074
rect 102428 585070 102456 585346
rect 98736 585064 98788 585070
rect 98736 585006 98788 585012
rect 102416 585064 102468 585070
rect 103532 585018 103560 585414
rect 102416 585006 102468 585012
rect 96528 583908 96580 583914
rect 96528 583850 96580 583856
rect 96540 581890 96568 583850
rect 97448 582752 97500 582758
rect 97448 582694 97500 582700
rect 97460 581890 97488 582694
rect 98748 581890 98776 585006
rect 103348 584990 103560 585018
rect 102600 584112 102652 584118
rect 102600 584054 102652 584060
rect 101312 583976 101364 583982
rect 101312 583918 101364 583924
rect 99288 583840 99340 583846
rect 99288 583782 99340 583788
rect 99300 581890 99328 583782
rect 101324 581890 101352 583918
rect 101862 582448 101918 582457
rect 101862 582383 101918 582392
rect 101876 581890 101904 582383
rect 102612 581890 102640 584054
rect 103348 581890 103376 584990
rect 104624 584044 104676 584050
rect 104624 583986 104676 583992
rect 95436 581862 95772 581890
rect 96462 581862 96568 581890
rect 97106 581862 97488 581890
rect 98394 581862 98776 581890
rect 99038 581862 99328 581890
rect 100970 581862 101352 581890
rect 101614 581862 101904 581890
rect 102258 581862 102640 581890
rect 102902 581862 103376 581890
rect 104440 581800 104492 581806
rect 100574 581768 100630 581777
rect 75512 581748 75808 581754
rect 75460 581742 75808 581748
rect 75472 581726 75808 581742
rect 84028 581738 84180 581754
rect 84016 581732 84180 581738
rect 72240 581674 72292 581680
rect 84068 581726 84180 581732
rect 85316 581726 85468 581754
rect 94976 581726 95128 581754
rect 97750 581738 97948 581754
rect 97750 581732 97960 581738
rect 97750 581726 97908 581732
rect 84016 581674 84068 581680
rect 100326 581726 100574 581754
rect 103546 581738 103928 581754
rect 104190 581748 104440 581754
rect 104190 581742 104492 581748
rect 104636 581754 104664 583986
rect 105544 583772 105596 583778
rect 105544 583714 105596 583720
rect 105556 581890 105584 583714
rect 105478 581862 105584 581890
rect 103546 581732 103940 581738
rect 103546 581726 103888 581732
rect 100574 581703 100630 581712
rect 97908 581674 97960 581680
rect 104190 581726 104480 581742
rect 104636 581726 104788 581754
rect 103888 581674 103940 581680
rect 69768 581318 70058 581346
rect 69768 579086 69796 581318
rect 69756 579080 69808 579086
rect 69756 579022 69808 579028
rect 105648 572898 105676 596146
rect 105636 572892 105688 572898
rect 105636 572834 105688 572840
rect 106186 572792 106242 572801
rect 106186 572727 106242 572736
rect 69756 558204 69808 558210
rect 69756 558146 69808 558152
rect 69768 557534 69796 558146
rect 69768 557506 70164 557534
rect 69202 545184 69258 545193
rect 69202 545119 69258 545128
rect 69664 541680 69716 541686
rect 69664 541622 69716 541628
rect 69296 533384 69348 533390
rect 69296 533326 69348 533332
rect 69202 486024 69258 486033
rect 69202 485959 69258 485968
rect 69110 482896 69166 482905
rect 69110 482831 69166 482840
rect 68926 451888 68982 451897
rect 68926 451823 68982 451832
rect 68756 451246 68876 451274
rect 68756 445097 68784 451246
rect 68742 445088 68798 445097
rect 68742 445023 68798 445032
rect 68388 402946 68692 402974
rect 68664 386050 68692 402946
rect 68834 401704 68890 401713
rect 68834 401639 68890 401648
rect 68744 386300 68796 386306
rect 68744 386242 68796 386248
rect 68756 386209 68784 386242
rect 68742 386200 68798 386209
rect 68742 386135 68798 386144
rect 68664 386022 68784 386050
rect 68756 383722 68784 386022
rect 68848 384849 68876 401639
rect 68834 384840 68890 384849
rect 68834 384775 68890 384784
rect 68744 383716 68796 383722
rect 68744 383658 68796 383664
rect 68756 383489 68784 383658
rect 68742 383480 68798 383489
rect 68742 383415 68798 383424
rect 67638 382528 67694 382537
rect 67638 382463 67694 382472
rect 67652 382294 67680 382463
rect 67640 382288 67692 382294
rect 67640 382230 67692 382236
rect 67640 380860 67692 380866
rect 67640 380802 67692 380808
rect 67652 380769 67680 380802
rect 68008 380792 68060 380798
rect 67638 380760 67694 380769
rect 68008 380734 68060 380740
rect 67638 380695 67694 380704
rect 67638 379808 67694 379817
rect 67638 379743 67694 379752
rect 67652 379574 67680 379743
rect 68020 379681 68048 380734
rect 68006 379672 68062 379681
rect 68006 379607 68062 379616
rect 67640 379568 67692 379574
rect 67640 379510 67692 379516
rect 67640 378820 67692 378826
rect 67640 378762 67692 378768
rect 67652 378729 67680 378762
rect 67638 378720 67694 378729
rect 67638 378655 67694 378664
rect 67638 377088 67694 377097
rect 67638 377023 67694 377032
rect 67652 376786 67680 377023
rect 67640 376780 67692 376786
rect 67640 376722 67692 376728
rect 67640 376644 67692 376650
rect 67640 376586 67692 376592
rect 67652 376009 67680 376586
rect 67638 376000 67694 376009
rect 67638 375935 67694 375944
rect 67640 375896 67692 375902
rect 67640 375838 67692 375844
rect 67652 374678 67680 375838
rect 67640 374672 67692 374678
rect 67638 374640 67640 374649
rect 67692 374640 67694 374649
rect 67638 374575 67694 374584
rect 67640 373992 67692 373998
rect 67640 373934 67692 373940
rect 67652 373289 67680 373934
rect 67638 373280 67694 373289
rect 67638 373215 67694 373224
rect 67640 373176 67692 373182
rect 67640 373118 67692 373124
rect 67652 372473 67680 373118
rect 67638 372464 67694 372473
rect 67638 372399 67694 372408
rect 67640 370660 67692 370666
rect 67640 370602 67692 370608
rect 67652 369753 67680 370602
rect 67732 370592 67784 370598
rect 67732 370534 67784 370540
rect 67744 370297 67772 370534
rect 67730 370288 67786 370297
rect 67730 370223 67786 370232
rect 67638 369744 67694 369753
rect 67638 369679 67694 369688
rect 67640 369164 67692 369170
rect 67640 369106 67692 369112
rect 67652 369073 67680 369106
rect 67638 369064 67694 369073
rect 67638 368999 67694 369008
rect 67916 367872 67968 367878
rect 67916 367814 67968 367820
rect 67928 367441 67956 367814
rect 67914 367432 67970 367441
rect 67914 367367 67970 367376
rect 68742 367432 68798 367441
rect 68742 367367 68798 367376
rect 67638 366480 67694 366489
rect 67638 366415 67694 366424
rect 68468 366444 68520 366450
rect 67652 366382 67680 366415
rect 68468 366386 68520 366392
rect 67640 366376 67692 366382
rect 67640 366318 67692 366324
rect 68480 365809 68508 366386
rect 68466 365800 68522 365809
rect 68466 365735 68522 365744
rect 67732 364336 67784 364342
rect 67732 364278 67784 364284
rect 67638 363760 67694 363769
rect 67638 363695 67694 363704
rect 67652 363662 67680 363695
rect 67640 363656 67692 363662
rect 67744 363633 67772 364278
rect 67640 363598 67692 363604
rect 67730 363624 67786 363633
rect 67730 363559 67786 363568
rect 67638 362400 67694 362409
rect 67560 362358 67638 362386
rect 67362 353424 67418 353433
rect 67362 353359 67418 353368
rect 67376 338910 67404 353359
rect 67364 338904 67416 338910
rect 67364 338846 67416 338852
rect 67560 323649 67588 362358
rect 67638 362335 67694 362344
rect 67640 361548 67692 361554
rect 67640 361490 67692 361496
rect 67652 361321 67680 361490
rect 67638 361312 67694 361321
rect 67638 361247 67694 361256
rect 67640 360868 67692 360874
rect 67640 360810 67692 360816
rect 67652 360641 67680 360810
rect 67638 360632 67694 360641
rect 67638 360567 67694 360576
rect 67638 359544 67694 359553
rect 68480 359514 68508 365735
rect 68560 365016 68612 365022
rect 68560 364958 68612 364964
rect 68572 364721 68600 364958
rect 68558 364712 68614 364721
rect 68558 364647 68614 364656
rect 68572 364334 68600 364647
rect 68572 364306 68692 364334
rect 68560 359576 68612 359582
rect 68560 359518 68612 359524
rect 67638 359479 67640 359488
rect 67692 359479 67694 359488
rect 68468 359508 68520 359514
rect 67640 359450 67692 359456
rect 68468 359450 68520 359456
rect 67638 358184 67694 358193
rect 67638 358119 67694 358128
rect 67652 358086 67680 358119
rect 67640 358080 67692 358086
rect 67640 358022 67692 358028
rect 67638 357504 67694 357513
rect 67638 357439 67640 357448
rect 67692 357439 67694 357448
rect 67640 357410 67692 357416
rect 67638 356960 67694 356969
rect 67638 356895 67694 356904
rect 67652 356726 67680 356895
rect 67640 356720 67692 356726
rect 67640 356662 67692 356668
rect 67640 356040 67692 356046
rect 67640 355982 67692 355988
rect 67652 355881 67680 355982
rect 67638 355872 67694 355881
rect 67638 355807 67694 355816
rect 67638 354784 67694 354793
rect 67638 354719 67640 354728
rect 67692 354719 67694 354728
rect 67640 354690 67692 354696
rect 68572 352753 68600 359518
rect 68558 352744 68614 352753
rect 68558 352679 68614 352688
rect 67640 352640 67692 352646
rect 67638 352608 67640 352617
rect 67692 352608 67694 352617
rect 68572 352578 68600 352679
rect 67638 352543 67694 352552
rect 68560 352572 68612 352578
rect 68560 352514 68612 352520
rect 68006 351248 68062 351257
rect 68006 351183 68008 351192
rect 68060 351183 68062 351192
rect 68008 351154 68060 351160
rect 67638 349888 67694 349897
rect 67638 349823 67640 349832
rect 67692 349823 67694 349832
rect 67640 349794 67692 349800
rect 67638 349208 67694 349217
rect 67638 349143 67640 349152
rect 67692 349143 67694 349152
rect 67640 349114 67692 349120
rect 67638 348528 67694 348537
rect 67638 348463 67640 348472
rect 67692 348463 67694 348472
rect 67640 348434 67692 348440
rect 67640 347744 67692 347750
rect 67640 347686 67692 347692
rect 67652 347313 67680 347686
rect 67638 347304 67694 347313
rect 67638 347239 67694 347248
rect 67638 345672 67694 345681
rect 67638 345607 67694 345616
rect 67652 345166 67680 345607
rect 67640 345160 67692 345166
rect 67640 345102 67692 345108
rect 68008 345024 68060 345030
rect 68664 345014 68692 364306
rect 68008 344966 68060 344972
rect 68572 344986 68692 345014
rect 67638 344448 67694 344457
rect 67638 344383 67694 344392
rect 67652 343670 67680 344383
rect 68020 344321 68048 344966
rect 68006 344312 68062 344321
rect 68006 344247 68062 344256
rect 67640 343664 67692 343670
rect 67640 343606 67692 343612
rect 67638 342952 67694 342961
rect 67638 342887 67694 342896
rect 67652 342310 67680 342887
rect 67640 342304 67692 342310
rect 67640 342246 67692 342252
rect 67638 341728 67694 341737
rect 67638 341663 67694 341672
rect 67652 340950 67680 341663
rect 67640 340944 67692 340950
rect 67640 340886 67692 340892
rect 68572 337414 68600 344986
rect 68652 341624 68704 341630
rect 68650 341592 68652 341601
rect 68704 341592 68706 341601
rect 68650 341527 68706 341536
rect 68652 340876 68704 340882
rect 68652 340818 68704 340824
rect 68664 340649 68692 340818
rect 68650 340640 68706 340649
rect 68650 340575 68706 340584
rect 68560 337408 68612 337414
rect 68560 337350 68612 337356
rect 68756 333266 68784 367367
rect 68940 359582 68968 451823
rect 69124 439074 69152 482831
rect 69216 439618 69244 485959
rect 69308 460934 69336 533326
rect 69676 497486 69704 541622
rect 69768 540110 70058 540138
rect 69768 533390 69796 540110
rect 70136 536858 70164 557506
rect 105726 543824 105782 543833
rect 105726 543759 105782 543768
rect 70412 540110 70702 540138
rect 70124 536852 70176 536858
rect 70124 536794 70176 536800
rect 69756 533384 69808 533390
rect 69756 533326 69808 533332
rect 70412 529310 70440 540110
rect 71332 536110 71360 540138
rect 71320 536104 71372 536110
rect 71320 536046 71372 536052
rect 70400 529304 70452 529310
rect 70400 529246 70452 529252
rect 71976 526454 72004 540138
rect 72620 537606 72648 540138
rect 73160 538960 73212 538966
rect 73160 538902 73212 538908
rect 73172 538082 73200 538902
rect 73160 538076 73212 538082
rect 73160 538018 73212 538024
rect 72608 537600 72660 537606
rect 72608 537542 72660 537548
rect 73172 536926 73200 538018
rect 73160 536920 73212 536926
rect 73160 536862 73212 536868
rect 72424 534948 72476 534954
rect 72424 534890 72476 534896
rect 71964 526448 72016 526454
rect 71964 526390 72016 526396
rect 69664 497480 69716 497486
rect 69664 497422 69716 497428
rect 72436 493746 72464 534890
rect 73264 534750 73292 540138
rect 73804 536920 73856 536926
rect 73804 536862 73856 536868
rect 73252 534744 73304 534750
rect 73252 534686 73304 534692
rect 73252 495576 73304 495582
rect 73252 495518 73304 495524
rect 70860 493740 70912 493746
rect 70860 493682 70912 493688
rect 72424 493740 72476 493746
rect 72424 493682 72476 493688
rect 70032 492856 70084 492862
rect 70032 492798 70084 492804
rect 69756 490612 69808 490618
rect 69756 490554 69808 490560
rect 69768 489977 69796 490554
rect 69754 489968 69810 489977
rect 70044 489940 70072 492798
rect 70400 492040 70452 492046
rect 70400 491982 70452 491988
rect 70412 489954 70440 491982
rect 70412 489926 70656 489954
rect 69754 489903 69810 489912
rect 70872 489870 70900 493682
rect 71780 493332 71832 493338
rect 71780 493274 71832 493280
rect 70952 491360 71004 491366
rect 70952 491302 71004 491308
rect 70964 489954 70992 491302
rect 71792 489954 71820 493274
rect 72240 491972 72292 491978
rect 72240 491914 72292 491920
rect 72252 489954 72280 491914
rect 70964 489926 71300 489954
rect 71792 489926 71944 489954
rect 72252 489926 72588 489954
rect 73264 489940 73292 495518
rect 73816 490822 73844 536862
rect 73908 536790 73936 540138
rect 73896 536784 73948 536790
rect 73896 536726 73948 536732
rect 74552 529242 74580 540138
rect 75196 534886 75224 540138
rect 76467 540110 76512 540138
rect 75920 536852 75972 536858
rect 75920 536794 75972 536800
rect 75184 534880 75236 534886
rect 75184 534822 75236 534828
rect 74540 529236 74592 529242
rect 74540 529178 74592 529184
rect 75828 497480 75880 497486
rect 75828 497422 75880 497428
rect 74540 495508 74592 495514
rect 74540 495450 74592 495456
rect 73804 490816 73856 490822
rect 73804 490758 73856 490764
rect 74552 489940 74580 495450
rect 74816 493400 74868 493406
rect 74816 493342 74868 493348
rect 74828 489954 74856 493342
rect 74828 489926 75164 489954
rect 75840 489940 75868 497422
rect 75932 490210 75960 536794
rect 76484 532166 76512 540110
rect 76472 532160 76524 532166
rect 76472 532102 76524 532108
rect 77128 529378 77156 540138
rect 77772 534954 77800 540138
rect 77760 534948 77812 534954
rect 77760 534890 77812 534896
rect 78416 534818 78444 540138
rect 78404 534812 78456 534818
rect 78404 534754 78456 534760
rect 79060 532030 79088 540138
rect 79324 537804 79376 537810
rect 79324 537746 79376 537752
rect 79048 532024 79100 532030
rect 79048 531966 79100 531972
rect 77116 529372 77168 529378
rect 77116 529314 77168 529320
rect 76104 495644 76156 495650
rect 76104 495586 76156 495592
rect 75920 490204 75972 490210
rect 75920 490146 75972 490152
rect 76116 489954 76144 495586
rect 79336 494086 79364 537746
rect 79704 499574 79732 540138
rect 80348 538121 80376 540138
rect 80334 538112 80390 538121
rect 80334 538047 80390 538056
rect 80348 537441 80376 538047
rect 80334 537432 80390 537441
rect 80334 537367 80390 537376
rect 79612 499546 79732 499574
rect 79324 494080 79376 494086
rect 79324 494022 79376 494028
rect 77760 492652 77812 492658
rect 77760 492594 77812 492600
rect 77070 490204 77122 490210
rect 77070 490146 77122 490152
rect 77082 489954 77110 490146
rect 76116 489926 76452 489954
rect 77082 489940 77340 489954
rect 77772 489940 77800 492594
rect 79612 490754 79640 499546
rect 80992 496126 81020 540138
rect 81636 537674 81664 540138
rect 82907 540110 82952 540138
rect 82268 538892 82320 538898
rect 82268 538834 82320 538840
rect 82280 538014 82308 538834
rect 82268 538008 82320 538014
rect 82268 537950 82320 537956
rect 81624 537668 81676 537674
rect 81624 537610 81676 537616
rect 82280 536858 82308 537950
rect 82924 537538 82952 540110
rect 82912 537532 82964 537538
rect 82912 537474 82964 537480
rect 82268 536852 82320 536858
rect 82268 536794 82320 536800
rect 82728 536852 82780 536858
rect 82728 536794 82780 536800
rect 81440 498228 81492 498234
rect 81440 498170 81492 498176
rect 81452 497486 81480 498170
rect 81440 497480 81492 497486
rect 81440 497422 81492 497428
rect 80980 496120 81032 496126
rect 80980 496062 81032 496068
rect 82268 494896 82320 494902
rect 82268 494838 82320 494844
rect 80980 494760 81032 494766
rect 80980 494702 81032 494708
rect 79968 494080 80020 494086
rect 79968 494022 80020 494028
rect 79692 493332 79744 493338
rect 79692 493274 79744 493280
rect 79600 490748 79652 490754
rect 79600 490690 79652 490696
rect 78036 490680 78088 490686
rect 78036 490622 78088 490628
rect 78048 489954 78076 490622
rect 77096 489938 77340 489940
rect 77096 489932 77352 489938
rect 77096 489926 77300 489932
rect 78048 489926 78384 489954
rect 79704 489940 79732 493274
rect 79980 492658 80008 494022
rect 79968 492652 80020 492658
rect 79968 492594 80020 492600
rect 80060 491428 80112 491434
rect 80060 491370 80112 491376
rect 80072 489954 80100 491370
rect 80072 489926 80316 489954
rect 80992 489940 81020 494702
rect 81624 493468 81676 493474
rect 81624 493410 81676 493416
rect 81636 489940 81664 493410
rect 82280 489940 82308 494838
rect 82740 494834 82768 536794
rect 83568 532098 83596 540138
rect 84108 536852 84160 536858
rect 84108 536794 84160 536800
rect 83556 532092 83608 532098
rect 83556 532034 83608 532040
rect 84120 500410 84148 536794
rect 84108 500404 84160 500410
rect 84108 500346 84160 500352
rect 84212 498846 84240 540138
rect 84856 536926 84884 540138
rect 84844 536920 84896 536926
rect 84844 536862 84896 536868
rect 85500 536858 85528 540138
rect 85488 536852 85540 536858
rect 85488 536794 85540 536800
rect 84200 498840 84252 498846
rect 86144 498817 86172 540138
rect 84200 498782 84252 498788
rect 86130 498808 86186 498817
rect 86130 498743 86186 498752
rect 83832 497480 83884 497486
rect 83832 497422 83884 497428
rect 83844 495446 83872 497422
rect 86788 496233 86816 540138
rect 87432 497622 87460 540138
rect 88076 538150 88104 540138
rect 89347 540110 89392 540138
rect 88064 538144 88116 538150
rect 88064 538086 88116 538092
rect 89364 532098 89392 540110
rect 90008 534750 90036 540138
rect 90364 536920 90416 536926
rect 90364 536862 90416 536868
rect 89996 534744 90048 534750
rect 89996 534686 90048 534692
rect 89352 532092 89404 532098
rect 89352 532034 89404 532040
rect 87420 497616 87472 497622
rect 87420 497558 87472 497564
rect 90376 497457 90404 536862
rect 90652 497554 90680 540138
rect 91296 538082 91324 540138
rect 91284 538076 91336 538082
rect 91284 538018 91336 538024
rect 91100 500336 91152 500342
rect 91100 500278 91152 500284
rect 91112 499574 91140 500278
rect 91940 500274 91968 540138
rect 92584 532001 92612 540138
rect 92570 531992 92626 532001
rect 92570 531927 92626 531936
rect 93228 500478 93256 540138
rect 93872 534818 93900 540138
rect 94516 537742 94544 540138
rect 95787 540110 95832 540138
rect 95056 538960 95108 538966
rect 95056 538902 95108 538908
rect 94504 537736 94556 537742
rect 94504 537678 94556 537684
rect 93860 534812 93912 534818
rect 93860 534754 93912 534760
rect 93768 532024 93820 532030
rect 93768 531966 93820 531972
rect 93216 500472 93268 500478
rect 93216 500414 93268 500420
rect 91744 500268 91796 500274
rect 91744 500210 91796 500216
rect 91928 500268 91980 500274
rect 91928 500210 91980 500216
rect 91112 499546 91508 499574
rect 90640 497548 90692 497554
rect 90640 497490 90692 497496
rect 90362 497448 90418 497457
rect 90362 497383 90418 497392
rect 86774 496224 86830 496233
rect 86774 496159 86830 496168
rect 88248 496188 88300 496194
rect 88248 496130 88300 496136
rect 83832 495440 83884 495446
rect 83832 495382 83884 495388
rect 82728 494828 82780 494834
rect 82728 494770 82780 494776
rect 82912 493400 82964 493406
rect 82912 493342 82964 493348
rect 82924 489940 82952 493342
rect 83844 489954 83872 495382
rect 85488 494216 85540 494222
rect 85488 494158 85540 494164
rect 84844 491564 84896 491570
rect 84844 491506 84896 491512
rect 83582 489926 83872 489954
rect 84856 489940 84884 491506
rect 85500 489940 85528 494158
rect 88260 493474 88288 496130
rect 89626 496088 89682 496097
rect 89626 496023 89682 496032
rect 89640 494222 89668 496023
rect 89628 494216 89680 494222
rect 89628 494158 89680 494164
rect 88248 493468 88300 493474
rect 88248 493410 88300 493416
rect 90272 493468 90324 493474
rect 90272 493410 90324 493416
rect 90284 492794 90312 493410
rect 90272 492788 90324 492794
rect 90272 492730 90324 492736
rect 89720 492720 89772 492726
rect 89720 492662 89772 492668
rect 88708 491632 88760 491638
rect 88708 491574 88760 491580
rect 86776 491428 86828 491434
rect 86776 491370 86828 491376
rect 86132 491360 86184 491366
rect 86132 491302 86184 491308
rect 86144 489940 86172 491302
rect 86788 489940 86816 491370
rect 87694 490648 87750 490657
rect 87694 490583 87750 490592
rect 87708 489954 87736 490583
rect 88248 490000 88300 490006
rect 87446 489926 87736 489954
rect 88090 489948 88248 489954
rect 88090 489942 88300 489948
rect 88090 489926 88288 489942
rect 88720 489940 88748 491574
rect 89732 489954 89760 492662
rect 90284 489954 90312 492730
rect 91284 492652 91336 492658
rect 91284 492594 91336 492600
rect 89732 489926 89976 489954
rect 90284 489926 90620 489954
rect 91296 489940 91324 492594
rect 91480 489954 91508 499546
rect 91756 492658 91784 500210
rect 93216 496120 93268 496126
rect 93216 496062 93268 496068
rect 91744 492652 91796 492658
rect 91744 492594 91796 492600
rect 92848 490680 92900 490686
rect 92848 490622 92900 490628
rect 92860 489954 92888 490622
rect 91480 489926 91908 489954
rect 92598 489926 92888 489954
rect 93228 489940 93256 496062
rect 93780 491366 93808 531966
rect 95068 499574 95096 538902
rect 95148 538892 95200 538898
rect 95148 538834 95200 538840
rect 94976 499546 95096 499574
rect 93768 491360 93820 491366
rect 93820 491308 93900 491314
rect 93768 491302 93900 491308
rect 93780 491286 93900 491302
rect 93872 490822 93900 491286
rect 93860 490816 93912 490822
rect 93860 490758 93912 490764
rect 94976 490618 95004 499546
rect 95160 495802 95188 538834
rect 95804 537674 95832 540110
rect 95792 537668 95844 537674
rect 95792 537610 95844 537616
rect 95068 495774 95188 495802
rect 95068 490657 95096 495774
rect 96448 495038 96476 540138
rect 97092 536897 97120 540138
rect 97078 536888 97134 536897
rect 97078 536823 97134 536832
rect 96436 495032 96488 495038
rect 96436 494974 96488 494980
rect 97736 494018 97764 540138
rect 98380 538218 98408 540138
rect 98368 538214 98420 538218
rect 98368 538212 98776 538214
rect 98420 538186 98776 538212
rect 98368 538154 98420 538160
rect 97908 536104 97960 536110
rect 97908 536046 97960 536052
rect 97724 494012 97776 494018
rect 97724 493954 97776 493960
rect 95240 493536 95292 493542
rect 95240 493478 95292 493484
rect 95252 492674 95280 493478
rect 95790 493368 95846 493377
rect 95790 493303 95846 493312
rect 95160 492646 95280 492674
rect 95054 490648 95110 490657
rect 94136 490612 94188 490618
rect 94136 490554 94188 490560
rect 94964 490612 95016 490618
rect 95054 490583 95110 490592
rect 94964 490554 95016 490560
rect 94148 489954 94176 490554
rect 93886 489926 94176 489954
rect 95160 489940 95188 492646
rect 95804 489940 95832 493303
rect 97724 492312 97776 492318
rect 97724 492254 97776 492260
rect 96436 492108 96488 492114
rect 96436 492050 96488 492056
rect 96448 489940 96476 492050
rect 97078 490512 97134 490521
rect 97078 490447 97134 490456
rect 97092 489940 97120 490447
rect 97736 489940 97764 492254
rect 97920 492114 97948 536046
rect 98644 534880 98696 534886
rect 98644 534822 98696 534828
rect 97908 492108 97960 492114
rect 97908 492050 97960 492056
rect 98656 491298 98684 534822
rect 98748 494970 98776 538186
rect 99024 538014 99052 540138
rect 99012 538008 99064 538014
rect 99012 537950 99064 537956
rect 99288 534948 99340 534954
rect 99288 534890 99340 534896
rect 98736 494964 98788 494970
rect 98736 494906 98788 494912
rect 99300 492318 99328 534890
rect 99668 528554 99696 540138
rect 99392 528526 99696 528554
rect 99288 492312 99340 492318
rect 99288 492254 99340 492260
rect 99300 492046 99328 492254
rect 99288 492040 99340 492046
rect 99288 491982 99340 491988
rect 99012 491496 99064 491502
rect 99012 491438 99064 491444
rect 98644 491292 98696 491298
rect 98644 491234 98696 491240
rect 99024 489940 99052 491438
rect 77300 489874 77352 489880
rect 69848 489864 69900 489870
rect 69848 489806 69900 489812
rect 70860 489864 70912 489870
rect 98736 489864 98788 489870
rect 70860 489806 70912 489812
rect 98394 489812 98736 489818
rect 98394 489806 98788 489812
rect 99288 489864 99340 489870
rect 99288 489806 99340 489812
rect 69860 489161 69888 489806
rect 98394 489790 98776 489806
rect 69846 489152 69902 489161
rect 69846 489087 69902 489096
rect 99300 488578 99328 489806
rect 99288 488572 99340 488578
rect 99288 488514 99340 488520
rect 99392 460934 99420 528526
rect 99656 491428 99708 491434
rect 99656 491370 99708 491376
rect 99668 489940 99696 491370
rect 100024 490816 100076 490822
rect 100024 490758 100076 490764
rect 69308 460906 69704 460934
rect 99392 460906 99512 460934
rect 69676 440722 69704 460906
rect 99378 443728 99434 443737
rect 99378 443663 99434 443672
rect 69676 440694 70058 440722
rect 72344 440706 72634 440722
rect 79336 440706 79824 440722
rect 71780 440700 71832 440706
rect 69204 439612 69256 439618
rect 69204 439554 69256 439560
rect 69112 439068 69164 439074
rect 69112 439010 69164 439016
rect 69112 437504 69164 437510
rect 69112 437446 69164 437452
rect 69124 437374 69152 437446
rect 69112 437368 69164 437374
rect 69112 437310 69164 437316
rect 69124 436529 69152 437310
rect 69110 436520 69166 436529
rect 69110 436455 69166 436464
rect 69676 431954 69704 440694
rect 71780 440642 71832 440648
rect 72332 440700 72634 440706
rect 72384 440694 72634 440700
rect 79324 440700 79824 440706
rect 72332 440642 72384 440648
rect 79376 440694 79824 440700
rect 93886 440706 94176 440722
rect 93886 440700 94188 440706
rect 93886 440694 94136 440700
rect 79324 440642 79376 440648
rect 70400 438660 70452 438666
rect 70400 438602 70452 438608
rect 70412 437238 70440 438602
rect 70400 437232 70452 437238
rect 70400 437174 70452 437180
rect 70412 436121 70440 437174
rect 70398 436112 70454 436121
rect 70398 436047 70454 436056
rect 70688 434654 70716 440028
rect 71042 438968 71098 438977
rect 71042 438903 71098 438912
rect 70676 434648 70728 434654
rect 70676 434590 70728 434596
rect 69308 431926 69704 431954
rect 69112 375352 69164 375358
rect 69112 375294 69164 375300
rect 69124 374241 69152 375294
rect 69110 374232 69166 374241
rect 69110 374167 69166 374176
rect 68928 359576 68980 359582
rect 68928 359518 68980 359524
rect 68836 359508 68888 359514
rect 68836 359450 68888 359456
rect 68744 333260 68796 333266
rect 68744 333202 68796 333208
rect 67546 323640 67602 323649
rect 67546 323575 67602 323584
rect 67548 320952 67600 320958
rect 67548 320894 67600 320900
rect 67456 313948 67508 313954
rect 67456 313890 67508 313896
rect 67270 312624 67326 312633
rect 67270 312559 67326 312568
rect 66168 311908 66220 311914
rect 66168 311850 66220 311856
rect 66076 298308 66128 298314
rect 66076 298250 66128 298256
rect 65982 296032 66038 296041
rect 65982 295967 66038 295976
rect 65524 294092 65576 294098
rect 65524 294034 65576 294040
rect 65536 292534 65564 294034
rect 65524 292528 65576 292534
rect 65524 292470 65576 292476
rect 66088 288318 66116 298250
rect 66180 288386 66208 311850
rect 67468 291145 67496 313890
rect 67454 291136 67510 291145
rect 67454 291071 67510 291080
rect 66902 289232 66958 289241
rect 66902 289167 66958 289176
rect 66168 288380 66220 288386
rect 66168 288322 66220 288328
rect 66076 288312 66128 288318
rect 66076 288254 66128 288260
rect 64604 273284 64656 273290
rect 64604 273226 64656 273232
rect 64512 248532 64564 248538
rect 64512 248474 64564 248480
rect 64524 178770 64552 248474
rect 64616 194138 64644 273226
rect 65984 271992 66036 271998
rect 65984 271934 66036 271940
rect 64696 271924 64748 271930
rect 64696 271866 64748 271872
rect 64604 194132 64656 194138
rect 64604 194074 64656 194080
rect 64708 182918 64736 271866
rect 65892 249076 65944 249082
rect 65892 249018 65944 249024
rect 64788 244316 64840 244322
rect 64788 244258 64840 244264
rect 64800 239494 64828 244258
rect 64788 239488 64840 239494
rect 64788 239430 64840 239436
rect 65904 196722 65932 249018
rect 65996 224262 66024 271934
rect 66916 262886 66944 289167
rect 67560 285433 67588 320894
rect 68848 320890 68876 359450
rect 68926 351248 68982 351257
rect 68926 351183 68982 351192
rect 68836 320884 68888 320890
rect 68836 320826 68888 320832
rect 68940 319462 68968 351183
rect 69020 340060 69072 340066
rect 69020 340002 69072 340008
rect 68928 319456 68980 319462
rect 68928 319398 68980 319404
rect 69032 300150 69060 340002
rect 69124 311137 69152 374167
rect 69308 364334 69336 431926
rect 71056 404326 71084 438903
rect 71332 438190 71360 440028
rect 71320 438184 71372 438190
rect 71320 438126 71372 438132
rect 70400 404320 70452 404326
rect 70400 404262 70452 404268
rect 71044 404320 71096 404326
rect 71044 404262 71096 404268
rect 70412 403034 70440 404262
rect 70400 403028 70452 403034
rect 70400 402970 70452 402976
rect 71792 402974 71820 440642
rect 71976 431954 72004 440028
rect 73264 437510 73292 440028
rect 73804 439068 73856 439074
rect 73804 439010 73856 439016
rect 73252 437504 73304 437510
rect 73252 437446 73304 437452
rect 71884 431934 72004 431954
rect 71872 431928 72004 431934
rect 71924 431926 72004 431928
rect 71872 431870 71924 431876
rect 70308 390040 70360 390046
rect 70308 389982 70360 389988
rect 69848 389972 69900 389978
rect 69848 389914 69900 389920
rect 69664 387388 69716 387394
rect 69664 387330 69716 387336
rect 69676 367810 69704 387330
rect 69860 385778 69888 389914
rect 70216 387864 70268 387870
rect 70216 387806 70268 387812
rect 70228 385914 70256 387806
rect 70058 385886 70256 385914
rect 69768 385750 69888 385778
rect 69768 370530 69796 385750
rect 70320 376038 70348 389982
rect 70412 385914 70440 402970
rect 71792 402946 71912 402974
rect 71780 389224 71832 389230
rect 71780 389166 71832 389172
rect 71792 385914 71820 389166
rect 71884 387326 71912 402946
rect 72424 390584 72476 390590
rect 72424 390526 72476 390532
rect 72436 389162 72464 390526
rect 72424 389156 72476 389162
rect 72424 389098 72476 389104
rect 71872 387320 71924 387326
rect 71872 387262 71924 387268
rect 72436 385914 72464 389098
rect 73816 388142 73844 439010
rect 73908 438258 73936 440028
rect 73896 438252 73948 438258
rect 73896 438194 73948 438200
rect 74552 434722 74580 440028
rect 75184 438864 75236 438870
rect 75184 438806 75236 438812
rect 75196 438161 75224 438806
rect 75182 438152 75238 438161
rect 75182 438087 75238 438096
rect 75840 437306 75868 440028
rect 74632 437300 74684 437306
rect 74632 437242 74684 437248
rect 75828 437300 75880 437306
rect 75828 437242 75880 437248
rect 74540 434716 74592 434722
rect 74540 434658 74592 434664
rect 74644 431954 74672 437242
rect 75184 436756 75236 436762
rect 75184 436698 75236 436704
rect 74552 431926 74672 431954
rect 74552 392698 74580 431926
rect 75196 402974 75224 436698
rect 76484 434586 76512 440028
rect 76564 439612 76616 439618
rect 76564 439554 76616 439560
rect 76472 434580 76524 434586
rect 76472 434522 76524 434528
rect 74828 402946 75224 402974
rect 76576 402974 76604 439554
rect 77128 438666 77156 440028
rect 77312 440014 77786 440042
rect 78430 440014 78628 440042
rect 77116 438660 77168 438666
rect 77116 438602 77168 438608
rect 77312 434625 77340 440014
rect 78600 436014 78628 440014
rect 79060 437442 79088 440028
rect 79324 439544 79376 439550
rect 79324 439486 79376 439492
rect 78680 437436 78732 437442
rect 78680 437378 78732 437384
rect 79048 437436 79100 437442
rect 79048 437378 79100 437384
rect 78588 436008 78640 436014
rect 78588 435950 78640 435956
rect 77944 435396 77996 435402
rect 77944 435338 77996 435344
rect 77298 434616 77354 434625
rect 77298 434551 77354 434560
rect 76576 402946 76696 402974
rect 74828 401674 74856 402946
rect 74816 401668 74868 401674
rect 74816 401610 74868 401616
rect 74540 392692 74592 392698
rect 74540 392634 74592 392640
rect 73528 388136 73580 388142
rect 73528 388078 73580 388084
rect 73804 388136 73856 388142
rect 73804 388078 73856 388084
rect 73540 385914 73568 388078
rect 74630 387968 74686 387977
rect 74630 387903 74686 387912
rect 74644 385914 74672 387903
rect 70412 385886 70702 385914
rect 71792 385886 71990 385914
rect 72436 385886 72634 385914
rect 73278 385886 73568 385914
rect 74566 385886 74672 385914
rect 74828 385914 74856 401610
rect 75460 391264 75512 391270
rect 75460 391206 75512 391212
rect 75472 390658 75500 391206
rect 75460 390652 75512 390658
rect 75460 390594 75512 390600
rect 75472 385914 75500 390594
rect 76668 386442 76696 402946
rect 77312 398138 77340 434551
rect 77300 398132 77352 398138
rect 77300 398074 77352 398080
rect 77956 397458 77984 435338
rect 78600 432002 78628 435950
rect 78588 431996 78640 432002
rect 78588 431938 78640 431944
rect 77944 397452 77996 397458
rect 77944 397394 77996 397400
rect 77956 390726 77984 397394
rect 77944 390720 77996 390726
rect 77944 390662 77996 390668
rect 76656 386436 76708 386442
rect 76656 386378 76708 386384
rect 76668 385914 76696 386378
rect 77956 385914 77984 390662
rect 78034 387832 78090 387841
rect 78034 387767 78090 387776
rect 74828 385886 75210 385914
rect 75472 385886 75854 385914
rect 76668 385886 77142 385914
rect 77786 385886 77984 385914
rect 78048 385914 78076 387767
rect 78692 387394 78720 437378
rect 79336 390046 79364 439486
rect 79796 439074 79824 440694
rect 79784 439068 79836 439074
rect 79784 439010 79836 439016
rect 80992 439006 81020 440028
rect 81452 440014 81650 440042
rect 81452 439550 81480 440014
rect 81440 439544 81492 439550
rect 81440 439486 81492 439492
rect 80980 439000 81032 439006
rect 80980 438942 81032 438948
rect 82280 438870 82308 440028
rect 82820 439068 82872 439074
rect 82820 439010 82872 439016
rect 82268 438864 82320 438870
rect 82268 438806 82320 438812
rect 80152 431996 80204 432002
rect 80152 431938 80204 431944
rect 82832 431954 82860 439010
rect 82924 438802 82952 440028
rect 82912 438796 82964 438802
rect 82912 438738 82964 438744
rect 83568 438734 83596 440028
rect 84212 438802 84240 440028
rect 84200 438796 84252 438802
rect 84200 438738 84252 438744
rect 83556 438728 83608 438734
rect 84856 438705 84884 440028
rect 86144 438870 86172 440028
rect 86132 438864 86184 438870
rect 86132 438806 86184 438812
rect 85580 438796 85632 438802
rect 85580 438738 85632 438744
rect 83556 438670 83608 438676
rect 84198 438696 84254 438705
rect 84198 438631 84254 438640
rect 84842 438696 84898 438705
rect 84842 438631 84898 438640
rect 84212 438002 84240 438631
rect 85592 438190 85620 438738
rect 85580 438184 85632 438190
rect 85580 438126 85632 438132
rect 84120 437974 84240 438002
rect 79324 390040 79376 390046
rect 79324 389982 79376 389988
rect 79324 389292 79376 389298
rect 79324 389234 79376 389240
rect 78680 387388 78732 387394
rect 78680 387330 78732 387336
rect 79336 385914 79364 389234
rect 80060 387932 80112 387938
rect 80060 387874 80112 387880
rect 80072 385914 80100 387874
rect 80164 386034 80192 431938
rect 82832 431926 82952 431954
rect 82820 395412 82872 395418
rect 82820 395354 82872 395360
rect 81440 395344 81492 395350
rect 81440 395286 81492 395292
rect 81452 390726 81480 395286
rect 82832 394806 82860 395354
rect 82820 394800 82872 394806
rect 82820 394742 82872 394748
rect 82924 393990 82952 431926
rect 84120 396846 84148 437974
rect 85028 437504 85080 437510
rect 84198 437472 84254 437481
rect 84198 437407 84254 437416
rect 85026 437472 85028 437481
rect 85080 437472 85082 437481
rect 85026 437407 85082 437416
rect 84108 396840 84160 396846
rect 84108 396782 84160 396788
rect 84212 395486 84240 437407
rect 85120 399492 85172 399498
rect 85120 399434 85172 399440
rect 84200 395480 84252 395486
rect 84200 395422 84252 395428
rect 83096 394800 83148 394806
rect 83096 394742 83148 394748
rect 82912 393984 82964 393990
rect 82912 393926 82964 393932
rect 83002 392592 83058 392601
rect 83002 392527 83058 392536
rect 81440 390720 81492 390726
rect 81440 390662 81492 390668
rect 82544 390720 82596 390726
rect 82544 390662 82596 390668
rect 80612 387252 80664 387258
rect 80612 387194 80664 387200
rect 80152 386028 80204 386034
rect 80152 385970 80204 385976
rect 80624 385914 80652 387194
rect 82556 385914 82584 390662
rect 83016 385914 83044 392527
rect 78048 385886 78430 385914
rect 79336 385886 79718 385914
rect 80072 385886 80362 385914
rect 80624 385886 81006 385914
rect 82294 385886 82584 385914
rect 82938 385886 83044 385914
rect 83108 385914 83136 394742
rect 84200 394732 84252 394738
rect 84200 394674 84252 394680
rect 84212 386050 84240 394674
rect 85132 393378 85160 399434
rect 85120 393372 85172 393378
rect 85120 393314 85172 393320
rect 84212 386022 84424 386050
rect 84396 385914 84424 386022
rect 85132 385914 85160 393314
rect 85592 389978 85620 438126
rect 86788 437510 86816 440028
rect 87432 438326 87460 440028
rect 87420 438320 87472 438326
rect 87420 438262 87472 438268
rect 88076 437510 88104 440028
rect 88720 439006 88748 440028
rect 88708 439000 88760 439006
rect 88708 438942 88760 438948
rect 88248 438660 88300 438666
rect 88248 438602 88300 438608
rect 88260 438326 88288 438602
rect 88248 438320 88300 438326
rect 88248 438262 88300 438268
rect 86776 437504 86828 437510
rect 86776 437446 86828 437452
rect 88064 437504 88116 437510
rect 88064 437446 88116 437452
rect 86224 399560 86276 399566
rect 86224 399502 86276 399508
rect 85580 389972 85632 389978
rect 85580 389914 85632 389920
rect 86236 386481 86264 399502
rect 88260 393990 88288 438262
rect 89364 437306 89392 440028
rect 89628 437504 89680 437510
rect 89628 437446 89680 437452
rect 89352 437300 89404 437306
rect 89352 437242 89404 437248
rect 89536 437300 89588 437306
rect 89536 437242 89588 437248
rect 89548 399634 89576 437242
rect 89640 436014 89668 437446
rect 90008 437442 90036 440028
rect 91296 438802 91324 440028
rect 91756 440014 91954 440042
rect 91284 438796 91336 438802
rect 91284 438738 91336 438744
rect 89996 437436 90048 437442
rect 89996 437378 90048 437384
rect 90364 437436 90416 437442
rect 90364 437378 90416 437384
rect 89628 436008 89680 436014
rect 89628 435950 89680 435956
rect 89536 399628 89588 399634
rect 89536 399570 89588 399576
rect 88340 396772 88392 396778
rect 88340 396714 88392 396720
rect 88352 396098 88380 396714
rect 88340 396092 88392 396098
rect 88340 396034 88392 396040
rect 88248 393984 88300 393990
rect 88248 393926 88300 393932
rect 88248 388544 88300 388550
rect 88248 388486 88300 388492
rect 87052 386504 87104 386510
rect 86222 386472 86278 386481
rect 87052 386446 87104 386452
rect 86222 386407 86278 386416
rect 86236 385914 86264 386407
rect 83108 385886 83582 385914
rect 84396 385886 84870 385914
rect 85132 385886 85514 385914
rect 86158 385886 86264 385914
rect 87064 385914 87092 386446
rect 88260 385914 88288 388486
rect 87064 385886 87446 385914
rect 88090 385886 88288 385914
rect 88352 385914 88380 396034
rect 89640 387258 89668 435950
rect 89720 396908 89772 396914
rect 89720 396850 89772 396856
rect 89732 395486 89760 396850
rect 89720 395480 89772 395486
rect 89720 395422 89772 395428
rect 90272 388612 90324 388618
rect 90272 388554 90324 388560
rect 89628 387252 89680 387258
rect 89628 387194 89680 387200
rect 90284 385914 90312 388554
rect 90376 387190 90404 437378
rect 91756 436082 91784 440014
rect 92584 436082 92612 440028
rect 93228 437238 93256 440028
rect 93964 438530 93992 440694
rect 94136 440642 94188 440648
rect 97448 440700 97500 440706
rect 97448 440642 97500 440648
rect 95332 440224 95384 440230
rect 95174 440172 95332 440178
rect 95174 440166 95384 440172
rect 95174 440150 95372 440166
rect 97460 440042 97488 440642
rect 97908 440156 97960 440162
rect 97908 440098 97960 440104
rect 97920 440042 97948 440098
rect 94530 440014 95004 440042
rect 97106 440028 97488 440042
rect 97750 440028 97948 440042
rect 94504 438864 94556 438870
rect 94504 438806 94556 438812
rect 93584 438524 93636 438530
rect 93584 438466 93636 438472
rect 93952 438524 94004 438530
rect 93952 438466 94004 438472
rect 93216 437232 93268 437238
rect 93216 437174 93268 437180
rect 91744 436076 91796 436082
rect 91744 436018 91796 436024
rect 92572 436076 92624 436082
rect 92572 436018 92624 436024
rect 91756 398138 91784 436018
rect 93596 403714 93624 438466
rect 93676 437232 93728 437238
rect 93676 437174 93728 437180
rect 93584 403708 93636 403714
rect 93584 403650 93636 403656
rect 93688 399566 93716 437174
rect 93768 436076 93820 436082
rect 93768 436018 93820 436024
rect 93676 399560 93728 399566
rect 93676 399502 93728 399508
rect 92664 399492 92716 399498
rect 92664 399434 92716 399440
rect 91744 398132 91796 398138
rect 91744 398074 91796 398080
rect 91100 393508 91152 393514
rect 91100 393450 91152 393456
rect 91008 388476 91060 388482
rect 91008 388418 91060 388424
rect 90364 387184 90416 387190
rect 90364 387126 90416 387132
rect 91020 385914 91048 388418
rect 88352 385886 88734 385914
rect 90022 385886 90312 385914
rect 90666 385886 91048 385914
rect 91112 385914 91140 393450
rect 91112 385886 91310 385914
rect 74644 385370 74672 385886
rect 92676 385778 92704 399434
rect 93780 396914 93808 436018
rect 94516 401033 94544 438806
rect 94976 437374 95004 440014
rect 95148 439612 95200 439618
rect 95148 439554 95200 439560
rect 95160 438870 95188 439554
rect 96448 438870 96476 440028
rect 97092 440014 97488 440028
rect 97736 440014 97948 440028
rect 96528 439544 96580 439550
rect 96528 439486 96580 439492
rect 95148 438864 95200 438870
rect 95148 438806 95200 438812
rect 96436 438864 96488 438870
rect 96436 438806 96488 438812
rect 95240 438796 95292 438802
rect 95240 438738 95292 438744
rect 94964 437368 95016 437374
rect 94964 437310 95016 437316
rect 94976 431954 95004 437310
rect 94976 431926 95188 431954
rect 94502 401024 94558 401033
rect 94502 400959 94558 400968
rect 93768 396908 93820 396914
rect 93768 396850 93820 396856
rect 94136 396772 94188 396778
rect 94136 396714 94188 396720
rect 93860 394120 93912 394126
rect 93860 394062 93912 394068
rect 92940 388000 92992 388006
rect 92940 387942 92992 387948
rect 92952 385914 92980 387942
rect 93872 386084 93900 394062
rect 93872 386056 93992 386084
rect 93964 385914 93992 386056
rect 92952 385886 93242 385914
rect 93886 385886 93992 385914
rect 94148 385914 94176 396714
rect 95160 395418 95188 431926
rect 95148 395412 95200 395418
rect 95148 395354 95200 395360
rect 95252 387122 95280 438738
rect 96448 431954 96476 438806
rect 96540 438802 96568 439486
rect 96620 438932 96672 438938
rect 96620 438874 96672 438880
rect 96528 438796 96580 438802
rect 96528 438738 96580 438744
rect 96448 431926 96568 431954
rect 96540 392698 96568 431926
rect 96632 400926 96660 438874
rect 97092 437889 97120 440014
rect 97264 439952 97316 439958
rect 97264 439894 97316 439900
rect 97078 437880 97134 437889
rect 97078 437815 97134 437824
rect 96620 400920 96672 400926
rect 96620 400862 96672 400868
rect 97276 398206 97304 439894
rect 97736 438938 97764 440014
rect 97724 438932 97776 438938
rect 97724 438874 97776 438880
rect 98380 438054 98408 440028
rect 99024 438870 99052 440028
rect 99012 438864 99064 438870
rect 99012 438806 99064 438812
rect 99392 438598 99420 443663
rect 99484 440298 99512 460906
rect 99930 442504 99986 442513
rect 99930 442439 99986 442448
rect 99944 440706 99972 442439
rect 99932 440700 99984 440706
rect 99932 440642 99984 440648
rect 99472 440292 99524 440298
rect 99472 440234 99524 440240
rect 99668 438977 99696 440028
rect 99654 438968 99710 438977
rect 99654 438903 99710 438912
rect 99380 438592 99432 438598
rect 99380 438534 99432 438540
rect 98368 438048 98420 438054
rect 98368 437990 98420 437996
rect 99288 438048 99340 438054
rect 99288 437990 99340 437996
rect 97264 398200 97316 398206
rect 97264 398142 97316 398148
rect 98000 395344 98052 395350
rect 98000 395286 98052 395292
rect 96712 394052 96764 394058
rect 96712 393994 96764 394000
rect 96528 392692 96580 392698
rect 96528 392634 96580 392640
rect 96528 391264 96580 391270
rect 96528 391206 96580 391212
rect 96158 389872 96214 389881
rect 96158 389807 96214 389816
rect 95240 387116 95292 387122
rect 95240 387058 95292 387064
rect 96172 385914 96200 389807
rect 96540 385914 96568 391206
rect 94148 385886 94530 385914
rect 95818 385886 96200 385914
rect 96462 385886 96568 385914
rect 96724 385914 96752 393994
rect 98012 385914 98040 395286
rect 99300 391338 99328 437990
rect 99288 391332 99340 391338
rect 99288 391274 99340 391280
rect 99380 389836 99432 389842
rect 99380 389778 99432 389784
rect 99392 388618 99420 389778
rect 99380 388612 99432 388618
rect 99380 388554 99432 388560
rect 100036 387938 100064 490758
rect 100312 473346 100340 540138
rect 100956 537985 100984 540138
rect 102227 540110 102272 540138
rect 100942 537976 100998 537985
rect 100942 537911 100998 537920
rect 102244 537606 102272 540110
rect 102232 537600 102284 537606
rect 102232 537542 102284 537548
rect 102888 537538 102916 540138
rect 103532 538218 103560 540138
rect 103520 538212 103572 538218
rect 103520 538154 103572 538160
rect 102876 537532 102928 537538
rect 102876 537474 102928 537480
rect 102048 536852 102100 536858
rect 102048 536794 102100 536800
rect 100668 491632 100720 491638
rect 100668 491574 100720 491580
rect 100680 491230 100708 491574
rect 101404 491292 101456 491298
rect 101404 491234 101456 491240
rect 100668 491224 100720 491230
rect 100668 491166 100720 491172
rect 100300 473340 100352 473346
rect 100300 473282 100352 473288
rect 100116 450560 100168 450566
rect 100116 450502 100168 450508
rect 100128 440230 100156 450502
rect 100116 440224 100168 440230
rect 100116 440166 100168 440172
rect 100680 398818 100708 491166
rect 100760 473340 100812 473346
rect 100760 473282 100812 473288
rect 100772 441153 100800 473282
rect 101034 446584 101090 446593
rect 101034 446519 101090 446528
rect 101048 445806 101076 446519
rect 101036 445800 101088 445806
rect 101036 445742 101088 445748
rect 100758 441144 100814 441153
rect 100758 441079 100814 441088
rect 100772 440366 100800 441079
rect 100760 440360 100812 440366
rect 100760 440302 100812 440308
rect 100852 440292 100904 440298
rect 100852 440234 100904 440240
rect 100864 440201 100892 440234
rect 100850 440192 100906 440201
rect 100850 440127 100906 440136
rect 100760 430636 100812 430642
rect 100760 430578 100812 430584
rect 100772 429894 100800 430578
rect 100760 429888 100812 429894
rect 100760 429830 100812 429836
rect 100668 398812 100720 398818
rect 100668 398754 100720 398760
rect 101416 393314 101444 491234
rect 101956 480956 102008 480962
rect 101956 480898 102008 480904
rect 101968 480185 101996 480898
rect 101954 480176 102010 480185
rect 101954 480111 102010 480120
rect 101956 451240 102008 451246
rect 101954 451208 101956 451217
rect 102008 451208 102010 451217
rect 101954 451143 102010 451152
rect 101968 430642 101996 451143
rect 102060 445806 102088 536794
rect 104176 528554 104204 540138
rect 104716 537736 104768 537742
rect 104716 537678 104768 537684
rect 104728 536178 104756 537678
rect 104716 536172 104768 536178
rect 104716 536114 104768 536120
rect 103716 528526 104204 528554
rect 102140 494012 102192 494018
rect 102140 493954 102192 493960
rect 102152 460934 102180 493954
rect 103426 488744 103482 488753
rect 103426 488679 103482 488688
rect 103440 488646 103468 488679
rect 103428 488640 103480 488646
rect 102874 488608 102930 488617
rect 103428 488582 103480 488588
rect 102874 488543 102930 488552
rect 102888 488442 102916 488543
rect 103336 488504 103388 488510
rect 103336 488446 103388 488452
rect 102876 488436 102928 488442
rect 102876 488378 102928 488384
rect 103348 488073 103376 488446
rect 103334 488064 103390 488073
rect 103334 487999 103390 488008
rect 103610 487248 103666 487257
rect 103610 487183 103666 487192
rect 103336 487144 103388 487150
rect 103336 487086 103388 487092
rect 103348 486577 103376 487086
rect 103334 486568 103390 486577
rect 103334 486503 103390 486512
rect 103428 486056 103480 486062
rect 103426 486024 103428 486033
rect 103480 486024 103482 486033
rect 103426 485959 103482 485968
rect 102232 485784 102284 485790
rect 102232 485726 102284 485732
rect 102244 485353 102272 485726
rect 102230 485344 102286 485353
rect 102230 485279 102286 485288
rect 102230 484664 102286 484673
rect 102230 484599 102286 484608
rect 102244 484430 102272 484599
rect 102232 484424 102284 484430
rect 102232 484366 102284 484372
rect 102230 483848 102286 483857
rect 102230 483783 102286 483792
rect 102244 483682 102272 483783
rect 102232 483676 102284 483682
rect 102232 483618 102284 483624
rect 102324 482996 102376 483002
rect 102324 482938 102376 482944
rect 102232 482656 102284 482662
rect 102336 482633 102364 482938
rect 102232 482598 102284 482604
rect 102322 482624 102378 482633
rect 102244 482497 102272 482598
rect 102322 482559 102378 482568
rect 102230 482488 102286 482497
rect 102230 482423 102286 482432
rect 102232 481636 102284 481642
rect 102232 481578 102284 481584
rect 102244 481545 102272 481578
rect 102324 481568 102376 481574
rect 102230 481536 102286 481545
rect 102324 481510 102376 481516
rect 102230 481471 102286 481480
rect 102336 481273 102364 481510
rect 102322 481264 102378 481273
rect 102322 481199 102378 481208
rect 102232 480208 102284 480214
rect 102232 480150 102284 480156
rect 102244 479913 102272 480150
rect 102230 479904 102286 479913
rect 102230 479839 102286 479848
rect 102874 477728 102930 477737
rect 102874 477663 102930 477672
rect 102888 477562 102916 477663
rect 102876 477556 102928 477562
rect 102876 477498 102928 477504
rect 102324 477488 102376 477494
rect 102324 477430 102376 477436
rect 102232 477420 102284 477426
rect 102232 477362 102284 477368
rect 102244 477057 102272 477362
rect 102230 477048 102286 477057
rect 102230 476983 102286 476992
rect 102336 476513 102364 477430
rect 102414 477184 102470 477193
rect 102414 477119 102470 477128
rect 102322 476504 102378 476513
rect 102322 476439 102378 476448
rect 102428 476066 102456 477119
rect 102416 476060 102468 476066
rect 102416 476002 102468 476008
rect 103336 476060 103388 476066
rect 103336 476002 103388 476008
rect 102232 475992 102284 475998
rect 102232 475934 102284 475940
rect 102244 475697 102272 475934
rect 102324 475924 102376 475930
rect 102324 475866 102376 475872
rect 102230 475688 102286 475697
rect 102230 475623 102286 475632
rect 102336 475153 102364 475866
rect 102322 475144 102378 475153
rect 102322 475079 102378 475088
rect 102232 474700 102284 474706
rect 102232 474642 102284 474648
rect 102244 474337 102272 474642
rect 102230 474328 102286 474337
rect 102230 474263 102286 474272
rect 102230 472968 102286 472977
rect 102230 472903 102286 472912
rect 102244 472666 102272 472903
rect 102324 472728 102376 472734
rect 102324 472670 102376 472676
rect 102232 472660 102284 472666
rect 102232 472602 102284 472608
rect 102336 472433 102364 472670
rect 102322 472424 102378 472433
rect 102322 472359 102378 472368
rect 102232 471980 102284 471986
rect 102232 471922 102284 471928
rect 102244 471617 102272 471922
rect 102230 471608 102286 471617
rect 102230 471543 102286 471552
rect 102784 471368 102836 471374
rect 102784 471310 102836 471316
rect 102796 470257 102824 471310
rect 103348 470594 103376 476002
rect 103426 474056 103482 474065
rect 103426 473991 103482 474000
rect 103440 472734 103468 473991
rect 103428 472728 103480 472734
rect 103428 472670 103480 472676
rect 103348 470566 103468 470594
rect 102782 470248 102838 470257
rect 102782 470183 102838 470192
rect 102232 469872 102284 469878
rect 102232 469814 102284 469820
rect 102244 469577 102272 469814
rect 102230 469568 102286 469577
rect 102230 469503 102286 469512
rect 102230 466848 102286 466857
rect 102230 466783 102286 466792
rect 102244 466478 102272 466783
rect 102232 466472 102284 466478
rect 102232 466414 102284 466420
rect 102230 466168 102286 466177
rect 102230 466103 102286 466112
rect 102244 465798 102272 466103
rect 102324 465860 102376 465866
rect 102324 465802 102376 465808
rect 102232 465792 102284 465798
rect 102232 465734 102284 465740
rect 102336 465497 102364 465802
rect 102322 465488 102378 465497
rect 102322 465423 102378 465432
rect 102232 463004 102284 463010
rect 102232 462946 102284 462952
rect 102244 462913 102272 462946
rect 102230 462904 102286 462913
rect 102230 462839 102286 462848
rect 102324 462324 102376 462330
rect 102324 462266 102376 462272
rect 102232 462256 102284 462262
rect 102232 462198 102284 462204
rect 102244 462097 102272 462198
rect 102230 462088 102286 462097
rect 102230 462023 102286 462032
rect 102336 461553 102364 462266
rect 102322 461544 102378 461553
rect 102322 461479 102378 461488
rect 102152 460906 102272 460934
rect 102138 460728 102194 460737
rect 102138 460663 102194 460672
rect 102152 460358 102180 460663
rect 102140 460352 102192 460358
rect 102140 460294 102192 460300
rect 102140 459536 102192 459542
rect 102140 459478 102192 459484
rect 102152 459377 102180 459478
rect 102138 459368 102194 459377
rect 102138 459303 102194 459312
rect 102138 458688 102194 458697
rect 102138 458623 102194 458632
rect 102152 458250 102180 458623
rect 102140 458244 102192 458250
rect 102140 458186 102192 458192
rect 102140 456748 102192 456754
rect 102140 456690 102192 456696
rect 102152 456657 102180 456690
rect 102138 456648 102194 456657
rect 102138 456583 102194 456592
rect 102138 454744 102194 454753
rect 102138 454679 102140 454688
rect 102192 454679 102194 454688
rect 102140 454650 102192 454656
rect 102140 454028 102192 454034
rect 102140 453970 102192 453976
rect 102152 453937 102180 453970
rect 102138 453928 102194 453937
rect 102138 453863 102194 453872
rect 102138 452024 102194 452033
rect 102138 451959 102140 451968
rect 102192 451959 102194 451968
rect 102140 451930 102192 451936
rect 102138 449848 102194 449857
rect 102138 449783 102140 449792
rect 102192 449783 102194 449792
rect 102140 449754 102192 449760
rect 102140 447976 102192 447982
rect 102140 447918 102192 447924
rect 102152 447817 102180 447918
rect 102138 447808 102194 447817
rect 102138 447743 102194 447752
rect 102048 445800 102100 445806
rect 102048 445742 102100 445748
rect 102140 445732 102192 445738
rect 102140 445674 102192 445680
rect 102152 445233 102180 445674
rect 102138 445224 102194 445233
rect 102138 445159 102194 445168
rect 102140 445052 102192 445058
rect 102140 444994 102192 445000
rect 102152 443737 102180 444994
rect 102138 443728 102194 443737
rect 102138 443663 102194 443672
rect 102138 442368 102194 442377
rect 102138 442303 102194 442312
rect 102152 441658 102180 442303
rect 102140 441652 102192 441658
rect 102140 441594 102192 441600
rect 102244 438054 102272 460906
rect 102324 460896 102376 460902
rect 102324 460838 102376 460844
rect 102336 460193 102364 460838
rect 102322 460184 102378 460193
rect 102322 460119 102378 460128
rect 102324 458176 102376 458182
rect 102324 458118 102376 458124
rect 102336 458017 102364 458118
rect 102322 458008 102378 458017
rect 102322 457943 102378 457952
rect 102876 455388 102928 455394
rect 102876 455330 102928 455336
rect 102888 454617 102916 455330
rect 102874 454608 102930 454617
rect 102874 454543 102930 454552
rect 103334 454608 103390 454617
rect 103334 454543 103390 454552
rect 102324 453960 102376 453966
rect 102324 453902 102376 453908
rect 102336 453393 102364 453902
rect 102322 453384 102378 453393
rect 102322 453319 102378 453328
rect 102508 451920 102560 451926
rect 102508 451862 102560 451868
rect 102520 450673 102548 451862
rect 102506 450664 102562 450673
rect 102506 450599 102562 450608
rect 102324 449880 102376 449886
rect 102324 449822 102376 449828
rect 102336 449313 102364 449822
rect 102322 449304 102378 449313
rect 102322 449239 102378 449248
rect 102322 447944 102378 447953
rect 102322 447879 102378 447888
rect 102336 447846 102364 447879
rect 102324 447840 102376 447846
rect 102324 447782 102376 447788
rect 102322 445768 102378 445777
rect 102322 445703 102378 445712
rect 102336 445330 102364 445703
rect 102324 445324 102376 445330
rect 102324 445266 102376 445272
rect 102324 444032 102376 444038
rect 102324 443974 102376 443980
rect 102336 443873 102364 443974
rect 102322 443864 102378 443873
rect 102322 443799 102378 443808
rect 102232 438048 102284 438054
rect 102232 437990 102284 437996
rect 101956 430636 102008 430642
rect 101956 430578 102008 430584
rect 101324 393286 101444 393314
rect 101324 389366 101352 393286
rect 103348 391241 103376 454543
rect 103334 391232 103390 391241
rect 103334 391167 103390 391176
rect 103440 390017 103468 470566
rect 103520 469940 103572 469946
rect 103520 469882 103572 469888
rect 103532 469033 103560 469882
rect 103518 469024 103574 469033
rect 103518 468959 103574 468968
rect 103520 465724 103572 465730
rect 103520 465666 103572 465672
rect 103532 464953 103560 465666
rect 103518 464944 103574 464953
rect 103518 464879 103574 464888
rect 103520 457496 103572 457502
rect 103520 457438 103572 457444
rect 103532 456113 103560 457438
rect 103518 456104 103574 456113
rect 103518 456039 103574 456048
rect 103624 440162 103652 487183
rect 103716 445738 103744 528526
rect 104716 483064 104768 483070
rect 104716 483006 104768 483012
rect 104728 482662 104756 483006
rect 104716 482656 104768 482662
rect 104716 482598 104768 482604
rect 104716 464160 104768 464166
rect 104714 464128 104716 464137
rect 104768 464128 104770 464137
rect 104714 464063 104770 464072
rect 104716 447908 104768 447914
rect 104716 447850 104768 447856
rect 103704 445732 103756 445738
rect 103704 445674 103756 445680
rect 104164 445732 104216 445738
rect 104164 445674 104216 445680
rect 103612 440156 103664 440162
rect 103612 440098 103664 440104
rect 104176 403646 104204 445674
rect 104256 430636 104308 430642
rect 104256 430578 104308 430584
rect 104164 403640 104216 403646
rect 104164 403582 104216 403588
rect 104164 398812 104216 398818
rect 104164 398754 104216 398760
rect 103796 395480 103848 395486
rect 103796 395422 103848 395428
rect 103520 394732 103572 394738
rect 103520 394674 103572 394680
rect 103426 390008 103482 390017
rect 103426 389943 103482 389952
rect 101312 389360 101364 389366
rect 101312 389302 101364 389308
rect 100024 387932 100076 387938
rect 100024 387874 100076 387880
rect 99288 387116 99340 387122
rect 99288 387058 99340 387064
rect 99300 385914 99328 387058
rect 100036 385914 100064 387874
rect 101324 385914 101352 389302
rect 101402 388920 101458 388929
rect 101402 388855 101458 388864
rect 101416 388006 101444 388855
rect 103532 388550 103560 394674
rect 103520 388544 103572 388550
rect 103520 388486 103572 388492
rect 102600 388408 102652 388414
rect 102600 388350 102652 388356
rect 101404 388000 101456 388006
rect 101404 387942 101456 387948
rect 96724 385886 97106 385914
rect 98012 385886 98394 385914
rect 99038 385886 99328 385914
rect 99682 385886 100064 385914
rect 100970 385886 101352 385914
rect 92598 385750 92704 385778
rect 101416 385778 101444 387942
rect 102612 385914 102640 388350
rect 103704 386504 103756 386510
rect 103704 386446 103756 386452
rect 103716 385914 103744 386446
rect 102258 385886 102640 385914
rect 103546 385886 103744 385914
rect 103808 385914 103836 395422
rect 104176 386510 104204 398754
rect 104268 398274 104296 430578
rect 104256 398268 104308 398274
rect 104256 398210 104308 398216
rect 104728 394738 104756 447850
rect 104820 446026 104848 540138
rect 105478 540110 105584 540138
rect 105556 536858 105584 540110
rect 105544 536852 105596 536858
rect 105544 536794 105596 536800
rect 104898 481536 104954 481545
rect 104898 481471 104954 481480
rect 104912 480321 104940 481471
rect 104898 480312 104954 480321
rect 104898 480247 104954 480256
rect 104912 480214 104940 480247
rect 104900 480208 104952 480214
rect 104900 480150 104952 480156
rect 105544 477624 105596 477630
rect 105544 477566 105596 477572
rect 105556 460358 105584 477566
rect 105636 466540 105688 466546
rect 105636 466482 105688 466488
rect 105544 460352 105596 460358
rect 105544 460294 105596 460300
rect 105358 450528 105414 450537
rect 105358 450463 105414 450472
rect 105372 449818 105400 450463
rect 105360 449812 105412 449818
rect 105360 449754 105412 449760
rect 104820 445998 104940 446026
rect 104912 445330 104940 445998
rect 104900 445324 104952 445330
rect 104900 445266 104952 445272
rect 104808 445120 104860 445126
rect 104808 445062 104860 445068
rect 104820 444038 104848 445062
rect 104808 444032 104860 444038
rect 104808 443974 104860 443980
rect 104716 394732 104768 394738
rect 104716 394674 104768 394680
rect 105556 392834 105584 460294
rect 105648 455394 105676 466482
rect 105636 455388 105688 455394
rect 105636 455330 105688 455336
rect 105740 451246 105768 543759
rect 105818 540424 105874 540433
rect 105818 540359 105874 540368
rect 105832 539578 105860 540359
rect 105820 539572 105872 539578
rect 105820 539514 105872 539520
rect 106200 481710 106228 572727
rect 106292 560425 106320 698906
rect 108960 586514 108988 702510
rect 108776 586486 108988 586514
rect 106648 584112 106700 584118
rect 106648 584054 106700 584060
rect 106922 584080 106978 584089
rect 106660 580990 106688 584054
rect 106922 584015 106978 584024
rect 106648 580984 106700 580990
rect 106648 580926 106700 580932
rect 106370 574696 106426 574705
rect 106370 574631 106426 574640
rect 106278 560416 106334 560425
rect 106278 560351 106334 560360
rect 106280 490680 106332 490686
rect 106280 490622 106332 490628
rect 106292 489870 106320 490622
rect 106280 489864 106332 489870
rect 106280 489806 106332 489812
rect 106280 487824 106332 487830
rect 106280 487766 106332 487772
rect 106292 486062 106320 487766
rect 106280 486056 106332 486062
rect 106280 485998 106332 486004
rect 106384 483002 106412 574631
rect 106936 566506 106964 584015
rect 107660 582480 107712 582486
rect 107660 582422 107712 582428
rect 107672 573345 107700 582422
rect 108672 581800 108724 581806
rect 108672 581742 108724 581748
rect 108684 581126 108712 581742
rect 108672 581120 108724 581126
rect 108672 581062 108724 581068
rect 108394 579456 108450 579465
rect 108394 579391 108450 579400
rect 108408 578338 108436 579391
rect 108396 578332 108448 578338
rect 108396 578274 108448 578280
rect 108776 577538 108804 586486
rect 109130 581768 109186 581777
rect 109130 581703 109186 581712
rect 108946 580816 109002 580825
rect 108946 580751 109002 580760
rect 108854 580136 108910 580145
rect 108854 580071 108910 580080
rect 108868 579578 108896 580071
rect 108960 579766 108988 580751
rect 108948 579760 109000 579766
rect 108948 579702 109000 579708
rect 108868 579550 109080 579578
rect 108946 578776 109002 578785
rect 108946 578711 109002 578720
rect 108960 578270 108988 578711
rect 108948 578264 109000 578270
rect 108948 578206 109000 578212
rect 108946 578096 109002 578105
rect 108946 578031 109002 578040
rect 108854 577552 108910 577561
rect 108776 577510 108854 577538
rect 108854 577487 108856 577496
rect 108908 577487 108910 577496
rect 108856 577458 108908 577464
rect 108960 576910 108988 578031
rect 108948 576904 109000 576910
rect 108948 576846 109000 576852
rect 108486 576736 108542 576745
rect 108486 576671 108542 576680
rect 108500 575550 108528 576671
rect 108946 576192 109002 576201
rect 108946 576127 108948 576136
rect 109000 576127 109002 576136
rect 108948 576098 109000 576104
rect 108488 575544 108540 575550
rect 108488 575486 108540 575492
rect 108946 574016 109002 574025
rect 108946 573951 109002 573960
rect 108960 573374 108988 573951
rect 108948 573368 109000 573374
rect 107658 573336 107714 573345
rect 108948 573310 109000 573316
rect 107658 573271 107714 573280
rect 107672 572762 107700 573271
rect 107660 572756 107712 572762
rect 107660 572698 107712 572704
rect 108946 571976 109002 571985
rect 108946 571911 109002 571920
rect 107842 571432 107898 571441
rect 108960 571402 108988 571911
rect 107842 571367 107898 571376
rect 108948 571396 109000 571402
rect 106924 566500 106976 566506
rect 106924 566442 106976 566448
rect 107750 557696 107806 557705
rect 107750 557631 107806 557640
rect 107658 556336 107714 556345
rect 107658 556271 107714 556280
rect 107014 551576 107070 551585
rect 107014 551511 107070 551520
rect 106922 542056 106978 542065
rect 106922 541991 106978 542000
rect 106372 482996 106424 483002
rect 106372 482938 106424 482944
rect 106188 481704 106240 481710
rect 106188 481646 106240 481652
rect 106200 481506 106228 481646
rect 106188 481500 106240 481506
rect 106188 481442 106240 481448
rect 106646 462224 106702 462233
rect 106646 462159 106702 462168
rect 106660 461009 106688 462159
rect 106646 461000 106702 461009
rect 106646 460935 106702 460944
rect 106660 460902 106688 460935
rect 106648 460896 106700 460902
rect 106648 460838 106700 460844
rect 106188 454844 106240 454850
rect 106188 454786 106240 454792
rect 105728 451240 105780 451246
rect 105728 451182 105780 451188
rect 105726 447264 105782 447273
rect 105726 447199 105782 447208
rect 105636 445324 105688 445330
rect 105636 445266 105688 445272
rect 105544 392828 105596 392834
rect 105544 392770 105596 392776
rect 104532 390108 104584 390114
rect 104532 390050 104584 390056
rect 104164 386504 104216 386510
rect 104164 386446 104216 386452
rect 104544 385914 104572 390050
rect 103808 385886 104190 385914
rect 104544 385886 104834 385914
rect 101416 385750 101614 385778
rect 105648 385762 105676 445266
rect 105740 438666 105768 447199
rect 105728 438660 105780 438666
rect 105728 438602 105780 438608
rect 106200 388521 106228 454786
rect 106936 449954 106964 541991
rect 107028 528630 107056 551511
rect 107016 528624 107068 528630
rect 107016 528566 107068 528572
rect 107384 489864 107436 489870
rect 107384 489806 107436 489812
rect 107016 459604 107068 459610
rect 107016 459546 107068 459552
rect 106924 449948 106976 449954
rect 106924 449890 106976 449896
rect 107028 447982 107056 459546
rect 107016 447976 107068 447982
rect 107016 447918 107068 447924
rect 107028 431954 107056 447918
rect 106936 431926 107056 431954
rect 106936 395321 106964 431926
rect 107396 402974 107424 489806
rect 107568 482996 107620 483002
rect 107568 482938 107620 482944
rect 107580 481778 107608 482938
rect 107568 481772 107620 481778
rect 107568 481714 107620 481720
rect 107672 464166 107700 556271
rect 107764 465866 107792 557631
rect 107856 552673 107884 571367
rect 108948 571338 109000 571344
rect 108854 570616 108910 570625
rect 108854 570551 108910 570560
rect 108868 570042 108896 570551
rect 108946 570072 109002 570081
rect 108856 570036 108908 570042
rect 108946 570007 109002 570016
rect 108856 569978 108908 569984
rect 108960 569974 108988 570007
rect 108948 569968 109000 569974
rect 108948 569910 109000 569916
rect 108946 569256 109002 569265
rect 108946 569191 109002 569200
rect 108960 568614 108988 569191
rect 108948 568608 109000 568614
rect 108948 568550 109000 568556
rect 108946 567896 109002 567905
rect 108946 567831 109002 567840
rect 108960 567594 108988 567831
rect 108948 567588 109000 567594
rect 108948 567530 109000 567536
rect 108948 567248 109000 567254
rect 108946 567216 108948 567225
rect 109000 567216 109002 567225
rect 108946 567151 109002 567160
rect 108394 566536 108450 566545
rect 108394 566471 108450 566480
rect 108408 565962 108436 566471
rect 108396 565956 108448 565962
rect 108396 565898 108448 565904
rect 108948 565888 109000 565894
rect 108946 565856 108948 565865
rect 109000 565856 109002 565865
rect 108946 565791 109002 565800
rect 108946 565176 109002 565185
rect 108946 565111 109002 565120
rect 108960 564466 108988 565111
rect 108948 564460 109000 564466
rect 108948 564402 109000 564408
rect 108396 564392 108448 564398
rect 108396 564334 108448 564340
rect 108408 563961 108436 564334
rect 108394 563952 108450 563961
rect 108394 563887 108450 563896
rect 108946 562456 109002 562465
rect 108946 562391 109002 562400
rect 108960 561746 108988 562391
rect 108948 561740 109000 561746
rect 108948 561682 109000 561688
rect 108946 561096 109002 561105
rect 108946 561031 109002 561040
rect 108210 560416 108266 560425
rect 108210 560351 108212 560360
rect 108264 560351 108266 560360
rect 108212 560322 108264 560328
rect 108960 560318 108988 561031
rect 108948 560312 109000 560318
rect 108948 560254 109000 560260
rect 108854 559736 108910 559745
rect 108854 559671 108910 559680
rect 108868 558958 108896 559671
rect 108946 559056 109002 559065
rect 108946 558991 108948 559000
rect 109000 558991 109002 559000
rect 108948 558962 109000 558968
rect 108856 558952 108908 558958
rect 108856 558894 108908 558900
rect 108946 558376 109002 558385
rect 108946 558311 109002 558320
rect 108960 557598 108988 558311
rect 108948 557592 109000 557598
rect 108948 557534 109000 557540
rect 108946 557016 109002 557025
rect 108946 556951 109002 556960
rect 108960 556238 108988 556951
rect 108948 556232 109000 556238
rect 108948 556174 109000 556180
rect 108856 556164 108908 556170
rect 108856 556106 108908 556112
rect 108868 555801 108896 556106
rect 108854 555792 108910 555801
rect 108854 555727 108910 555736
rect 108946 554296 109002 554305
rect 108946 554231 109002 554240
rect 108960 553450 108988 554231
rect 108948 553444 109000 553450
rect 108948 553386 109000 553392
rect 108118 552936 108174 552945
rect 108118 552871 108174 552880
rect 107842 552664 107898 552673
rect 107842 552599 107898 552608
rect 107934 546816 107990 546825
rect 107934 546751 107990 546760
rect 107842 540696 107898 540705
rect 107842 540631 107898 540640
rect 107856 539646 107884 540631
rect 107844 539640 107896 539646
rect 107844 539582 107896 539588
rect 107948 539458 107976 546751
rect 107856 539430 107976 539458
rect 107856 466546 107884 539430
rect 108132 539322 108160 552871
rect 108946 550896 109002 550905
rect 108946 550831 109002 550840
rect 108960 550662 108988 550831
rect 108948 550656 109000 550662
rect 108948 550598 109000 550604
rect 108854 550216 108910 550225
rect 108854 550151 108910 550160
rect 108868 549370 108896 550151
rect 108946 549536 109002 549545
rect 108946 549471 109002 549480
rect 108856 549364 108908 549370
rect 108856 549306 108908 549312
rect 108960 549302 108988 549471
rect 108948 549296 109000 549302
rect 108948 549238 109000 549244
rect 108946 548856 109002 548865
rect 108946 548791 109002 548800
rect 108960 547942 108988 548791
rect 108948 547936 109000 547942
rect 108948 547878 109000 547884
rect 108946 547496 109002 547505
rect 108946 547431 109002 547440
rect 108960 546514 108988 547431
rect 108948 546508 109000 546514
rect 108948 546450 109000 546456
rect 108946 546136 109002 546145
rect 108946 546071 109002 546080
rect 108960 545766 108988 546071
rect 108948 545760 109000 545766
rect 108948 545702 109000 545708
rect 108946 545456 109002 545465
rect 108946 545391 109002 545400
rect 108960 545154 108988 545391
rect 108948 545148 109000 545154
rect 108948 545090 109000 545096
rect 108946 543416 109002 543425
rect 108946 543351 109002 543360
rect 108960 542434 108988 543351
rect 108948 542428 109000 542434
rect 108948 542370 109000 542376
rect 108946 540016 109002 540025
rect 108946 539951 109002 539960
rect 108960 539714 108988 539951
rect 108948 539708 109000 539714
rect 108948 539650 109000 539656
rect 107948 539294 108160 539322
rect 107948 477630 107976 539294
rect 109052 488442 109080 579550
rect 109144 538966 109172 581703
rect 109684 541000 109736 541006
rect 109684 540942 109736 540948
rect 109132 538960 109184 538966
rect 109132 538902 109184 538908
rect 109696 538218 109724 540942
rect 110340 539714 110368 703054
rect 111708 702908 111760 702914
rect 111708 702850 111760 702856
rect 110512 583908 110564 583914
rect 110512 583850 110564 583856
rect 110420 572756 110472 572762
rect 110420 572698 110472 572704
rect 110328 539708 110380 539714
rect 110328 539650 110380 539656
rect 109684 538212 109736 538218
rect 109684 538154 109736 538160
rect 109132 536172 109184 536178
rect 109132 536114 109184 536120
rect 109040 488436 109092 488442
rect 109040 488378 109092 488384
rect 109052 487898 109080 488378
rect 109040 487892 109092 487898
rect 109040 487834 109092 487840
rect 107936 477624 107988 477630
rect 107936 477566 107988 477572
rect 109040 472728 109092 472734
rect 109040 472670 109092 472676
rect 108302 471880 108358 471889
rect 108302 471815 108358 471824
rect 108316 471073 108344 471815
rect 109052 471306 109080 472670
rect 109040 471300 109092 471306
rect 109040 471242 109092 471248
rect 108302 471064 108358 471073
rect 108302 470999 108358 471008
rect 107844 466540 107896 466546
rect 107844 466482 107896 466488
rect 107752 465860 107804 465866
rect 107752 465802 107804 465808
rect 107660 464160 107712 464166
rect 107660 464102 107712 464108
rect 107568 462392 107620 462398
rect 107568 462334 107620 462340
rect 107580 462262 107608 462334
rect 107568 462256 107620 462262
rect 107568 462198 107620 462204
rect 108212 458856 108264 458862
rect 108212 458798 108264 458804
rect 108224 458182 108252 458798
rect 108212 458176 108264 458182
rect 108212 458118 108264 458124
rect 108212 454776 108264 454782
rect 108212 454718 108264 454724
rect 108224 453966 108252 454718
rect 108212 453960 108264 453966
rect 108212 453902 108264 453908
rect 107396 402946 107516 402974
rect 106922 395312 106978 395321
rect 106922 395247 106978 395256
rect 107016 388544 107068 388550
rect 106186 388512 106242 388521
rect 107016 388486 107068 388492
rect 106186 388447 106242 388456
rect 106200 388414 106228 388447
rect 106188 388408 106240 388414
rect 106188 388350 106240 388356
rect 106188 387864 106240 387870
rect 106188 387806 106240 387812
rect 106200 385914 106228 387806
rect 107028 385914 107056 388486
rect 107488 385914 107516 402946
rect 108316 387190 108344 470999
rect 108396 466608 108448 466614
rect 108396 466550 108448 466556
rect 108408 437306 108436 466550
rect 108486 465760 108542 465769
rect 108486 465695 108542 465704
rect 108396 437300 108448 437306
rect 108396 437242 108448 437248
rect 108500 437238 108528 465695
rect 109144 450566 109172 536114
rect 109776 491972 109828 491978
rect 109776 491914 109828 491920
rect 109684 490612 109736 490618
rect 109684 490554 109736 490560
rect 109132 450560 109184 450566
rect 109132 450502 109184 450508
rect 108488 437232 108540 437238
rect 108488 437174 108540 437180
rect 108762 388376 108818 388385
rect 108762 388311 108818 388320
rect 108776 387870 108804 388311
rect 109696 388074 109724 490554
rect 109788 394670 109816 491914
rect 110432 481642 110460 572698
rect 110524 493474 110552 583850
rect 110604 572892 110656 572898
rect 110604 572834 110656 572840
rect 110616 556170 110644 572834
rect 110604 556164 110656 556170
rect 110604 556106 110656 556112
rect 110616 555490 110644 556106
rect 110604 555484 110656 555490
rect 110604 555426 110656 555432
rect 111720 544513 111748 702850
rect 117228 702772 117280 702778
rect 117228 702714 117280 702720
rect 113088 702704 113140 702710
rect 113088 702646 113140 702652
rect 111798 583944 111854 583953
rect 111798 583879 111854 583888
rect 111706 544504 111762 544513
rect 111706 544439 111762 544448
rect 110604 500404 110656 500410
rect 110604 500346 110656 500352
rect 110512 493468 110564 493474
rect 110512 493410 110564 493416
rect 110512 491496 110564 491502
rect 110512 491438 110564 491444
rect 110524 491298 110552 491438
rect 110512 491292 110564 491298
rect 110512 491234 110564 491240
rect 110420 481636 110472 481642
rect 110420 481578 110472 481584
rect 110616 439618 110644 500346
rect 111812 494902 111840 583879
rect 111892 578332 111944 578338
rect 111892 578274 111944 578280
rect 111800 494896 111852 494902
rect 111800 494838 111852 494844
rect 111812 494737 111840 494838
rect 111798 494728 111854 494737
rect 111798 494663 111854 494672
rect 111064 492040 111116 492046
rect 111064 491982 111116 491988
rect 110604 439612 110656 439618
rect 110604 439554 110656 439560
rect 109776 394664 109828 394670
rect 109776 394606 109828 394612
rect 110880 394188 110932 394194
rect 110880 394130 110932 394136
rect 110892 393446 110920 394130
rect 110880 393440 110932 393446
rect 110880 393382 110932 393388
rect 110328 392760 110380 392766
rect 110328 392702 110380 392708
rect 109684 388068 109736 388074
rect 109684 388010 109736 388016
rect 108764 387864 108816 387870
rect 108764 387806 108816 387812
rect 108304 387184 108356 387190
rect 108304 387126 108356 387132
rect 109696 385914 109724 388010
rect 110340 385914 110368 392702
rect 106122 385886 106228 385914
rect 106766 385886 107056 385914
rect 107410 385886 107516 385914
rect 109342 385886 109724 385914
rect 109986 385886 110368 385914
rect 110892 385914 110920 393382
rect 111076 392086 111104 491982
rect 111708 491292 111760 491298
rect 111708 491234 111760 491240
rect 111156 481636 111208 481642
rect 111156 481578 111208 481584
rect 111168 480282 111196 481578
rect 111156 480276 111208 480282
rect 111156 480218 111208 480224
rect 111064 392080 111116 392086
rect 111064 392022 111116 392028
rect 111720 389638 111748 491234
rect 111800 489932 111852 489938
rect 111800 489874 111852 489880
rect 111812 389842 111840 489874
rect 111904 488510 111932 578274
rect 111984 565956 112036 565962
rect 111984 565898 112036 565904
rect 111892 488504 111944 488510
rect 111892 488446 111944 488452
rect 111904 487966 111932 488446
rect 111892 487960 111944 487966
rect 111892 487902 111944 487908
rect 111892 477556 111944 477562
rect 111892 477498 111944 477504
rect 111904 477358 111932 477498
rect 111892 477352 111944 477358
rect 111892 477294 111944 477300
rect 111996 477170 112024 565898
rect 113100 545766 113128 702646
rect 116124 588600 116176 588606
rect 116124 588542 116176 588548
rect 114560 585336 114612 585342
rect 114560 585278 114612 585284
rect 113364 583976 113416 583982
rect 113364 583918 113416 583924
rect 113272 581188 113324 581194
rect 113272 581130 113324 581136
rect 113088 545760 113140 545766
rect 113088 545702 113140 545708
rect 113284 534954 113312 581130
rect 113272 534948 113324 534954
rect 113272 534890 113324 534896
rect 113272 532092 113324 532098
rect 113272 532034 113324 532040
rect 112076 497616 112128 497622
rect 112076 497558 112128 497564
rect 111904 477142 112024 477170
rect 111904 475930 111932 477142
rect 111892 475924 111944 475930
rect 111892 475866 111944 475872
rect 111904 475386 111932 475866
rect 111892 475380 111944 475386
rect 111892 475322 111944 475328
rect 112088 436014 112116 497558
rect 113180 495032 113232 495038
rect 113180 494974 113232 494980
rect 113088 484356 113140 484362
rect 113088 484298 113140 484304
rect 113100 479505 113128 484298
rect 113086 479496 113142 479505
rect 113086 479431 113142 479440
rect 113088 477352 113140 477358
rect 113088 477294 113140 477300
rect 113100 474026 113128 477294
rect 113088 474020 113140 474026
rect 113088 473962 113140 473968
rect 113088 443692 113140 443698
rect 113088 443634 113140 443640
rect 112076 436008 112128 436014
rect 112076 435950 112128 435956
rect 111984 394664 112036 394670
rect 111984 394606 112036 394612
rect 111800 389836 111852 389842
rect 111800 389778 111852 389784
rect 111708 389632 111760 389638
rect 111708 389574 111760 389580
rect 111996 385914 112024 394606
rect 113100 388482 113128 443634
rect 113192 442513 113220 494974
rect 113284 466614 113312 532034
rect 113376 493474 113404 583918
rect 113824 567588 113876 567594
rect 113824 567530 113876 567536
rect 113364 493468 113416 493474
rect 113364 493410 113416 493416
rect 113364 480276 113416 480282
rect 113364 480218 113416 480224
rect 113272 466608 113324 466614
rect 113272 466550 113324 466556
rect 113178 442504 113234 442513
rect 113178 442439 113234 442448
rect 113088 388476 113140 388482
rect 113088 388418 113140 388424
rect 112810 387968 112866 387977
rect 112810 387903 112866 387912
rect 112824 385914 112852 387903
rect 110892 385886 111274 385914
rect 111918 385886 112208 385914
rect 112562 385886 112852 385914
rect 105636 385756 105688 385762
rect 105636 385698 105688 385704
rect 74814 385384 74870 385393
rect 74644 385342 74814 385370
rect 107488 385370 107516 385886
rect 112180 385422 112208 385886
rect 113376 385694 113404 480218
rect 113836 477562 113864 567530
rect 114572 491230 114600 585278
rect 114652 583772 114704 583778
rect 114652 583714 114704 583720
rect 114664 491434 114692 583714
rect 114836 580984 114888 580990
rect 114836 580926 114888 580932
rect 114744 539708 114796 539714
rect 114744 539650 114796 539656
rect 114652 491428 114704 491434
rect 114652 491370 114704 491376
rect 114560 491224 114612 491230
rect 114560 491166 114612 491172
rect 114376 488504 114428 488510
rect 114376 488446 114428 488452
rect 114388 487257 114416 488446
rect 114374 487248 114430 487257
rect 114374 487183 114430 487192
rect 113824 477556 113876 477562
rect 113824 477498 113876 477504
rect 114756 459610 114784 539650
rect 114848 536110 114876 580926
rect 115940 577516 115992 577522
rect 115940 577458 115992 577464
rect 114836 536104 114888 536110
rect 114836 536046 114888 536052
rect 114928 498228 114980 498234
rect 114928 498170 114980 498176
rect 114836 490612 114888 490618
rect 114836 490554 114888 490560
rect 114848 490006 114876 490554
rect 114836 490000 114888 490006
rect 114836 489942 114888 489948
rect 114744 459604 114796 459610
rect 114744 459546 114796 459552
rect 114848 454850 114876 489942
rect 114836 454844 114888 454850
rect 114836 454786 114888 454792
rect 114940 447914 114968 498170
rect 115480 491428 115532 491434
rect 115480 491370 115532 491376
rect 115492 491230 115520 491370
rect 115480 491224 115532 491230
rect 115480 491166 115532 491172
rect 115848 489184 115900 489190
rect 115848 489126 115900 489132
rect 115860 488646 115888 489126
rect 115848 488640 115900 488646
rect 115848 488582 115900 488588
rect 115860 483002 115888 488582
rect 115952 485790 115980 577458
rect 116032 557592 116084 557598
rect 116032 557534 116084 557540
rect 115940 485784 115992 485790
rect 115940 485726 115992 485732
rect 115848 482996 115900 483002
rect 115848 482938 115900 482944
rect 115296 481772 115348 481778
rect 115296 481714 115348 481720
rect 114928 447908 114980 447914
rect 114928 447850 114980 447856
rect 115308 402974 115336 481714
rect 116044 465798 116072 557534
rect 116136 536178 116164 588542
rect 116216 585268 116268 585274
rect 116216 585210 116268 585216
rect 116228 538898 116256 585210
rect 117240 564534 117268 702714
rect 130384 630692 130436 630698
rect 130384 630634 130436 630640
rect 124220 589348 124272 589354
rect 124220 589290 124272 589296
rect 121460 587172 121512 587178
rect 121460 587114 121512 587120
rect 120172 586628 120224 586634
rect 120172 586570 120224 586576
rect 118700 586560 118752 586566
rect 118700 586502 118752 586508
rect 117412 582684 117464 582690
rect 117412 582626 117464 582632
rect 117320 575544 117372 575550
rect 117320 575486 117372 575492
rect 117228 564528 117280 564534
rect 117228 564470 117280 564476
rect 117240 564398 117268 564470
rect 117228 564392 117280 564398
rect 117228 564334 117280 564340
rect 116216 538892 116268 538898
rect 116216 538834 116268 538840
rect 116124 536172 116176 536178
rect 116124 536114 116176 536120
rect 116124 500472 116176 500478
rect 116124 500414 116176 500420
rect 116032 465792 116084 465798
rect 116032 465734 116084 465740
rect 115848 458176 115900 458182
rect 115848 458118 115900 458124
rect 115308 402946 115428 402974
rect 113640 392080 113692 392086
rect 113640 392022 113692 392028
rect 113652 389230 113680 392022
rect 114836 389632 114888 389638
rect 114836 389574 114888 389580
rect 114282 389328 114338 389337
rect 114282 389263 114284 389272
rect 114336 389263 114338 389272
rect 114284 389234 114336 389240
rect 113640 389224 113692 389230
rect 113640 389166 113692 389172
rect 113652 385778 113680 389166
rect 114296 385778 114324 389234
rect 114848 385914 114876 389574
rect 115294 385928 115350 385937
rect 114848 385886 115294 385914
rect 115294 385863 115350 385872
rect 113652 385750 113850 385778
rect 114296 385750 114494 385778
rect 113364 385688 113416 385694
rect 113364 385630 113416 385636
rect 112168 385416 112220 385422
rect 107120 385354 107516 385370
rect 74814 385319 74870 385328
rect 107108 385348 107516 385354
rect 107160 385342 107516 385348
rect 108698 385354 108988 385370
rect 112168 385358 112220 385364
rect 108698 385348 109000 385354
rect 108698 385342 108948 385348
rect 107108 385290 107160 385296
rect 108948 385290 109000 385296
rect 115400 378593 115428 402946
rect 115572 389496 115624 389502
rect 115572 389438 115624 389444
rect 115584 385778 115612 389438
rect 115584 385750 115782 385778
rect 115386 378584 115442 378593
rect 115386 378519 115442 378528
rect 115294 377904 115350 377913
rect 115216 377862 115294 377890
rect 70308 376032 70360 376038
rect 70308 375974 70360 375980
rect 69756 370524 69808 370530
rect 69756 370466 69808 370472
rect 69664 367804 69716 367810
rect 69664 367746 69716 367752
rect 115216 364334 115244 377862
rect 115294 377839 115350 377848
rect 69308 364306 69704 364334
rect 115216 364306 115336 364334
rect 69202 352744 69258 352753
rect 69202 352679 69258 352688
rect 69216 329186 69244 352679
rect 69676 345014 69704 364306
rect 69676 344986 69796 345014
rect 69768 340082 69796 344986
rect 115308 344593 115336 364306
rect 115860 357406 115888 458118
rect 115938 452024 115994 452033
rect 115938 451959 115940 451968
rect 115992 451959 115994 451968
rect 115940 451930 115992 451936
rect 116136 440910 116164 500414
rect 116216 487960 116268 487966
rect 116216 487902 116268 487908
rect 116124 440904 116176 440910
rect 116124 440846 116176 440852
rect 116124 392488 116176 392494
rect 116124 392430 116176 392436
rect 116032 384396 116084 384402
rect 116032 384338 116084 384344
rect 116044 384033 116072 384338
rect 116030 384024 116086 384033
rect 116030 383959 116086 383968
rect 115938 370288 115994 370297
rect 115938 370223 115994 370232
rect 115952 369986 115980 370223
rect 115940 369980 115992 369986
rect 115940 369922 115992 369928
rect 115848 357400 115900 357406
rect 115848 357342 115900 357348
rect 115294 344584 115350 344593
rect 115294 344519 115350 344528
rect 69768 340066 70058 340082
rect 69756 340060 70058 340066
rect 69808 340054 70058 340060
rect 70412 340054 70702 340082
rect 69756 340002 69808 340008
rect 70412 333985 70440 340054
rect 71332 338065 71360 340068
rect 71686 339960 71742 339969
rect 71742 339930 71820 339946
rect 71742 339924 71832 339930
rect 71742 339918 71780 339924
rect 71686 339895 71742 339904
rect 71780 339866 71832 339872
rect 71318 338056 71374 338065
rect 71318 337991 71374 338000
rect 71332 337385 71360 337991
rect 71318 337376 71374 337385
rect 71318 337311 71374 337320
rect 71976 336666 72004 340068
rect 72424 339924 72476 339930
rect 72424 339866 72476 339872
rect 71964 336660 72016 336666
rect 71964 336602 72016 336608
rect 70398 333976 70454 333985
rect 70398 333911 70454 333920
rect 70412 333305 70440 333911
rect 70398 333296 70454 333305
rect 70398 333231 70454 333240
rect 69204 329180 69256 329186
rect 69204 329122 69256 329128
rect 71044 326392 71096 326398
rect 71044 326334 71096 326340
rect 69204 316056 69256 316062
rect 69204 315998 69256 316004
rect 69110 311128 69166 311137
rect 69110 311063 69166 311072
rect 69020 300144 69072 300150
rect 69020 300086 69072 300092
rect 68926 298208 68982 298217
rect 68926 298143 68982 298152
rect 67638 291136 67694 291145
rect 67638 291071 67694 291080
rect 67652 290494 67680 291071
rect 67640 290488 67692 290494
rect 67640 290430 67692 290436
rect 67638 288824 67694 288833
rect 67638 288759 67694 288768
rect 67652 288454 67680 288759
rect 67640 288448 67692 288454
rect 67640 288390 67692 288396
rect 67730 288416 67786 288425
rect 67730 288351 67732 288360
rect 67784 288351 67786 288360
rect 67732 288322 67784 288328
rect 68192 288312 68244 288318
rect 68192 288254 68244 288260
rect 68204 288153 68232 288254
rect 68190 288144 68246 288153
rect 68190 288079 68246 288088
rect 68940 286113 68968 298143
rect 69112 292800 69164 292806
rect 69112 292742 69164 292748
rect 69124 287065 69152 292742
rect 69110 287056 69166 287065
rect 69110 286991 69166 287000
rect 68926 286104 68982 286113
rect 68926 286039 68982 286048
rect 67546 285424 67602 285433
rect 67546 285359 67602 285368
rect 67638 284472 67694 284481
rect 67638 284407 67694 284416
rect 67652 284374 67680 284407
rect 67640 284368 67692 284374
rect 67640 284310 67692 284316
rect 67732 284300 67784 284306
rect 67732 284242 67784 284248
rect 67744 283393 67772 284242
rect 68834 283792 68890 283801
rect 68834 283727 68890 283736
rect 67730 283384 67786 283393
rect 67730 283319 67786 283328
rect 67730 280528 67786 280537
rect 67730 280463 67786 280472
rect 67638 280392 67694 280401
rect 67638 280327 67694 280336
rect 67652 280294 67680 280327
rect 67640 280288 67692 280294
rect 67640 280230 67692 280236
rect 67744 280226 67772 280463
rect 67732 280220 67784 280226
rect 67732 280162 67784 280168
rect 67638 279168 67694 279177
rect 67638 279103 67694 279112
rect 67652 278798 67680 279103
rect 67640 278792 67692 278798
rect 67640 278734 67692 278740
rect 67638 277808 67694 277817
rect 67638 277743 67694 277752
rect 67652 277438 67680 277743
rect 68282 277672 68338 277681
rect 68282 277607 68338 277616
rect 67640 277432 67692 277438
rect 67640 277374 67692 277380
rect 67730 276448 67786 276457
rect 67730 276383 67786 276392
rect 67638 276312 67694 276321
rect 67638 276247 67694 276256
rect 67652 276146 67680 276247
rect 67640 276140 67692 276146
rect 67640 276082 67692 276088
rect 67744 276078 67772 276383
rect 67732 276072 67784 276078
rect 67732 276014 67784 276020
rect 67730 275088 67786 275097
rect 67730 275023 67786 275032
rect 67638 274952 67694 274961
rect 67638 274887 67694 274896
rect 67652 274786 67680 274887
rect 67640 274780 67692 274786
rect 67640 274722 67692 274728
rect 67744 274718 67772 275023
rect 67732 274712 67784 274718
rect 67732 274654 67784 274660
rect 67638 273320 67694 273329
rect 67638 273255 67640 273264
rect 67692 273255 67694 273264
rect 67640 273226 67692 273232
rect 67638 272368 67694 272377
rect 67638 272303 67694 272312
rect 67652 271930 67680 272303
rect 68098 272232 68154 272241
rect 68098 272167 68154 272176
rect 68112 271998 68140 272167
rect 68100 271992 68152 271998
rect 68100 271934 68152 271940
rect 67640 271924 67692 271930
rect 67640 271866 67692 271872
rect 67730 271552 67786 271561
rect 67730 271487 67786 271496
rect 67640 271176 67692 271182
rect 67638 271144 67640 271153
rect 67692 271144 67694 271153
rect 67638 271079 67694 271088
rect 67744 270570 67772 271487
rect 67732 270564 67784 270570
rect 67732 270506 67784 270512
rect 67730 269648 67786 269657
rect 67730 269583 67786 269592
rect 67638 269512 67694 269521
rect 67638 269447 67694 269456
rect 67652 269142 67680 269447
rect 67744 269210 67772 269583
rect 67732 269204 67784 269210
rect 67732 269146 67784 269152
rect 67640 269136 67692 269142
rect 67640 269078 67692 269084
rect 67732 269068 67784 269074
rect 67732 269010 67784 269016
rect 67454 268832 67510 268841
rect 67454 268767 67510 268776
rect 66904 262880 66956 262886
rect 66904 262822 66956 262828
rect 67362 245712 67418 245721
rect 67362 245647 67418 245656
rect 66168 243024 66220 243030
rect 66168 242966 66220 242972
rect 66076 241528 66128 241534
rect 66076 241470 66128 241476
rect 65984 224256 66036 224262
rect 65984 224198 66036 224204
rect 65892 196716 65944 196722
rect 65892 196658 65944 196664
rect 66088 191282 66116 241470
rect 66180 236774 66208 242966
rect 66168 236768 66220 236774
rect 66168 236710 66220 236716
rect 67376 200870 67404 245647
rect 67468 229906 67496 268767
rect 67744 268433 67772 269010
rect 67730 268424 67786 268433
rect 67730 268359 67786 268368
rect 67730 266928 67786 266937
rect 67730 266863 67786 266872
rect 67638 266792 67694 266801
rect 67638 266727 67694 266736
rect 67652 266558 67680 266727
rect 67640 266552 67692 266558
rect 67640 266494 67692 266500
rect 67744 266422 67772 266863
rect 67732 266416 67784 266422
rect 67732 266358 67784 266364
rect 67640 265668 67692 265674
rect 67640 265610 67692 265616
rect 67652 265441 67680 265610
rect 67730 265568 67786 265577
rect 67730 265503 67786 265512
rect 67638 265432 67694 265441
rect 67638 265367 67694 265376
rect 67744 264994 67772 265503
rect 67732 264988 67784 264994
rect 67732 264930 67784 264936
rect 67640 264920 67692 264926
rect 67638 264888 67640 264897
rect 67692 264888 67694 264897
rect 67638 264823 67694 264832
rect 67730 262848 67786 262857
rect 67730 262783 67786 262792
rect 67744 262342 67772 262783
rect 67732 262336 67784 262342
rect 67638 262304 67694 262313
rect 67732 262278 67784 262284
rect 67638 262239 67640 262248
rect 67692 262239 67694 262248
rect 67640 262210 67692 262216
rect 67730 261488 67786 261497
rect 67730 261423 67786 261432
rect 67744 260914 67772 261423
rect 67732 260908 67784 260914
rect 67732 260850 67784 260856
rect 67640 260840 67692 260846
rect 67638 260808 67640 260817
rect 67692 260808 67694 260817
rect 67638 260743 67694 260752
rect 67638 259584 67694 259593
rect 67638 259519 67694 259528
rect 67652 259486 67680 259519
rect 67640 259480 67692 259486
rect 67640 259422 67692 259428
rect 67730 258632 67786 258641
rect 67730 258567 67786 258576
rect 67638 258224 67694 258233
rect 67638 258159 67640 258168
rect 67692 258159 67694 258168
rect 67640 258130 67692 258136
rect 67744 258126 67772 258567
rect 67732 258120 67784 258126
rect 67732 258062 67784 258068
rect 67730 257272 67786 257281
rect 67730 257207 67786 257216
rect 67638 256864 67694 256873
rect 67638 256799 67640 256808
rect 67692 256799 67694 256808
rect 67640 256770 67692 256776
rect 67744 256766 67772 257207
rect 67732 256760 67784 256766
rect 67732 256702 67784 256708
rect 67638 255912 67694 255921
rect 67638 255847 67694 255856
rect 67652 255406 67680 255847
rect 67640 255400 67692 255406
rect 67640 255342 67692 255348
rect 67730 255368 67786 255377
rect 67730 255303 67732 255312
rect 67784 255303 67786 255312
rect 67732 255274 67784 255280
rect 67640 255264 67692 255270
rect 67638 255232 67640 255241
rect 67692 255232 67694 255241
rect 67638 255167 67694 255176
rect 67640 254584 67692 254590
rect 67638 254552 67640 254561
rect 67692 254552 67694 254561
rect 67638 254487 67694 254496
rect 68098 252648 68154 252657
rect 68098 252583 68154 252592
rect 67638 251832 67694 251841
rect 67638 251767 67694 251776
rect 67652 251258 67680 251767
rect 67640 251252 67692 251258
rect 67640 251194 67692 251200
rect 67730 250472 67786 250481
rect 67730 250407 67786 250416
rect 67638 249928 67694 249937
rect 67744 249898 67772 250407
rect 67638 249863 67694 249872
rect 67732 249892 67784 249898
rect 67652 249830 67680 249863
rect 67732 249834 67784 249840
rect 67640 249824 67692 249830
rect 67640 249766 67692 249772
rect 67730 249112 67786 249121
rect 68112 249082 68140 252583
rect 68296 249150 68324 277607
rect 68284 249144 68336 249150
rect 68284 249086 68336 249092
rect 67730 249047 67786 249056
rect 68100 249076 68152 249082
rect 67638 248568 67694 248577
rect 67638 248503 67640 248512
rect 67692 248503 67694 248512
rect 67640 248474 67692 248480
rect 67744 248470 67772 249047
rect 68100 249018 68152 249024
rect 67732 248464 67784 248470
rect 67732 248406 67784 248412
rect 67730 247752 67786 247761
rect 67730 247687 67786 247696
rect 67638 247208 67694 247217
rect 67744 247178 67772 247687
rect 67638 247143 67694 247152
rect 67732 247172 67784 247178
rect 67652 247110 67680 247143
rect 67732 247114 67784 247120
rect 67640 247104 67692 247110
rect 67640 247046 67692 247052
rect 67638 244624 67694 244633
rect 67638 244559 67694 244568
rect 67652 244322 67680 244559
rect 67640 244316 67692 244322
rect 67640 244258 67692 244264
rect 67730 243672 67786 243681
rect 67730 243607 67786 243616
rect 67638 243264 67694 243273
rect 67638 243199 67694 243208
rect 67652 242962 67680 243199
rect 67744 243030 67772 243607
rect 67732 243024 67784 243030
rect 67732 242966 67784 242972
rect 67640 242956 67692 242962
rect 67640 242898 67692 242904
rect 68190 241632 68246 241641
rect 68190 241567 68246 241576
rect 68204 241534 68232 241567
rect 68192 241528 68244 241534
rect 68192 241470 68244 241476
rect 67638 240952 67694 240961
rect 67638 240887 67694 240896
rect 67652 234569 67680 240887
rect 68848 239465 68876 283727
rect 69216 282169 69244 315998
rect 69846 296848 69902 296857
rect 69846 296783 69902 296792
rect 69860 290873 69888 296783
rect 70676 296744 70728 296750
rect 70676 296686 70728 296692
rect 70032 294704 70084 294710
rect 70032 294646 70084 294652
rect 70044 291924 70072 294646
rect 70688 291963 70716 296686
rect 71056 292369 71084 326334
rect 72436 315314 72464 339866
rect 73280 339810 73308 340068
rect 73280 339782 73384 339810
rect 72516 336660 72568 336666
rect 72516 336602 72568 336608
rect 72528 324970 72556 336602
rect 73356 336462 73384 339782
rect 73908 339425 73936 340068
rect 73894 339416 73950 339425
rect 73894 339351 73950 339360
rect 73908 338065 73936 339351
rect 73894 338056 73950 338065
rect 73894 337991 73950 338000
rect 74446 338056 74502 338065
rect 74446 337991 74502 338000
rect 73344 336456 73396 336462
rect 73344 336398 73396 336404
rect 73356 336025 73384 336398
rect 73342 336016 73398 336025
rect 73342 335951 73398 335960
rect 72516 324964 72568 324970
rect 72516 324906 72568 324912
rect 73160 323604 73212 323610
rect 73160 323546 73212 323552
rect 72516 316736 72568 316742
rect 72516 316678 72568 316684
rect 72424 315308 72476 315314
rect 72424 315250 72476 315256
rect 71780 300960 71832 300966
rect 71780 300902 71832 300908
rect 71320 294364 71372 294370
rect 71320 294306 71372 294312
rect 71042 292360 71098 292369
rect 71042 292295 71098 292304
rect 71332 291963 71360 294306
rect 71792 291977 71820 300902
rect 72528 294370 72556 316678
rect 72608 295316 72660 295322
rect 72608 295258 72660 295264
rect 72516 294364 72568 294370
rect 72516 294306 72568 294312
rect 71792 291949 71990 291977
rect 72620 291963 72648 295258
rect 73172 294370 73200 323546
rect 74460 308514 74488 337991
rect 74552 337890 74580 340068
rect 75840 339454 75868 340068
rect 75918 339688 75974 339697
rect 75918 339623 75974 339632
rect 75184 339448 75236 339454
rect 75184 339390 75236 339396
rect 75828 339448 75880 339454
rect 75828 339390 75880 339396
rect 74540 337884 74592 337890
rect 74540 337826 74592 337832
rect 74448 308508 74500 308514
rect 74448 308450 74500 308456
rect 74540 306400 74592 306406
rect 74540 306342 74592 306348
rect 73252 303816 73304 303822
rect 73252 303758 73304 303764
rect 73160 294364 73212 294370
rect 73160 294306 73212 294312
rect 73264 291963 73292 303758
rect 73620 294364 73672 294370
rect 73620 294306 73672 294312
rect 73632 291977 73660 294306
rect 73632 291949 73922 291977
rect 74552 291963 74580 306342
rect 75196 302938 75224 339390
rect 75276 337884 75328 337890
rect 75276 337826 75328 337832
rect 75288 318102 75316 337826
rect 75276 318096 75328 318102
rect 75276 318038 75328 318044
rect 75932 312497 75960 339623
rect 76484 337958 76512 340068
rect 77128 339697 77156 340068
rect 77114 339688 77170 339697
rect 77114 339623 77170 339632
rect 78416 339522 78444 340068
rect 78404 339516 78456 339522
rect 78404 339458 78456 339464
rect 77944 338904 77996 338910
rect 77944 338846 77996 338852
rect 76472 337952 76524 337958
rect 76472 337894 76524 337900
rect 76484 335354 76512 337894
rect 76484 335326 76604 335354
rect 76576 326534 76604 335326
rect 76564 326528 76616 326534
rect 76564 326470 76616 326476
rect 75918 312488 75974 312497
rect 75918 312423 75974 312432
rect 75920 309188 75972 309194
rect 75920 309130 75972 309136
rect 75276 303000 75328 303006
rect 75276 302942 75328 302948
rect 75184 302932 75236 302938
rect 75184 302874 75236 302880
rect 75288 295322 75316 302942
rect 75276 295316 75328 295322
rect 75276 295258 75328 295264
rect 75826 294400 75882 294409
rect 75826 294335 75882 294344
rect 75184 292732 75236 292738
rect 75184 292674 75236 292680
rect 75196 291963 75224 292674
rect 75840 291963 75868 294335
rect 75932 291977 75960 309130
rect 77298 299568 77354 299577
rect 77298 299503 77354 299512
rect 77116 294636 77168 294642
rect 77116 294578 77168 294584
rect 75932 291949 76498 291977
rect 77128 291963 77156 294578
rect 77312 291977 77340 299503
rect 77956 294273 77984 338846
rect 78416 338842 78444 339458
rect 78404 338836 78456 338842
rect 78404 338778 78456 338784
rect 79060 338094 79088 340068
rect 79658 339810 79686 340068
rect 79336 339782 79686 339810
rect 79048 338088 79100 338094
rect 79048 338030 79100 338036
rect 79060 337482 79088 338030
rect 79048 337476 79100 337482
rect 79048 337418 79100 337424
rect 78034 337376 78090 337385
rect 78034 337311 78090 337320
rect 78048 327758 78076 337311
rect 79336 336530 79364 339782
rect 79324 336524 79376 336530
rect 79324 336466 79376 336472
rect 78036 327752 78088 327758
rect 78036 327694 78088 327700
rect 79336 306374 79364 336466
rect 80992 335102 81020 340068
rect 81636 335306 81664 340068
rect 82280 338094 82308 340068
rect 83522 339810 83550 340068
rect 83476 339782 83550 339810
rect 82268 338088 82320 338094
rect 82268 338030 82320 338036
rect 83476 336598 83504 339782
rect 84212 338026 84240 340068
rect 84200 338020 84252 338026
rect 84200 337962 84252 337968
rect 84856 337550 84884 340068
rect 86160 339810 86188 340068
rect 86160 339782 86264 339810
rect 84844 337544 84896 337550
rect 84844 337486 84896 337492
rect 83464 336592 83516 336598
rect 83464 336534 83516 336540
rect 81624 335300 81676 335306
rect 81624 335242 81676 335248
rect 80980 335096 81032 335102
rect 80980 335038 81032 335044
rect 80992 330449 81020 335038
rect 81636 334014 81664 335242
rect 81624 334008 81676 334014
rect 81624 333950 81676 333956
rect 82084 334008 82136 334014
rect 82084 333950 82136 333956
rect 80978 330440 81034 330449
rect 80978 330375 81034 330384
rect 82096 325038 82124 333950
rect 82084 325032 82136 325038
rect 82084 324974 82136 324980
rect 80060 314016 80112 314022
rect 80060 313958 80112 313964
rect 79336 306346 79456 306374
rect 79230 302288 79286 302297
rect 79230 302223 79286 302232
rect 77942 294264 77998 294273
rect 77942 294199 77998 294208
rect 77312 291949 77786 291977
rect 77956 291938 77984 294199
rect 79048 294092 79100 294098
rect 79048 294034 79100 294040
rect 79060 291963 79088 294034
rect 79244 291938 79272 302223
rect 79428 293185 79456 306346
rect 79414 293176 79470 293185
rect 79414 293111 79470 293120
rect 80072 291977 80100 313958
rect 81440 313336 81492 313342
rect 81440 313278 81492 313284
rect 81452 306374 81480 313278
rect 83476 308446 83504 336534
rect 86236 333946 86264 339782
rect 86788 335238 86816 340068
rect 87432 339454 87460 340068
rect 87420 339448 87472 339454
rect 87420 339390 87472 339396
rect 87696 339448 87748 339454
rect 87696 339390 87748 339396
rect 87604 338768 87656 338774
rect 87604 338710 87656 338716
rect 86776 335232 86828 335238
rect 86776 335174 86828 335180
rect 86788 334694 86816 335174
rect 86316 334688 86368 334694
rect 86316 334630 86368 334636
rect 86776 334688 86828 334694
rect 86776 334630 86828 334636
rect 86224 333940 86276 333946
rect 86224 333882 86276 333888
rect 84292 316124 84344 316130
rect 84292 316066 84344 316072
rect 83464 308440 83516 308446
rect 83464 308382 83516 308388
rect 81452 306346 81940 306374
rect 81532 301164 81584 301170
rect 81532 301106 81584 301112
rect 80978 296984 81034 296993
rect 80978 296919 81034 296928
rect 80072 291949 80362 291977
rect 80992 291963 81020 296919
rect 81544 291977 81572 301106
rect 81544 291949 81650 291977
rect 81912 291938 81940 306346
rect 83556 296948 83608 296954
rect 83556 296890 83608 296896
rect 82912 295656 82964 295662
rect 82912 295598 82964 295604
rect 82924 291963 82952 295598
rect 83568 291963 83596 296890
rect 84304 294370 84332 316066
rect 84384 309936 84436 309942
rect 84384 309878 84436 309884
rect 84292 294364 84344 294370
rect 84292 294306 84344 294312
rect 84396 291938 84424 309878
rect 85580 305108 85632 305114
rect 85580 305050 85632 305056
rect 85212 294364 85264 294370
rect 85212 294306 85264 294312
rect 85224 291977 85252 294306
rect 85224 291949 85514 291977
rect 85592 291938 85620 305050
rect 86236 300218 86264 333882
rect 86328 322250 86356 334630
rect 86316 322244 86368 322250
rect 86316 322186 86368 322192
rect 87616 311234 87644 338710
rect 87708 333334 87736 339390
rect 87696 333328 87748 333334
rect 87696 333270 87748 333276
rect 88720 329798 88748 340068
rect 89318 339810 89346 340068
rect 88996 339782 89346 339810
rect 88996 331226 89024 339782
rect 88984 331220 89036 331226
rect 88984 331162 89036 331168
rect 88708 329792 88760 329798
rect 88708 329734 88760 329740
rect 87604 311228 87656 311234
rect 87604 311170 87656 311176
rect 88996 309777 89024 331162
rect 90008 321570 90036 340068
rect 89996 321564 90048 321570
rect 89996 321506 90048 321512
rect 91296 318782 91324 340068
rect 91940 327894 91968 340068
rect 92480 336728 92532 336734
rect 92480 336670 92532 336676
rect 92492 336054 92520 336670
rect 92480 336048 92532 336054
rect 92480 335990 92532 335996
rect 92584 329730 92612 340068
rect 93124 338836 93176 338842
rect 93124 338778 93176 338784
rect 92572 329724 92624 329730
rect 92572 329666 92624 329672
rect 91928 327888 91980 327894
rect 91928 327830 91980 327836
rect 91284 318776 91336 318782
rect 91284 318718 91336 318724
rect 91100 314696 91152 314702
rect 91100 314638 91152 314644
rect 91112 314022 91140 314638
rect 93136 314022 93164 338778
rect 93228 336054 93256 340068
rect 93952 337544 94004 337550
rect 93952 337486 94004 337492
rect 93216 336048 93268 336054
rect 93216 335990 93268 335996
rect 93768 319592 93820 319598
rect 93768 319534 93820 319540
rect 91100 314016 91152 314022
rect 91100 313958 91152 313964
rect 93124 314016 93176 314022
rect 93124 313958 93176 313964
rect 88982 309768 89038 309777
rect 88982 309703 89038 309712
rect 88340 307828 88392 307834
rect 88340 307770 88392 307776
rect 87512 302320 87564 302326
rect 87512 302262 87564 302268
rect 86316 302252 86368 302258
rect 86316 302194 86368 302200
rect 86224 300212 86276 300218
rect 86224 300154 86276 300160
rect 86328 291977 86356 302194
rect 87420 298376 87472 298382
rect 87420 298318 87472 298324
rect 86328 291949 86802 291977
rect 87432 291963 87460 298318
rect 87524 291977 87552 302262
rect 87524 291949 88090 291977
rect 88352 291938 88380 307770
rect 92664 303884 92716 303890
rect 92664 303826 92716 303832
rect 90272 301232 90324 301238
rect 90272 301174 90324 301180
rect 88984 299532 89036 299538
rect 88984 299474 89036 299480
rect 88996 291977 89024 299474
rect 89994 295488 90050 295497
rect 89994 295423 90050 295432
rect 88996 291949 89378 291977
rect 90008 291963 90036 295423
rect 90284 291977 90312 301174
rect 91928 295520 91980 295526
rect 91928 295462 91980 295468
rect 91284 294772 91336 294778
rect 91284 294714 91336 294720
rect 90284 291949 90666 291977
rect 91296 291963 91324 294714
rect 91940 291963 91968 295462
rect 92572 292596 92624 292602
rect 92572 292538 92624 292544
rect 92584 291963 92612 292538
rect 92676 291977 92704 303826
rect 93780 292602 93808 319534
rect 93964 294370 93992 337486
rect 94516 335170 94544 340068
rect 95114 339810 95142 340068
rect 94608 339782 95142 339810
rect 94504 335164 94556 335170
rect 94504 335106 94556 335112
rect 94608 307766 94636 339782
rect 95148 333328 95200 333334
rect 95148 333270 95200 333276
rect 94228 307760 94280 307766
rect 94228 307702 94280 307708
rect 94596 307760 94648 307766
rect 94596 307702 94648 307708
rect 94240 307193 94268 307702
rect 94226 307184 94282 307193
rect 94226 307119 94282 307128
rect 95160 303686 95188 333270
rect 95804 324290 95832 340068
rect 97092 333946 97120 340068
rect 97736 339522 97764 340068
rect 97724 339516 97776 339522
rect 97724 339458 97776 339464
rect 97080 333940 97132 333946
rect 97080 333882 97132 333888
rect 97092 332790 97120 333882
rect 97080 332784 97132 332790
rect 97080 332726 97132 332732
rect 95792 324284 95844 324290
rect 95792 324226 95844 324232
rect 97736 305658 97764 339458
rect 97908 332784 97960 332790
rect 97908 332726 97960 332732
rect 97920 307154 97948 332726
rect 97908 307148 97960 307154
rect 97908 307090 97960 307096
rect 98380 306338 98408 340068
rect 99668 339386 99696 340068
rect 99656 339380 99708 339386
rect 99656 339322 99708 339328
rect 100312 338026 100340 340068
rect 100668 339380 100720 339386
rect 100668 339322 100720 339328
rect 100300 338020 100352 338026
rect 100300 337962 100352 337968
rect 100024 334688 100076 334694
rect 100024 334630 100076 334636
rect 98644 331968 98696 331974
rect 98644 331910 98696 331916
rect 98368 306332 98420 306338
rect 98368 306274 98420 306280
rect 97724 305652 97776 305658
rect 97724 305594 97776 305600
rect 98656 303958 98684 331910
rect 98644 303952 98696 303958
rect 98644 303894 98696 303900
rect 98656 303686 98684 303894
rect 94044 303680 94096 303686
rect 94044 303622 94096 303628
rect 95148 303680 95200 303686
rect 95148 303622 95200 303628
rect 98000 303680 98052 303686
rect 98000 303622 98052 303628
rect 98644 303680 98696 303686
rect 98644 303622 98696 303628
rect 93952 294364 94004 294370
rect 93952 294306 94004 294312
rect 93860 292868 93912 292874
rect 93860 292810 93912 292816
rect 93768 292596 93820 292602
rect 93768 292538 93820 292544
rect 92676 291949 93242 291977
rect 93872 291963 93900 292810
rect 94056 291977 94084 303622
rect 97356 299600 97408 299606
rect 97356 299542 97408 299548
rect 94780 294364 94832 294370
rect 94780 294306 94832 294312
rect 94056 291949 94530 291977
rect 94792 291938 94820 294306
rect 97080 294160 97132 294166
rect 95790 294128 95846 294137
rect 97080 294102 97132 294108
rect 95790 294063 95846 294072
rect 95804 291963 95832 294063
rect 96436 294024 96488 294030
rect 96436 293966 96488 293972
rect 96448 291963 96476 293966
rect 97092 292670 97120 294102
rect 97080 292664 97132 292670
rect 97080 292606 97132 292612
rect 97092 291963 97120 292606
rect 97368 291938 97396 299542
rect 98012 291977 98040 303622
rect 98644 301096 98696 301102
rect 98644 301038 98696 301044
rect 98012 291949 98394 291977
rect 98656 291938 98684 301038
rect 100036 296886 100064 334630
rect 100680 304638 100708 339322
rect 100956 320142 100984 340068
rect 100944 320136 100996 320142
rect 100944 320078 100996 320084
rect 101404 319524 101456 319530
rect 101404 319466 101456 319472
rect 101416 311302 101444 319466
rect 102244 317422 102272 340068
rect 102888 335170 102916 340068
rect 103532 337618 103560 340068
rect 104820 339425 104848 340068
rect 104806 339416 104862 339425
rect 104806 339351 104862 339360
rect 104820 338881 104848 339351
rect 104806 338872 104862 338881
rect 104806 338807 104862 338816
rect 103520 337612 103572 337618
rect 103520 337554 103572 337560
rect 104164 336048 104216 336054
rect 104164 335990 104216 335996
rect 102876 335164 102928 335170
rect 102876 335106 102928 335112
rect 103428 335164 103480 335170
rect 103428 335106 103480 335112
rect 102232 317416 102284 317422
rect 102232 317358 102284 317364
rect 101404 311296 101456 311302
rect 101404 311238 101456 311244
rect 100668 304632 100720 304638
rect 100668 304574 100720 304580
rect 100852 299668 100904 299674
rect 100852 299610 100904 299616
rect 100024 296880 100076 296886
rect 100024 296822 100076 296828
rect 99656 296812 99708 296818
rect 99656 296754 99708 296760
rect 99668 291963 99696 296754
rect 100036 294370 100064 296822
rect 100024 294364 100076 294370
rect 100024 294306 100076 294312
rect 100864 291977 100892 299610
rect 103440 296002 103468 335106
rect 104176 297430 104204 335990
rect 105464 331226 105492 340068
rect 106124 339810 106152 340068
rect 106124 339782 106228 339810
rect 106200 338094 106228 339782
rect 107396 339289 107424 340068
rect 107382 339280 107438 339289
rect 107382 339215 107438 339224
rect 107566 339280 107622 339289
rect 107566 339215 107622 339224
rect 106188 338088 106240 338094
rect 106188 338030 106240 338036
rect 105452 331220 105504 331226
rect 105452 331162 105504 331168
rect 106096 327956 106148 327962
rect 106096 327898 106148 327904
rect 104256 316056 104308 316062
rect 104256 315998 104308 316004
rect 104268 309126 104296 315998
rect 104900 309868 104952 309874
rect 104900 309810 104952 309816
rect 104256 309120 104308 309126
rect 104256 309062 104308 309068
rect 104256 304632 104308 304638
rect 104256 304574 104308 304580
rect 104164 297424 104216 297430
rect 104164 297366 104216 297372
rect 103428 295996 103480 296002
rect 103428 295938 103480 295944
rect 104268 295594 104296 304574
rect 104256 295588 104308 295594
rect 104256 295530 104308 295536
rect 104808 295588 104860 295594
rect 104808 295530 104860 295536
rect 102232 295452 102284 295458
rect 102232 295394 102284 295400
rect 101588 294364 101640 294370
rect 101588 294306 101640 294312
rect 100864 291949 100970 291977
rect 101600 291963 101628 294306
rect 102244 291963 102272 295394
rect 102876 294228 102928 294234
rect 102876 294170 102928 294176
rect 102888 291963 102916 294170
rect 103520 292664 103572 292670
rect 103520 292606 103572 292612
rect 103532 291963 103560 292606
rect 104820 291963 104848 295530
rect 104912 294370 104940 309810
rect 106108 301374 106136 327898
rect 106200 307086 106228 338030
rect 106188 307080 106240 307086
rect 106188 307022 106240 307028
rect 106832 303068 106884 303074
rect 106832 303010 106884 303016
rect 104992 301368 105044 301374
rect 104992 301310 105044 301316
rect 106096 301368 106148 301374
rect 106096 301310 106148 301316
rect 104900 294364 104952 294370
rect 104900 294306 104952 294312
rect 105004 291938 105032 301310
rect 106108 300898 106136 301310
rect 106096 300892 106148 300898
rect 106096 300834 106148 300840
rect 106740 298240 106792 298246
rect 106740 298182 106792 298188
rect 105820 294364 105872 294370
rect 105820 294306 105872 294312
rect 105832 291977 105860 294306
rect 105832 291949 106122 291977
rect 106752 291963 106780 298182
rect 106844 291977 106872 303010
rect 107580 297498 107608 339215
rect 108040 336734 108068 340068
rect 108638 339810 108666 340068
rect 108316 339782 108666 339810
rect 108028 336728 108080 336734
rect 108028 336670 108080 336676
rect 108040 329118 108068 336670
rect 108316 332586 108344 339782
rect 109972 335238 110000 340068
rect 109960 335232 110012 335238
rect 109960 335174 110012 335180
rect 108304 332580 108356 332586
rect 108304 332522 108356 332528
rect 108028 329112 108080 329118
rect 108028 329054 108080 329060
rect 108316 316742 108344 332522
rect 110616 322930 110644 340068
rect 110604 322924 110656 322930
rect 110604 322866 110656 322872
rect 111260 318714 111288 340068
rect 112548 327078 112576 340068
rect 113208 339833 113236 340068
rect 113194 339824 113250 339833
rect 113192 339768 113194 339810
rect 113192 339759 113250 339768
rect 112536 327072 112588 327078
rect 112536 327014 112588 327020
rect 111248 318708 111300 318714
rect 111248 318650 111300 318656
rect 108304 316736 108356 316742
rect 108304 316678 108356 316684
rect 113192 316130 113220 339759
rect 113836 337958 113864 340068
rect 113824 337952 113876 337958
rect 113824 337894 113876 337900
rect 113836 333334 113864 337894
rect 114468 337612 114520 337618
rect 114468 337554 114520 337560
rect 114480 336054 114508 337554
rect 115124 336666 115152 340068
rect 115216 340054 115782 340082
rect 115112 336660 115164 336666
rect 115112 336602 115164 336608
rect 114468 336048 114520 336054
rect 114468 335990 114520 335996
rect 115216 335306 115244 340054
rect 115296 336660 115348 336666
rect 115296 336602 115348 336608
rect 115204 335300 115256 335306
rect 115204 335242 115256 335248
rect 113824 333328 113876 333334
rect 113824 333270 113876 333276
rect 115204 330540 115256 330546
rect 115204 330482 115256 330488
rect 113180 316124 113232 316130
rect 113180 316066 113232 316072
rect 113192 309806 113220 316066
rect 113180 309800 113232 309806
rect 113180 309742 113232 309748
rect 113824 307080 113876 307086
rect 113824 307022 113876 307028
rect 108394 301608 108450 301617
rect 108394 301543 108450 301552
rect 107568 297492 107620 297498
rect 107568 297434 107620 297440
rect 108028 294092 108080 294098
rect 108028 294034 108080 294040
rect 106844 291949 107410 291977
rect 108040 291963 108068 294034
rect 108408 291977 108436 301543
rect 109040 301028 109092 301034
rect 109040 300970 109092 300976
rect 109052 291977 109080 300970
rect 112444 299736 112496 299742
rect 112444 299678 112496 299684
rect 111248 298172 111300 298178
rect 111248 298114 111300 298120
rect 110604 296880 110656 296886
rect 110604 296822 110656 296828
rect 109960 294296 110012 294302
rect 109960 294238 110012 294244
rect 108408 291949 108698 291977
rect 109052 291949 109342 291977
rect 109972 291963 110000 294238
rect 110616 291963 110644 296822
rect 111260 291963 111288 298114
rect 112456 294710 112484 299678
rect 113836 298450 113864 307022
rect 114560 305040 114612 305046
rect 114560 304982 114612 304988
rect 113824 298444 113876 298450
rect 113824 298386 113876 298392
rect 113836 296714 113864 298386
rect 113744 296686 113864 296714
rect 112444 294704 112496 294710
rect 112444 294646 112496 294652
rect 111890 292768 111946 292777
rect 111890 292703 111946 292712
rect 111904 291963 111932 292703
rect 113744 291977 113772 296686
rect 114466 295352 114522 295361
rect 114466 295287 114522 295296
rect 113824 294024 113876 294030
rect 113824 293966 113876 293972
rect 113206 291949 113772 291977
rect 113836 291963 113864 293966
rect 114480 291963 114508 295287
rect 114572 291977 114600 304982
rect 115216 296714 115244 330482
rect 115308 319598 115336 336602
rect 115952 323610 115980 369922
rect 116044 327962 116072 383959
rect 116136 370025 116164 392430
rect 116228 383625 116256 487902
rect 117228 485784 117280 485790
rect 117226 485752 117228 485761
rect 117280 485752 117282 485761
rect 117226 485687 117282 485696
rect 117332 484362 117360 575486
rect 117424 534886 117452 582626
rect 117964 567248 118016 567254
rect 117964 567190 118016 567196
rect 117412 534880 117464 534886
rect 117412 534822 117464 534828
rect 117320 484356 117372 484362
rect 117320 484298 117372 484304
rect 117688 482996 117740 483002
rect 117688 482938 117740 482944
rect 117320 474020 117372 474026
rect 117320 473962 117372 473968
rect 116584 465860 116636 465866
rect 116584 465802 116636 465808
rect 116214 383616 116270 383625
rect 116214 383551 116270 383560
rect 116228 382294 116256 383551
rect 116216 382288 116268 382294
rect 116216 382230 116268 382236
rect 116122 370016 116178 370025
rect 116122 369951 116178 369960
rect 116596 362030 116624 465802
rect 116676 465792 116728 465798
rect 116676 465734 116728 465740
rect 116688 462262 116716 465734
rect 116676 462256 116728 462262
rect 116676 462198 116728 462204
rect 117332 387705 117360 473962
rect 117502 398032 117558 398041
rect 117502 397967 117558 397976
rect 117318 387696 117374 387705
rect 117318 387631 117374 387640
rect 117412 387184 117464 387190
rect 117412 387126 117464 387132
rect 117228 385688 117280 385694
rect 117228 385630 117280 385636
rect 117240 383654 117268 385630
rect 117240 383626 117360 383654
rect 117332 376145 117360 383626
rect 117318 376136 117374 376145
rect 117318 376071 117374 376080
rect 117424 363662 117452 387126
rect 117412 363656 117464 363662
rect 117412 363598 117464 363604
rect 117424 363225 117452 363598
rect 117410 363216 117466 363225
rect 117410 363151 117466 363160
rect 116584 362024 116636 362030
rect 116584 361966 116636 361972
rect 117320 362024 117372 362030
rect 117320 361966 117372 361972
rect 117332 357105 117360 361966
rect 117412 357400 117464 357406
rect 117412 357342 117464 357348
rect 117318 357096 117374 357105
rect 117318 357031 117374 357040
rect 117424 348945 117452 357342
rect 117516 355745 117544 397967
rect 117596 392828 117648 392834
rect 117596 392770 117648 392776
rect 117608 364334 117636 392770
rect 117700 384985 117728 482938
rect 117976 476134 118004 567190
rect 118712 493338 118740 586502
rect 118792 582616 118844 582622
rect 118792 582558 118844 582564
rect 118804 497486 118832 582558
rect 120080 550656 120132 550662
rect 120080 550598 120132 550604
rect 119344 545760 119396 545766
rect 119344 545702 119396 545708
rect 118884 498840 118936 498846
rect 118884 498782 118936 498788
rect 118792 497480 118844 497486
rect 118792 497422 118844 497428
rect 118700 493332 118752 493338
rect 118700 493274 118752 493280
rect 118792 491224 118844 491230
rect 118792 491166 118844 491172
rect 118700 477556 118752 477562
rect 118700 477498 118752 477504
rect 117964 476128 118016 476134
rect 117964 476070 118016 476076
rect 117976 475998 118004 476070
rect 117964 475992 118016 475998
rect 117964 475934 118016 475940
rect 118712 392494 118740 477498
rect 118804 422278 118832 491166
rect 118896 438190 118924 498782
rect 119356 454073 119384 545702
rect 120092 458182 120120 550598
rect 120184 494766 120212 586570
rect 121472 585410 121500 587114
rect 122840 585472 122892 585478
rect 122840 585414 122892 585420
rect 121460 585404 121512 585410
rect 121460 585346 121512 585352
rect 120264 582752 120316 582758
rect 120264 582694 120316 582700
rect 120172 494760 120224 494766
rect 120172 494702 120224 494708
rect 120276 492658 120304 582694
rect 120448 497548 120500 497554
rect 120448 497490 120500 497496
rect 120356 494828 120408 494834
rect 120356 494770 120408 494776
rect 120264 492652 120316 492658
rect 120264 492594 120316 492600
rect 120276 492386 120304 492594
rect 120264 492380 120316 492386
rect 120264 492322 120316 492328
rect 120080 458176 120132 458182
rect 120080 458118 120132 458124
rect 118974 454064 119030 454073
rect 118974 453999 118976 454008
rect 119028 453999 119030 454008
rect 119342 454064 119398 454073
rect 119342 453999 119398 454008
rect 118976 453970 119028 453976
rect 120368 438977 120396 494770
rect 120460 439550 120488 497490
rect 121472 489870 121500 585346
rect 121552 585200 121604 585206
rect 121552 585142 121604 585148
rect 121564 493406 121592 585142
rect 121644 566500 121696 566506
rect 121644 566442 121696 566448
rect 121656 496194 121684 566442
rect 122104 538892 122156 538898
rect 122104 538834 122156 538840
rect 122116 538286 122144 538834
rect 122104 538280 122156 538286
rect 122104 538222 122156 538228
rect 121644 496188 121696 496194
rect 121644 496130 121696 496136
rect 121644 494964 121696 494970
rect 121644 494906 121696 494912
rect 121552 493400 121604 493406
rect 121552 493342 121604 493348
rect 121552 492380 121604 492386
rect 121552 492322 121604 492328
rect 121460 489864 121512 489870
rect 121460 489806 121512 489812
rect 121460 475380 121512 475386
rect 121460 475322 121512 475328
rect 120724 462256 120776 462262
rect 120724 462198 120776 462204
rect 120448 439544 120500 439550
rect 120448 439486 120500 439492
rect 120354 438968 120410 438977
rect 120354 438903 120410 438912
rect 118884 438184 118936 438190
rect 118884 438126 118936 438132
rect 118792 422272 118844 422278
rect 118792 422214 118844 422220
rect 118700 392488 118752 392494
rect 118700 392430 118752 392436
rect 118804 389978 118832 422214
rect 120172 391332 120224 391338
rect 120172 391274 120224 391280
rect 120080 390788 120132 390794
rect 120080 390730 120132 390736
rect 118792 389972 118844 389978
rect 118792 389914 118844 389920
rect 118804 389502 118832 389914
rect 120092 389910 120120 390730
rect 120080 389904 120132 389910
rect 120080 389846 120132 389852
rect 118792 389496 118844 389502
rect 118792 389438 118844 389444
rect 119436 388068 119488 388074
rect 119436 388010 119488 388016
rect 119344 388000 119396 388006
rect 119344 387942 119396 387948
rect 118700 387252 118752 387258
rect 118700 387194 118752 387200
rect 117686 384976 117742 384985
rect 117686 384911 117742 384920
rect 118606 384976 118662 384985
rect 118606 384911 118662 384920
rect 118620 384334 118648 384911
rect 118608 384328 118660 384334
rect 118608 384270 118660 384276
rect 118606 382256 118662 382265
rect 118606 382191 118608 382200
rect 118660 382191 118662 382200
rect 118608 382162 118660 382168
rect 118608 381608 118660 381614
rect 118606 381576 118608 381585
rect 118660 381576 118662 381585
rect 118606 381511 118662 381520
rect 118606 380896 118662 380905
rect 118606 380831 118662 380840
rect 118620 379642 118648 380831
rect 118608 379636 118660 379642
rect 118608 379578 118660 379584
rect 118516 379568 118568 379574
rect 118514 379536 118516 379545
rect 118568 379536 118570 379545
rect 118514 379471 118570 379480
rect 118608 378888 118660 378894
rect 118606 378856 118608 378865
rect 118660 378856 118662 378865
rect 118606 378791 118662 378800
rect 117872 378208 117924 378214
rect 117870 378176 117872 378185
rect 117924 378176 117926 378185
rect 117870 378111 117926 378120
rect 118608 376848 118660 376854
rect 118606 376816 118608 376825
rect 118660 376816 118662 376825
rect 118606 376751 118662 376760
rect 118606 375456 118662 375465
rect 118606 375391 118608 375400
rect 118660 375391 118662 375400
rect 118608 375362 118660 375368
rect 118148 375352 118200 375358
rect 118148 375294 118200 375300
rect 118160 374105 118188 375294
rect 118146 374096 118202 374105
rect 118146 374031 118202 374040
rect 118330 373416 118386 373425
rect 118330 373351 118386 373360
rect 118344 372706 118372 373351
rect 118514 372736 118570 372745
rect 118332 372700 118384 372706
rect 118514 372671 118570 372680
rect 118332 372642 118384 372648
rect 118528 372638 118556 372671
rect 118516 372632 118568 372638
rect 118516 372574 118568 372580
rect 118146 371376 118202 371385
rect 118146 371311 118202 371320
rect 118160 371278 118188 371311
rect 118148 371272 118200 371278
rect 118148 371214 118200 371220
rect 118146 370016 118202 370025
rect 118146 369951 118202 369960
rect 118160 369918 118188 369951
rect 118148 369912 118200 369918
rect 118148 369854 118200 369860
rect 118606 368656 118662 368665
rect 118606 368591 118662 368600
rect 118620 368558 118648 368591
rect 118608 368552 118660 368558
rect 118608 368494 118660 368500
rect 118606 367976 118662 367985
rect 118606 367911 118662 367920
rect 118620 367878 118648 367911
rect 118608 367872 118660 367878
rect 118608 367814 118660 367820
rect 118606 367296 118662 367305
rect 118606 367231 118608 367240
rect 118660 367231 118662 367240
rect 118608 367202 118660 367208
rect 118608 366444 118660 366450
rect 118608 366386 118660 366392
rect 118620 365945 118648 366386
rect 118606 365936 118662 365945
rect 118606 365871 118662 365880
rect 118514 365256 118570 365265
rect 118514 365191 118570 365200
rect 118528 364410 118556 365191
rect 118608 365084 118660 365090
rect 118608 365026 118660 365032
rect 118620 364585 118648 365026
rect 118606 364576 118662 364585
rect 118606 364511 118662 364520
rect 118516 364404 118568 364410
rect 118516 364346 118568 364352
rect 117608 364306 117728 364334
rect 117502 355736 117558 355745
rect 117502 355671 117558 355680
rect 117504 354612 117556 354618
rect 117504 354554 117556 354560
rect 117516 354385 117544 354554
rect 117502 354376 117558 354385
rect 117502 354311 117558 354320
rect 117504 353252 117556 353258
rect 117504 353194 117556 353200
rect 117516 353025 117544 353194
rect 117502 353016 117558 353025
rect 117502 352951 117558 352960
rect 117700 351665 117728 364306
rect 118608 362908 118660 362914
rect 118608 362850 118660 362856
rect 118620 362545 118648 362850
rect 118606 362536 118662 362545
rect 118606 362471 118662 362480
rect 118608 362228 118660 362234
rect 118608 362170 118660 362176
rect 118620 361865 118648 362170
rect 118606 361856 118662 361865
rect 118606 361791 118662 361800
rect 118054 361176 118110 361185
rect 118054 361111 118110 361120
rect 118068 360262 118096 361111
rect 118056 360256 118108 360262
rect 118056 360198 118108 360204
rect 117964 360188 118016 360194
rect 117964 360130 118016 360136
rect 117976 359145 118004 360130
rect 118608 360120 118660 360126
rect 118608 360062 118660 360068
rect 118620 359825 118648 360062
rect 118606 359816 118662 359825
rect 118606 359751 118662 359760
rect 117962 359136 118018 359145
rect 117962 359071 118018 359080
rect 118608 358760 118660 358766
rect 118608 358702 118660 358708
rect 118620 358465 118648 358702
rect 118606 358456 118662 358465
rect 118606 358391 118662 358400
rect 118608 357400 118660 357406
rect 118608 357342 118660 357348
rect 118238 357096 118294 357105
rect 118238 357031 118294 357040
rect 118252 356726 118280 357031
rect 118240 356720 118292 356726
rect 118240 356662 118292 356668
rect 118620 356425 118648 357342
rect 118606 356416 118662 356425
rect 118606 356351 118662 356360
rect 118608 354680 118660 354686
rect 118608 354622 118660 354628
rect 118620 353705 118648 354622
rect 118606 353696 118662 353705
rect 118606 353631 118662 353640
rect 118056 351892 118108 351898
rect 118056 351834 118108 351840
rect 117686 351656 117742 351665
rect 117686 351591 117742 351600
rect 118068 350985 118096 351834
rect 118606 351656 118662 351665
rect 118606 351591 118662 351600
rect 118620 351218 118648 351591
rect 118608 351212 118660 351218
rect 118608 351154 118660 351160
rect 118054 350976 118110 350985
rect 118054 350911 118110 350920
rect 117502 350296 117558 350305
rect 117502 350231 117558 350240
rect 117516 349178 117544 350231
rect 117504 349172 117556 349178
rect 117504 349114 117556 349120
rect 117410 348936 117466 348945
rect 117410 348871 117466 348880
rect 118514 348936 118570 348945
rect 118514 348871 118570 348880
rect 118528 348430 118556 348871
rect 118516 348424 118568 348430
rect 118516 348366 118568 348372
rect 117962 348256 118018 348265
rect 117962 348191 118018 348200
rect 117976 345030 118004 348191
rect 118608 347744 118660 347750
rect 118608 347686 118660 347692
rect 118620 347585 118648 347686
rect 118606 347576 118662 347585
rect 118606 347511 118662 347520
rect 118608 346384 118660 346390
rect 118608 346326 118660 346332
rect 118514 346216 118570 346225
rect 118514 346151 118570 346160
rect 118528 345778 118556 346151
rect 118516 345772 118568 345778
rect 118516 345714 118568 345720
rect 117964 345024 118016 345030
rect 117964 344966 118016 344972
rect 117870 344856 117926 344865
rect 117870 344791 117926 344800
rect 117884 343670 117912 344791
rect 117872 343664 117924 343670
rect 117872 343606 117924 343612
rect 118054 342136 118110 342145
rect 118054 342071 118110 342080
rect 118068 340950 118096 342071
rect 118056 340944 118108 340950
rect 118056 340886 118108 340892
rect 117964 340876 118016 340882
rect 117964 340818 118016 340824
rect 117976 340105 118004 340818
rect 116122 340096 116178 340105
rect 116122 340031 116178 340040
rect 117962 340096 118018 340105
rect 117962 340031 118018 340040
rect 116032 327956 116084 327962
rect 116032 327898 116084 327904
rect 115940 323604 115992 323610
rect 115940 323546 115992 323552
rect 116136 320958 116164 340031
rect 118528 335354 118556 345714
rect 118620 345545 118648 346326
rect 118606 345536 118662 345545
rect 118606 345471 118662 345480
rect 118606 343496 118662 343505
rect 118606 343431 118662 343440
rect 118620 342922 118648 343431
rect 118608 342916 118660 342922
rect 118608 342858 118660 342864
rect 118606 342816 118662 342825
rect 118606 342751 118662 342760
rect 118620 342242 118648 342751
rect 118608 342236 118660 342242
rect 118608 342178 118660 342184
rect 118608 340808 118660 340814
rect 118606 340776 118608 340785
rect 118660 340776 118662 340785
rect 118606 340711 118662 340720
rect 118528 335326 118648 335354
rect 116124 320952 116176 320958
rect 116124 320894 116176 320900
rect 115296 319592 115348 319598
rect 115296 319534 115348 319540
rect 115296 318096 115348 318102
rect 115296 318038 115348 318044
rect 115308 305046 115336 318038
rect 116584 311296 116636 311302
rect 116584 311238 116636 311244
rect 115848 311160 115900 311166
rect 115848 311102 115900 311108
rect 115860 309942 115888 311102
rect 115848 309936 115900 309942
rect 115848 309878 115900 309884
rect 115296 305040 115348 305046
rect 115296 304982 115348 304988
rect 116596 303754 116624 311238
rect 115940 303748 115992 303754
rect 115940 303690 115992 303696
rect 116584 303748 116636 303754
rect 116584 303690 116636 303696
rect 115216 296686 115336 296714
rect 115308 292641 115336 296686
rect 115294 292632 115350 292641
rect 115294 292567 115350 292576
rect 115754 292632 115810 292641
rect 115754 292567 115810 292576
rect 114572 291949 115138 291977
rect 115768 291963 115796 292567
rect 115952 291977 115980 303690
rect 118330 298344 118386 298353
rect 118330 298279 118386 298288
rect 117044 295384 117096 295390
rect 117044 295326 117096 295332
rect 115952 291949 116426 291977
rect 117056 291963 117084 295326
rect 118344 291963 118372 298279
rect 118620 293078 118648 335326
rect 118712 318782 118740 387194
rect 119356 360913 119384 387942
rect 119448 376009 119476 388010
rect 119528 387932 119580 387938
rect 119528 387874 119580 387880
rect 119540 378826 119568 387874
rect 119528 378820 119580 378826
rect 119528 378762 119580 378768
rect 119528 377460 119580 377466
rect 119528 377402 119580 377408
rect 119540 376854 119568 377402
rect 119528 376848 119580 376854
rect 119528 376790 119580 376796
rect 119434 376000 119490 376009
rect 119434 375935 119490 375944
rect 119540 368393 119568 376790
rect 120184 373994 120212 391274
rect 120736 390794 120764 462198
rect 120816 396840 120868 396846
rect 120816 396782 120868 396788
rect 120724 390788 120776 390794
rect 120724 390730 120776 390736
rect 120092 373966 120212 373994
rect 119526 368384 119582 368393
rect 119526 368319 119582 368328
rect 119988 362228 120040 362234
rect 119988 362170 120040 362176
rect 119342 360904 119398 360913
rect 119342 360839 119398 360848
rect 118790 355736 118846 355745
rect 118790 355671 118846 355680
rect 118804 354006 118832 355671
rect 119344 355360 119396 355366
rect 119344 355302 119396 355308
rect 118792 354000 118844 354006
rect 118792 353942 118844 353948
rect 119356 338065 119384 355302
rect 119436 349172 119488 349178
rect 119436 349114 119488 349120
rect 119342 338056 119398 338065
rect 119342 337991 119398 338000
rect 119448 336666 119476 349114
rect 119436 336660 119488 336666
rect 119436 336602 119488 336608
rect 119448 334626 119476 336602
rect 119436 334620 119488 334626
rect 119436 334562 119488 334568
rect 118700 318776 118752 318782
rect 118700 318718 118752 318724
rect 118712 318102 118740 318718
rect 118700 318096 118752 318102
rect 118700 318038 118752 318044
rect 118700 307080 118752 307086
rect 118700 307022 118752 307028
rect 118712 306374 118740 307022
rect 118712 306346 119200 306374
rect 118608 293072 118660 293078
rect 118608 293014 118660 293020
rect 119066 292088 119122 292097
rect 119066 292023 119122 292032
rect 119080 291977 119108 292023
rect 117962 291952 118018 291961
rect 77956 291910 78418 291938
rect 79244 291910 79706 291938
rect 81912 291910 82282 291938
rect 84292 291916 84344 291922
rect 84226 291864 84292 291870
rect 84396 291910 84858 291938
rect 85592 291910 86146 291938
rect 88352 291910 88722 291938
rect 94792 291910 95162 291938
rect 97368 291910 97738 291938
rect 98656 291910 99026 291938
rect 104440 291916 104492 291922
rect 84226 291858 84344 291864
rect 104190 291864 104440 291870
rect 105004 291910 105466 291938
rect 112812 291916 112864 291922
rect 104190 291858 104492 291864
rect 112562 291864 112812 291870
rect 117714 291910 117962 291938
rect 119002 291949 119108 291977
rect 119172 291938 119200 306346
rect 119172 291910 119646 291938
rect 119712 291916 119764 291922
rect 117962 291887 118018 291896
rect 112562 291858 112864 291864
rect 119712 291858 119764 291864
rect 84226 291842 84332 291858
rect 104190 291842 104480 291858
rect 112562 291842 112852 291858
rect 119724 291310 119752 291858
rect 119712 291304 119764 291310
rect 119712 291246 119764 291252
rect 69846 290864 69902 290873
rect 69846 290799 69902 290808
rect 69202 282160 69258 282169
rect 69202 282095 69258 282104
rect 68926 263664 68982 263673
rect 68926 263599 68982 263608
rect 68834 239456 68890 239465
rect 68834 239391 68890 239400
rect 67638 234560 67694 234569
rect 67638 234495 67694 234504
rect 67456 229900 67508 229906
rect 67456 229842 67508 229848
rect 67364 200864 67416 200870
rect 67364 200806 67416 200812
rect 68940 199345 68968 263599
rect 120000 259350 120028 362170
rect 120092 335170 120120 373966
rect 120172 372700 120224 372706
rect 120172 372642 120224 372648
rect 120184 371210 120212 372642
rect 120172 371204 120224 371210
rect 120172 371146 120224 371152
rect 120172 369980 120224 369986
rect 120172 369922 120224 369928
rect 120184 367062 120212 369922
rect 120172 367056 120224 367062
rect 120172 366998 120224 367004
rect 120828 365702 120856 396782
rect 121368 386368 121420 386374
rect 121368 386310 121420 386316
rect 120816 365696 120868 365702
rect 120816 365638 120868 365644
rect 120724 365016 120776 365022
rect 120724 364958 120776 364964
rect 120736 364410 120764 364958
rect 120724 364404 120776 364410
rect 120724 364346 120776 364352
rect 120080 335164 120132 335170
rect 120080 335106 120132 335112
rect 120080 293072 120132 293078
rect 120080 293014 120132 293020
rect 119988 259344 120040 259350
rect 119988 259286 120040 259292
rect 69018 253192 69074 253201
rect 69018 253127 69074 253136
rect 69032 252618 69060 253127
rect 69020 252612 69072 252618
rect 69020 252554 69072 252560
rect 69032 213246 69060 252554
rect 69110 251288 69166 251297
rect 69110 251223 69166 251232
rect 69124 232626 69152 251223
rect 120092 251025 120120 293014
rect 120736 287054 120764 364346
rect 121276 305720 121328 305726
rect 121276 305662 121328 305668
rect 120736 287026 120948 287054
rect 120920 284374 120948 287026
rect 120908 284368 120960 284374
rect 120906 284336 120908 284345
rect 120960 284336 120962 284345
rect 120906 284271 120962 284280
rect 121288 257145 121316 305662
rect 121274 257136 121330 257145
rect 121274 257071 121276 257080
rect 121328 257071 121330 257080
rect 121276 257042 121328 257048
rect 121288 257011 121316 257042
rect 120078 251016 120134 251025
rect 120078 250951 120134 250960
rect 120092 249898 120120 250951
rect 120080 249892 120132 249898
rect 120080 249834 120132 249840
rect 69202 245032 69258 245041
rect 69202 244967 69258 244976
rect 69216 237386 69244 244967
rect 69846 242312 69902 242321
rect 69846 242247 69902 242256
rect 69860 240106 69888 242247
rect 69848 240100 69900 240106
rect 69848 240042 69900 240048
rect 69952 240094 70058 240122
rect 119646 240094 119752 240122
rect 69952 238202 69980 240094
rect 69940 238196 69992 238202
rect 69940 238138 69992 238144
rect 70688 238134 70716 240037
rect 71320 239850 71348 240037
rect 71240 239822 71348 239850
rect 70676 238128 70728 238134
rect 70676 238070 70728 238076
rect 69204 237380 69256 237386
rect 69204 237322 69256 237328
rect 69112 232620 69164 232626
rect 69112 232562 69164 232568
rect 71240 219434 71268 239822
rect 71976 238754 72004 240037
rect 70412 219406 71268 219434
rect 71792 238726 72004 238754
rect 70412 216073 70440 219406
rect 70398 216064 70454 216073
rect 70398 215999 70454 216008
rect 69020 213240 69072 213246
rect 69020 213182 69072 213188
rect 68926 199336 68982 199345
rect 68926 199271 68982 199280
rect 66076 191276 66128 191282
rect 66076 191218 66128 191224
rect 71792 188426 71820 238726
rect 72620 238610 72648 240037
rect 73252 239850 73280 240037
rect 73896 239850 73924 240037
rect 73172 239822 73280 239850
rect 73816 239822 73924 239850
rect 72608 238604 72660 238610
rect 72608 238546 72660 238552
rect 72620 238066 72648 238546
rect 72608 238060 72660 238066
rect 72608 238002 72660 238008
rect 71780 188420 71832 188426
rect 71780 188362 71832 188368
rect 73172 186998 73200 239822
rect 73816 219434 73844 239822
rect 74552 239442 74580 240037
rect 74552 239414 74764 239442
rect 74632 239352 74684 239358
rect 74632 239294 74684 239300
rect 74448 231872 74500 231878
rect 74500 231826 74580 231854
rect 74448 231814 74500 231820
rect 73264 219406 73844 219434
rect 73264 189854 73292 219406
rect 73252 189848 73304 189854
rect 73252 189790 73304 189796
rect 73160 186992 73212 186998
rect 73160 186934 73212 186940
rect 74552 185609 74580 231826
rect 74644 217462 74672 239294
rect 74736 225622 74764 239414
rect 75196 231878 75224 240037
rect 75840 239358 75868 240037
rect 75920 239828 75972 239834
rect 75920 239770 75972 239776
rect 75828 239352 75880 239358
rect 75828 239294 75880 239300
rect 75184 231872 75236 231878
rect 75184 231814 75236 231820
rect 74724 225616 74776 225622
rect 74724 225558 74776 225564
rect 74632 217456 74684 217462
rect 74632 217398 74684 217404
rect 74538 185600 74594 185609
rect 74538 185535 74594 185544
rect 75932 184278 75960 239770
rect 76484 238754 76512 240037
rect 77116 239834 77144 240037
rect 77104 239828 77156 239834
rect 77104 239770 77156 239776
rect 77300 239828 77352 239834
rect 77300 239770 77352 239776
rect 76484 238726 76604 238754
rect 76576 237289 76604 238726
rect 76562 237280 76618 237289
rect 76562 237215 76618 237224
rect 76576 220153 76604 237215
rect 76562 220144 76618 220153
rect 76562 220079 76618 220088
rect 77312 189922 77340 239770
rect 77772 238754 77800 240037
rect 78404 239834 78432 240037
rect 78392 239828 78444 239834
rect 78392 239770 78444 239776
rect 78312 239488 78364 239494
rect 78312 239430 78364 239436
rect 77404 238726 77800 238754
rect 77404 209001 77432 238726
rect 78324 232694 78352 239430
rect 79060 238754 79088 240037
rect 79692 239850 79720 240037
rect 78692 238726 79088 238754
rect 79612 239822 79720 239850
rect 80060 239828 80112 239834
rect 78312 232688 78364 232694
rect 78312 232630 78364 232636
rect 77390 208992 77446 209001
rect 77390 208927 77446 208936
rect 77300 189916 77352 189922
rect 77300 189858 77352 189864
rect 75920 184272 75972 184278
rect 75920 184214 75972 184220
rect 64696 182912 64748 182918
rect 78692 182889 78720 238726
rect 79612 219434 79640 239822
rect 80060 239770 80112 239776
rect 78784 219406 79640 219434
rect 78784 206310 78812 219406
rect 78772 206304 78824 206310
rect 78772 206246 78824 206252
rect 80072 185706 80100 239770
rect 80348 238754 80376 240037
rect 80980 239834 81008 240037
rect 80968 239828 81020 239834
rect 80968 239770 81020 239776
rect 80164 238726 80376 238754
rect 80164 202162 80192 238726
rect 81636 237318 81664 240037
rect 82280 238754 82308 240037
rect 82912 239850 82940 240037
rect 83556 239850 83584 240037
rect 82004 238726 82308 238754
rect 82832 239822 82940 239850
rect 83476 239822 83584 239850
rect 81624 237312 81676 237318
rect 81624 237254 81676 237260
rect 81636 236026 81664 237254
rect 81624 236020 81676 236026
rect 81624 235962 81676 235968
rect 82004 219434 82032 238726
rect 82084 236020 82136 236026
rect 82084 235962 82136 235968
rect 81544 219406 82032 219434
rect 81544 215286 81572 219406
rect 81532 215280 81584 215286
rect 81532 215222 81584 215228
rect 80152 202156 80204 202162
rect 80152 202098 80204 202104
rect 82096 199442 82124 235962
rect 82832 205630 82860 239822
rect 83476 230450 83504 239822
rect 84212 233850 84240 240037
rect 84856 238754 84884 240037
rect 84304 238726 84884 238754
rect 84200 233844 84252 233850
rect 84200 233786 84252 233792
rect 84304 233730 84332 238726
rect 85500 237454 85528 240037
rect 86144 238678 86172 240037
rect 86788 238746 86816 240037
rect 86960 239828 87012 239834
rect 86960 239770 87012 239776
rect 86776 238740 86828 238746
rect 86776 238682 86828 238688
rect 86132 238672 86184 238678
rect 86132 238614 86184 238620
rect 86144 237969 86172 238614
rect 86788 238338 86816 238682
rect 86776 238332 86828 238338
rect 86776 238274 86828 238280
rect 86316 238060 86368 238066
rect 86316 238002 86368 238008
rect 86130 237960 86186 237969
rect 86130 237895 86186 237904
rect 85488 237448 85540 237454
rect 85488 237390 85540 237396
rect 86224 237448 86276 237454
rect 86224 237390 86276 237396
rect 84212 233702 84332 233730
rect 82912 230444 82964 230450
rect 82912 230386 82964 230392
rect 83464 230444 83516 230450
rect 83464 230386 83516 230392
rect 82924 222698 82952 230386
rect 82912 222692 82964 222698
rect 82912 222634 82964 222640
rect 83464 222692 83516 222698
rect 83464 222634 83516 222640
rect 82924 222222 82952 222634
rect 82912 222216 82964 222222
rect 82912 222158 82964 222164
rect 82820 205624 82872 205630
rect 82820 205566 82872 205572
rect 82084 199436 82136 199442
rect 82084 199378 82136 199384
rect 83476 196654 83504 222634
rect 83464 196648 83516 196654
rect 83464 196590 83516 196596
rect 84212 185842 84240 233702
rect 84292 233640 84344 233646
rect 84292 233582 84344 233588
rect 84304 192545 84332 233582
rect 86236 202230 86264 237390
rect 86328 221474 86356 238002
rect 86316 221468 86368 221474
rect 86316 221410 86368 221416
rect 86972 203794 87000 239770
rect 87432 238754 87460 240037
rect 88064 239834 88092 240037
rect 88052 239828 88104 239834
rect 88052 239770 88104 239776
rect 88248 239420 88300 239426
rect 88248 239362 88300 239368
rect 87064 238726 87460 238754
rect 88260 238746 88288 239362
rect 88720 238754 88748 240037
rect 89352 239850 89380 240037
rect 88248 238740 88300 238746
rect 87064 215937 87092 238726
rect 88248 238682 88300 238688
rect 88352 238726 88748 238754
rect 89272 239822 89380 239850
rect 89720 239828 89772 239834
rect 87050 215928 87106 215937
rect 87050 215863 87106 215872
rect 86960 203788 87012 203794
rect 86960 203730 87012 203736
rect 86224 202224 86276 202230
rect 86224 202166 86276 202172
rect 84290 192536 84346 192545
rect 84290 192471 84346 192480
rect 88352 191146 88380 238726
rect 89272 230382 89300 239822
rect 89720 239770 89772 239776
rect 89260 230376 89312 230382
rect 89260 230318 89312 230324
rect 89732 194206 89760 239770
rect 90008 238754 90036 240037
rect 90640 239834 90668 240037
rect 90628 239828 90680 239834
rect 90628 239770 90680 239776
rect 89824 238726 90036 238754
rect 89824 218822 89852 238726
rect 91296 234433 91324 240037
rect 91940 238754 91968 240037
rect 92572 239850 92600 240037
rect 93216 239850 93244 240037
rect 91756 238726 91968 238754
rect 92492 239822 92600 239850
rect 93136 239822 93244 239850
rect 91756 234530 91784 238726
rect 91744 234524 91796 234530
rect 91744 234466 91796 234472
rect 91282 234424 91338 234433
rect 91282 234359 91338 234368
rect 91756 224942 91784 234466
rect 91744 224936 91796 224942
rect 91744 224878 91796 224884
rect 89812 218816 89864 218822
rect 89812 218758 89864 218764
rect 92492 195498 92520 239822
rect 93136 219434 93164 239822
rect 93872 239442 93900 240037
rect 93872 239414 94084 239442
rect 93952 239352 94004 239358
rect 93952 239294 94004 239300
rect 93768 231872 93820 231878
rect 93820 231826 93900 231854
rect 93768 231814 93820 231820
rect 92584 219406 93164 219434
rect 92584 205018 92612 219406
rect 92572 205012 92624 205018
rect 92572 204954 92624 204960
rect 92480 195492 92532 195498
rect 92480 195434 92532 195440
rect 89720 194200 89772 194206
rect 89720 194142 89772 194148
rect 93872 194070 93900 231826
rect 93964 198082 93992 239294
rect 94056 227050 94084 239414
rect 94516 231878 94544 240037
rect 95160 239358 95188 240037
rect 95240 239828 95292 239834
rect 95240 239770 95292 239776
rect 95148 239352 95200 239358
rect 95148 239294 95200 239300
rect 94504 231872 94556 231878
rect 94504 231814 94556 231820
rect 94044 227044 94096 227050
rect 94044 226986 94096 226992
rect 93952 198076 94004 198082
rect 93952 198018 94004 198024
rect 93860 194064 93912 194070
rect 93860 194006 93912 194012
rect 88340 191140 88392 191146
rect 88340 191082 88392 191088
rect 95252 187066 95280 239770
rect 95804 235793 95832 240037
rect 96436 239834 96464 240037
rect 96424 239828 96476 239834
rect 96424 239770 96476 239776
rect 96620 239828 96672 239834
rect 96620 239770 96672 239776
rect 95790 235784 95846 235793
rect 95790 235719 95846 235728
rect 95240 187060 95292 187066
rect 95240 187002 95292 187008
rect 84200 185836 84252 185842
rect 84200 185778 84252 185784
rect 80060 185700 80112 185706
rect 80060 185642 80112 185648
rect 64696 182854 64748 182860
rect 78678 182880 78734 182889
rect 78678 182815 78734 182824
rect 96632 181558 96660 239770
rect 97092 238754 97120 240037
rect 97724 239834 97752 240037
rect 97712 239828 97764 239834
rect 97712 239770 97764 239776
rect 96724 238726 97120 238754
rect 96724 201074 96752 238726
rect 98380 238649 98408 240037
rect 99024 238754 99052 240037
rect 99668 238754 99696 240037
rect 99024 238726 99328 238754
rect 98366 238640 98422 238649
rect 98366 238575 98422 238584
rect 98828 238332 98880 238338
rect 98828 238274 98880 238280
rect 98840 238066 98868 238274
rect 98828 238060 98880 238066
rect 98828 238002 98880 238008
rect 99196 238060 99248 238066
rect 99196 238002 99248 238008
rect 98642 235784 98698 235793
rect 98642 235719 98698 235728
rect 98656 228410 98684 235719
rect 98644 228404 98696 228410
rect 98644 228346 98696 228352
rect 96712 201068 96764 201074
rect 96712 201010 96764 201016
rect 99208 200802 99236 238002
rect 99300 237318 99328 238726
rect 99392 238726 99696 238754
rect 99288 237312 99340 237318
rect 99288 237254 99340 237260
rect 99196 200796 99248 200802
rect 99196 200738 99248 200744
rect 99300 193934 99328 237254
rect 99288 193928 99340 193934
rect 99288 193870 99340 193876
rect 99392 188562 99420 238726
rect 100312 238270 100340 240037
rect 100956 238754 100984 240037
rect 101588 239850 101616 240037
rect 102232 239850 102260 240037
rect 100772 238726 100984 238754
rect 101508 239822 101616 239850
rect 102152 239822 102260 239850
rect 100300 238264 100352 238270
rect 100300 238206 100352 238212
rect 100772 206378 100800 238726
rect 101508 231198 101536 239822
rect 101496 231192 101548 231198
rect 101496 231134 101548 231140
rect 100760 206372 100812 206378
rect 100760 206314 100812 206320
rect 102152 191350 102180 239822
rect 102888 237454 102916 240037
rect 103532 238746 103560 240037
rect 104176 239442 104204 240037
rect 104808 239850 104836 240037
rect 103992 239414 104204 239442
rect 104728 239822 104836 239850
rect 104900 239828 104952 239834
rect 103992 238754 104020 239414
rect 104728 238754 104756 239822
rect 104900 239770 104952 239776
rect 103520 238740 103572 238746
rect 103520 238682 103572 238688
rect 103624 238726 104020 238754
rect 104084 238726 104756 238754
rect 103532 237522 103560 238682
rect 103520 237516 103572 237522
rect 103520 237458 103572 237464
rect 102876 237448 102928 237454
rect 102876 237390 102928 237396
rect 103624 222873 103652 238726
rect 103610 222864 103666 222873
rect 103610 222799 103666 222808
rect 104084 219434 104112 238726
rect 104164 237516 104216 237522
rect 104164 237458 104216 237464
rect 103716 219406 104112 219434
rect 102140 191344 102192 191350
rect 102140 191286 102192 191292
rect 99380 188556 99432 188562
rect 99380 188498 99432 188504
rect 103428 187808 103480 187814
rect 103428 187750 103480 187756
rect 100668 184952 100720 184958
rect 100668 184894 100720 184900
rect 96620 181552 96672 181558
rect 96620 181494 96672 181500
rect 97356 179512 97408 179518
rect 97356 179454 97408 179460
rect 64512 178764 64564 178770
rect 64512 178706 64564 178712
rect 97368 177041 97396 179454
rect 97354 177032 97410 177041
rect 97354 176967 97410 176976
rect 100680 176769 100708 184894
rect 103440 176769 103468 187750
rect 103716 184414 103744 219406
rect 104176 217326 104204 237458
rect 104164 217320 104216 217326
rect 104164 217262 104216 217268
rect 104912 201006 104940 239770
rect 105464 238338 105492 240037
rect 106096 239834 106124 240037
rect 106084 239828 106136 239834
rect 106084 239770 106136 239776
rect 106752 238754 106780 240037
rect 106292 238726 106780 238754
rect 105452 238332 105504 238338
rect 105452 238274 105504 238280
rect 105544 237448 105596 237454
rect 105544 237390 105596 237396
rect 104900 201000 104952 201006
rect 104900 200942 104952 200948
rect 105556 196790 105584 237390
rect 106292 212537 106320 238726
rect 107396 235929 107424 240037
rect 107382 235920 107438 235929
rect 107382 235855 107438 235864
rect 107396 232558 107424 235855
rect 108040 233918 108068 240037
rect 108672 239850 108700 240037
rect 109960 239850 109988 240037
rect 108592 239822 108700 239850
rect 109880 239822 109988 239850
rect 108028 233912 108080 233918
rect 108028 233854 108080 233860
rect 107384 232552 107436 232558
rect 107384 232494 107436 232500
rect 108592 219434 108620 239822
rect 109880 238754 109908 239822
rect 109696 238726 109908 238754
rect 109696 233238 109724 238726
rect 110616 235958 110644 240037
rect 111260 238754 111288 240037
rect 111892 239850 111920 240037
rect 110892 238726 111288 238754
rect 111812 239822 111920 239850
rect 110604 235952 110656 235958
rect 110604 235894 110656 235900
rect 109684 233232 109736 233238
rect 109684 233174 109736 233180
rect 107672 219406 108620 219434
rect 106278 212528 106334 212537
rect 106278 212463 106334 212472
rect 105544 196784 105596 196790
rect 105544 196726 105596 196732
rect 106188 189236 106240 189242
rect 106188 189178 106240 189184
rect 104808 189168 104860 189174
rect 104808 189110 104860 189116
rect 103704 184408 103756 184414
rect 103704 184350 103756 184356
rect 104820 177721 104848 189110
rect 106200 177721 106228 189178
rect 107672 182850 107700 219406
rect 109696 209846 109724 233174
rect 110892 219434 110920 238726
rect 111064 235952 111116 235958
rect 111064 235894 111116 235900
rect 110432 219406 110920 219434
rect 109684 209840 109736 209846
rect 109684 209782 109736 209788
rect 108948 190528 109000 190534
rect 108948 190470 109000 190476
rect 107660 182844 107712 182850
rect 107660 182786 107712 182792
rect 108960 177721 108988 190470
rect 104806 177712 104862 177721
rect 104806 177647 104862 177656
rect 106186 177712 106242 177721
rect 106186 177647 106242 177656
rect 108946 177712 109002 177721
rect 108946 177647 109002 177656
rect 109408 176792 109460 176798
rect 100666 176760 100722 176769
rect 100666 176695 100722 176704
rect 102046 176760 102102 176769
rect 102046 176695 102048 176704
rect 102100 176695 102102 176704
rect 103426 176760 103482 176769
rect 109408 176734 109460 176740
rect 103426 176695 103482 176704
rect 102048 176666 102100 176672
rect 98368 175976 98420 175982
rect 109420 175953 109448 176734
rect 109696 176050 109724 209782
rect 110432 196858 110460 219406
rect 110420 196852 110472 196858
rect 110420 196794 110472 196800
rect 109776 178220 109828 178226
rect 109776 178162 109828 178168
rect 109788 176769 109816 178162
rect 111076 176866 111104 235894
rect 111812 207738 111840 239822
rect 112548 238814 112576 240037
rect 111892 238808 111944 238814
rect 111892 238750 111944 238756
rect 112536 238808 112588 238814
rect 112536 238750 112588 238756
rect 111904 228478 111932 238750
rect 111892 228472 111944 228478
rect 111892 228414 111944 228420
rect 113192 209166 113220 240037
rect 113836 237289 113864 240037
rect 114480 238746 114508 240037
rect 114560 239828 114612 239834
rect 114560 239770 114612 239776
rect 114468 238740 114520 238746
rect 114468 238682 114520 238688
rect 113822 237280 113878 237289
rect 113822 237215 113878 237224
rect 113836 236065 113864 237215
rect 113822 236056 113878 236065
rect 113822 235991 113878 236000
rect 114466 236056 114522 236065
rect 114466 235991 114522 236000
rect 113180 209160 113232 209166
rect 113180 209102 113232 209108
rect 111800 207732 111852 207738
rect 111800 207674 111852 207680
rect 114480 203862 114508 235991
rect 114468 203856 114520 203862
rect 114468 203798 114520 203804
rect 114572 203726 114600 239770
rect 115124 238754 115152 240037
rect 115756 239834 115784 240037
rect 115744 239828 115796 239834
rect 115744 239770 115796 239776
rect 116412 239442 116440 240037
rect 114664 238726 115152 238754
rect 115952 239414 116440 239442
rect 114664 219337 114692 238726
rect 114650 219328 114706 219337
rect 114650 219263 114706 219272
rect 114560 203720 114612 203726
rect 114560 203662 114612 203668
rect 115952 182986 115980 239414
rect 117056 238814 117084 240037
rect 117700 239970 117728 240037
rect 117688 239964 117740 239970
rect 117688 239906 117740 239912
rect 118332 239850 118360 240037
rect 118252 239822 118360 239850
rect 116032 238808 116084 238814
rect 116032 238750 116084 238756
rect 117044 238808 117096 238814
rect 117044 238750 117096 238756
rect 116044 199510 116072 238750
rect 118252 222154 118280 239822
rect 118988 234598 119016 240037
rect 119724 238754 119752 240094
rect 119080 238726 119752 238754
rect 118976 234592 119028 234598
rect 118976 234534 119028 234540
rect 118988 234190 119016 234534
rect 118976 234184 119028 234190
rect 118976 234126 119028 234132
rect 118240 222148 118292 222154
rect 118240 222090 118292 222096
rect 119080 219434 119108 238726
rect 119344 234184 119396 234190
rect 119344 234126 119396 234132
rect 118712 219406 119108 219434
rect 116032 199504 116084 199510
rect 116032 199446 116084 199452
rect 118712 188494 118740 219406
rect 119356 206281 119384 234126
rect 119342 206272 119398 206281
rect 119342 206207 119398 206216
rect 120092 203590 120120 249834
rect 121380 247625 121408 386310
rect 121472 367878 121500 475322
rect 121564 388385 121592 492322
rect 121656 460934 121684 494906
rect 121656 460906 121776 460934
rect 121642 439512 121698 439521
rect 121642 439447 121698 439456
rect 121656 439006 121684 439447
rect 121644 439000 121696 439006
rect 121644 438942 121696 438948
rect 121748 438870 121776 460906
rect 122116 439521 122144 538222
rect 122852 490521 122880 585414
rect 122932 582548 122984 582554
rect 122932 582490 122984 582496
rect 122944 491570 122972 582490
rect 123116 576156 123168 576162
rect 123116 576098 123168 576104
rect 123128 576065 123156 576098
rect 123114 576056 123170 576065
rect 123114 575991 123170 576000
rect 123128 575550 123156 575991
rect 123116 575544 123168 575550
rect 123116 575486 123168 575492
rect 123024 537668 123076 537674
rect 123024 537610 123076 537616
rect 122932 491564 122984 491570
rect 122932 491506 122984 491512
rect 122838 490512 122894 490521
rect 122838 490447 122894 490456
rect 122944 488578 122972 491506
rect 122932 488572 122984 488578
rect 122932 488514 122984 488520
rect 122932 487892 122984 487898
rect 122932 487834 122984 487840
rect 122840 449948 122892 449954
rect 122840 449890 122892 449896
rect 122102 439512 122158 439521
rect 122102 439447 122158 439456
rect 121736 438864 121788 438870
rect 121736 438806 121788 438812
rect 121644 404388 121696 404394
rect 121644 404330 121696 404336
rect 121656 397458 121684 404330
rect 121644 397452 121696 397458
rect 121644 397394 121696 397400
rect 121550 388376 121606 388385
rect 121550 388311 121606 388320
rect 121564 386374 121592 388311
rect 122196 388136 122248 388142
rect 122196 388078 122248 388084
rect 121552 386368 121604 386374
rect 121552 386310 121604 386316
rect 122104 385348 122156 385354
rect 122104 385290 122156 385296
rect 121552 378208 121604 378214
rect 121552 378150 121604 378156
rect 121564 377602 121592 378150
rect 121552 377596 121604 377602
rect 121552 377538 121604 377544
rect 121460 367872 121512 367878
rect 121460 367814 121512 367820
rect 121460 365696 121512 365702
rect 121460 365638 121512 365644
rect 121472 364410 121500 365638
rect 121460 364404 121512 364410
rect 121460 364346 121512 364352
rect 121472 339454 121500 364346
rect 121460 339448 121512 339454
rect 121460 339390 121512 339396
rect 122012 329792 122064 329798
rect 122010 329760 122012 329769
rect 122064 329760 122066 329769
rect 122010 329695 122066 329704
rect 121460 329180 121512 329186
rect 121460 329122 121512 329128
rect 121472 286686 121500 329122
rect 122024 328506 122052 329695
rect 122012 328500 122064 328506
rect 122012 328442 122064 328448
rect 122116 326398 122144 385290
rect 122208 349858 122236 388078
rect 122288 385688 122340 385694
rect 122288 385630 122340 385636
rect 122300 385354 122328 385630
rect 122288 385348 122340 385354
rect 122288 385290 122340 385296
rect 122196 349852 122248 349858
rect 122196 349794 122248 349800
rect 122852 336598 122880 449890
rect 122944 384402 122972 487834
rect 123036 438802 123064 537610
rect 124232 532030 124260 589290
rect 125600 586696 125652 586702
rect 125600 586638 125652 586644
rect 124864 568608 124916 568614
rect 124864 568550 124916 568556
rect 124404 534744 124456 534750
rect 124404 534686 124456 534692
rect 124220 532024 124272 532030
rect 124220 531966 124272 531972
rect 124312 500268 124364 500274
rect 124312 500210 124364 500216
rect 123116 494080 123168 494086
rect 123116 494022 123168 494028
rect 123128 443698 123156 494022
rect 123206 483712 123262 483721
rect 123206 483647 123208 483656
rect 123260 483647 123262 483656
rect 123208 483618 123260 483624
rect 123116 443692 123168 443698
rect 123116 443634 123168 443640
rect 124220 438864 124272 438870
rect 124220 438806 124272 438812
rect 123024 438796 123076 438802
rect 123024 438738 123076 438744
rect 123024 392692 123076 392698
rect 123024 392634 123076 392640
rect 122932 384396 122984 384402
rect 122932 384338 122984 384344
rect 122932 367260 122984 367266
rect 122932 367202 122984 367208
rect 122840 336592 122892 336598
rect 122840 336534 122892 336540
rect 122196 326528 122248 326534
rect 122196 326470 122248 326476
rect 122104 326392 122156 326398
rect 122104 326334 122156 326340
rect 121552 308508 121604 308514
rect 121552 308450 121604 308456
rect 121564 306374 121592 308450
rect 121564 306346 121776 306374
rect 121552 291848 121604 291854
rect 121550 291816 121552 291825
rect 121604 291816 121606 291825
rect 121550 291751 121606 291760
rect 121642 291136 121698 291145
rect 121642 291071 121698 291080
rect 121550 290456 121606 290465
rect 121550 290391 121606 290400
rect 121564 289950 121592 290391
rect 121552 289944 121604 289950
rect 121552 289886 121604 289892
rect 121656 289882 121684 291071
rect 121644 289876 121696 289882
rect 121644 289818 121696 289824
rect 121748 289785 121776 306346
rect 121826 296032 121882 296041
rect 121826 295967 121882 295976
rect 121734 289776 121790 289785
rect 121734 289711 121790 289720
rect 121748 289202 121776 289711
rect 121736 289196 121788 289202
rect 121736 289138 121788 289144
rect 121840 289134 121868 295967
rect 121828 289128 121880 289134
rect 121642 289096 121698 289105
rect 121828 289070 121880 289076
rect 122012 289128 122064 289134
rect 122012 289070 122064 289076
rect 121642 289031 121698 289040
rect 121656 288454 121684 289031
rect 121644 288448 121696 288454
rect 121644 288390 121696 288396
rect 121552 288380 121604 288386
rect 121552 288322 121604 288328
rect 121564 287745 121592 288322
rect 121550 287736 121606 287745
rect 121550 287671 121606 287680
rect 121550 287056 121606 287065
rect 122024 287054 122052 289070
rect 122024 287026 122144 287054
rect 121550 286991 121606 287000
rect 121460 286680 121512 286686
rect 121460 286622 121512 286628
rect 121460 286544 121512 286550
rect 121460 286486 121512 286492
rect 121472 285705 121500 286486
rect 121564 286482 121592 286991
rect 121644 286680 121696 286686
rect 121644 286622 121696 286628
rect 121552 286476 121604 286482
rect 121552 286418 121604 286424
rect 121656 286414 121684 286622
rect 121644 286408 121696 286414
rect 121642 286376 121644 286385
rect 121696 286376 121698 286385
rect 121642 286311 121698 286320
rect 121656 286285 121684 286311
rect 121458 285696 121514 285705
rect 121458 285631 121514 285640
rect 121458 285016 121514 285025
rect 121458 284951 121514 284960
rect 121472 284442 121500 284951
rect 121460 284436 121512 284442
rect 121460 284378 121512 284384
rect 121458 282976 121514 282985
rect 121458 282911 121460 282920
rect 121512 282911 121514 282920
rect 121460 282882 121512 282888
rect 121458 281616 121514 281625
rect 121458 281551 121460 281560
rect 121512 281551 121514 281560
rect 121460 281522 121512 281528
rect 121458 280256 121514 280265
rect 121458 280191 121460 280200
rect 121512 280191 121514 280200
rect 121460 280162 121512 280168
rect 121550 279576 121606 279585
rect 121550 279511 121606 279520
rect 121458 278896 121514 278905
rect 121564 278866 121592 279511
rect 121458 278831 121514 278840
rect 121552 278860 121604 278866
rect 121472 278798 121500 278831
rect 121552 278802 121604 278808
rect 121460 278792 121512 278798
rect 121460 278734 121512 278740
rect 121550 278216 121606 278225
rect 121550 278151 121606 278160
rect 121458 277536 121514 277545
rect 121458 277471 121460 277480
rect 121512 277471 121514 277480
rect 121460 277442 121512 277448
rect 121564 277438 121592 278151
rect 121552 277432 121604 277438
rect 121552 277374 121604 277380
rect 121642 276312 121698 276321
rect 121642 276247 121698 276256
rect 121458 276176 121514 276185
rect 121458 276111 121460 276120
rect 121512 276111 121514 276120
rect 121460 276082 121512 276088
rect 121552 276072 121604 276078
rect 121552 276014 121604 276020
rect 121564 275505 121592 276014
rect 121550 275496 121606 275505
rect 121550 275431 121606 275440
rect 121458 274816 121514 274825
rect 121458 274751 121514 274760
rect 121472 274718 121500 274751
rect 121460 274712 121512 274718
rect 121460 274654 121512 274660
rect 121458 273456 121514 273465
rect 121458 273391 121514 273400
rect 121472 273290 121500 273391
rect 121460 273284 121512 273290
rect 121460 273226 121512 273232
rect 121458 272776 121514 272785
rect 121458 272711 121514 272720
rect 121472 272542 121500 272711
rect 121460 272536 121512 272542
rect 121460 272478 121512 272484
rect 121458 272096 121514 272105
rect 121458 272031 121514 272040
rect 121472 271930 121500 272031
rect 121460 271924 121512 271930
rect 121460 271866 121512 271872
rect 121458 271416 121514 271425
rect 121458 271351 121514 271360
rect 121472 270570 121500 271351
rect 121460 270564 121512 270570
rect 121460 270506 121512 270512
rect 121458 270056 121514 270065
rect 121458 269991 121514 270000
rect 121472 269210 121500 269991
rect 121550 269376 121606 269385
rect 121550 269311 121606 269320
rect 121460 269204 121512 269210
rect 121460 269146 121512 269152
rect 121564 269142 121592 269311
rect 121552 269136 121604 269142
rect 121552 269078 121604 269084
rect 121460 269068 121512 269074
rect 121460 269010 121512 269016
rect 121472 268705 121500 269010
rect 121458 268696 121514 268705
rect 121458 268631 121514 268640
rect 121656 268546 121684 276247
rect 121918 276040 121974 276049
rect 121918 275975 121974 275984
rect 121932 272513 121960 275975
rect 122116 274145 122144 287026
rect 122208 277394 122236 326470
rect 122944 294302 122972 367202
rect 123036 338026 123064 392634
rect 123114 378992 123170 379001
rect 123114 378927 123170 378936
rect 123128 378894 123156 378927
rect 123116 378888 123168 378894
rect 123116 378830 123168 378836
rect 123024 338020 123076 338026
rect 123024 337962 123076 337968
rect 122932 294296 122984 294302
rect 122932 294238 122984 294244
rect 122286 288416 122342 288425
rect 122286 288351 122342 288360
rect 122300 286346 122328 288351
rect 122288 286340 122340 286346
rect 122288 286282 122340 286288
rect 122208 277366 122328 277394
rect 122300 276078 122328 277366
rect 122288 276072 122340 276078
rect 122288 276014 122340 276020
rect 122102 274136 122158 274145
rect 122102 274071 122158 274080
rect 121918 272504 121974 272513
rect 121918 272439 121974 272448
rect 121472 268518 121684 268546
rect 121472 257922 121500 268518
rect 121550 268016 121606 268025
rect 121550 267951 121606 267960
rect 121564 267782 121592 267951
rect 121552 267776 121604 267782
rect 121552 267718 121604 267724
rect 121642 267336 121698 267345
rect 121642 267271 121698 267280
rect 121550 266656 121606 266665
rect 121550 266591 121606 266600
rect 121564 266422 121592 266591
rect 121656 266490 121684 267271
rect 121644 266484 121696 266490
rect 121644 266426 121696 266432
rect 121552 266416 121604 266422
rect 121552 266358 121604 266364
rect 121642 265976 121698 265985
rect 121642 265911 121698 265920
rect 121550 265296 121606 265305
rect 121550 265231 121606 265240
rect 121564 265062 121592 265231
rect 121552 265056 121604 265062
rect 121552 264998 121604 265004
rect 121656 264994 121684 265911
rect 121644 264988 121696 264994
rect 121644 264930 121696 264936
rect 121642 263936 121698 263945
rect 121642 263871 121698 263880
rect 121656 263634 121684 263871
rect 121644 263628 121696 263634
rect 121644 263570 121696 263576
rect 123036 263566 123064 337962
rect 123128 337550 123156 378830
rect 124128 367804 124180 367810
rect 124128 367746 124180 367752
rect 124140 367266 124168 367746
rect 124128 367260 124180 367266
rect 124128 367202 124180 367208
rect 123116 337544 123168 337550
rect 123116 337486 123168 337492
rect 124232 336598 124260 438806
rect 124324 436082 124352 500210
rect 124416 437442 124444 534686
rect 124876 478922 124904 568550
rect 124956 528624 125008 528630
rect 124956 528566 125008 528572
rect 124864 478916 124916 478922
rect 124864 478858 124916 478864
rect 124876 477426 124904 478858
rect 124864 477420 124916 477426
rect 124864 477362 124916 477368
rect 124968 459610 124996 528566
rect 125612 490618 125640 586638
rect 128360 583840 128412 583846
rect 128360 583782 128412 583788
rect 126980 579760 127032 579766
rect 126980 579702 127032 579708
rect 126888 574048 126940 574054
rect 126888 573990 126940 573996
rect 126900 573374 126928 573990
rect 126152 573368 126204 573374
rect 126152 573310 126204 573316
rect 126888 573368 126940 573374
rect 126888 573310 126940 573316
rect 126164 572801 126192 573310
rect 126150 572792 126206 572801
rect 126150 572727 126206 572736
rect 125968 555484 126020 555490
rect 125968 555426 126020 555432
rect 125784 534812 125836 534818
rect 125784 534754 125836 534760
rect 125600 490612 125652 490618
rect 125600 490554 125652 490560
rect 125690 484392 125746 484401
rect 125690 484327 125746 484336
rect 125704 483070 125732 484327
rect 125692 483064 125744 483070
rect 125692 483006 125744 483012
rect 125508 467152 125560 467158
rect 125508 467094 125560 467100
rect 125520 466478 125548 467094
rect 125508 466472 125560 466478
rect 125508 466414 125560 466420
rect 124956 459604 125008 459610
rect 124956 459546 125008 459552
rect 124404 437436 124456 437442
rect 124404 437378 124456 437384
rect 124312 436076 124364 436082
rect 124312 436018 124364 436024
rect 124312 393984 124364 393990
rect 124312 393926 124364 393932
rect 123484 336592 123536 336598
rect 123484 336534 123536 336540
rect 124220 336592 124272 336598
rect 124220 336534 124272 336540
rect 123496 336054 123524 336534
rect 123484 336048 123536 336054
rect 123484 335990 123536 335996
rect 123496 272542 123524 335990
rect 124220 331900 124272 331906
rect 124220 331842 124272 331848
rect 123668 294296 123720 294302
rect 123668 294238 123720 294244
rect 123576 274780 123628 274786
rect 123576 274722 123628 274728
rect 123484 272536 123536 272542
rect 123484 272478 123536 272484
rect 121552 263560 121604 263566
rect 121552 263502 121604 263508
rect 123024 263560 123076 263566
rect 123024 263502 123076 263508
rect 121564 263265 121592 263502
rect 121550 263256 121606 263265
rect 121550 263191 121606 263200
rect 121550 262576 121606 262585
rect 121550 262511 121606 262520
rect 121564 262342 121592 262511
rect 121552 262336 121604 262342
rect 121552 262278 121604 262284
rect 121552 262200 121604 262206
rect 121552 262142 121604 262148
rect 121564 261225 121592 262142
rect 121642 261896 121698 261905
rect 121642 261831 121698 261840
rect 121550 261216 121606 261225
rect 121550 261151 121606 261160
rect 121656 260914 121684 261831
rect 121644 260908 121696 260914
rect 121644 260850 121696 260856
rect 121552 260840 121604 260846
rect 121552 260782 121604 260788
rect 121564 260545 121592 260782
rect 121550 260536 121606 260545
rect 121550 260471 121606 260480
rect 121550 259856 121606 259865
rect 121550 259791 121606 259800
rect 121564 259554 121592 259791
rect 121552 259548 121604 259554
rect 121552 259490 121604 259496
rect 121552 259412 121604 259418
rect 121552 259354 121604 259360
rect 121564 258505 121592 259354
rect 121644 259344 121696 259350
rect 121644 259286 121696 259292
rect 121550 258496 121606 258505
rect 121550 258431 121606 258440
rect 121460 257916 121512 257922
rect 121460 257858 121512 257864
rect 121458 257816 121514 257825
rect 121458 257751 121514 257760
rect 121472 256766 121500 257751
rect 121656 257258 121684 259286
rect 121734 259176 121790 259185
rect 121734 259111 121790 259120
rect 121748 258126 121776 259111
rect 121736 258120 121788 258126
rect 121736 258062 121788 258068
rect 121736 257916 121788 257922
rect 121736 257858 121788 257864
rect 121564 257230 121684 257258
rect 121460 256760 121512 256766
rect 121460 256702 121512 256708
rect 121458 256456 121514 256465
rect 121458 256391 121514 256400
rect 121472 255270 121500 256391
rect 121460 255264 121512 255270
rect 121460 255206 121512 255212
rect 121458 254416 121514 254425
rect 121458 254351 121514 254360
rect 121472 253978 121500 254351
rect 121460 253972 121512 253978
rect 121460 253914 121512 253920
rect 121458 253056 121514 253065
rect 121458 252991 121514 253000
rect 121472 252618 121500 252991
rect 121460 252612 121512 252618
rect 121460 252554 121512 252560
rect 121458 251696 121514 251705
rect 121458 251631 121514 251640
rect 121472 251258 121500 251631
rect 121460 251252 121512 251258
rect 121460 251194 121512 251200
rect 121458 250336 121514 250345
rect 121458 250271 121514 250280
rect 121472 249830 121500 250271
rect 121460 249824 121512 249830
rect 121460 249766 121512 249772
rect 121458 248976 121514 248985
rect 121458 248911 121514 248920
rect 121472 248470 121500 248911
rect 121460 248464 121512 248470
rect 121460 248406 121512 248412
rect 121564 248414 121592 257230
rect 121644 257100 121696 257106
rect 121644 257042 121696 257048
rect 121656 256018 121684 257042
rect 121644 256012 121696 256018
rect 121644 255954 121696 255960
rect 121642 255096 121698 255105
rect 121642 255031 121698 255040
rect 121656 254046 121684 255031
rect 121644 254040 121696 254046
rect 121644 253982 121696 253988
rect 121642 253736 121698 253745
rect 121642 253671 121698 253680
rect 121656 252686 121684 253671
rect 121644 252680 121696 252686
rect 121644 252622 121696 252628
rect 121748 252385 121776 257858
rect 122840 255808 122892 255814
rect 122746 255776 122802 255785
rect 122802 255756 122840 255762
rect 122802 255750 122892 255756
rect 122802 255734 122880 255750
rect 122746 255711 122802 255720
rect 121734 252376 121790 252385
rect 121734 252311 121790 252320
rect 121748 251870 121776 252311
rect 121736 251864 121788 251870
rect 121736 251806 121788 251812
rect 122840 249892 122892 249898
rect 122840 249834 122892 249840
rect 121642 249656 121698 249665
rect 121642 249591 121698 249600
rect 121656 249422 121684 249591
rect 121644 249416 121696 249422
rect 121644 249358 121696 249364
rect 122748 249416 122800 249422
rect 122748 249358 122800 249364
rect 121564 248386 121684 248414
rect 121458 248296 121514 248305
rect 121458 248231 121514 248240
rect 121366 247616 121422 247625
rect 121366 247551 121422 247560
rect 121380 246922 121408 247551
rect 121472 247110 121500 248231
rect 121460 247104 121512 247110
rect 121460 247046 121512 247052
rect 121550 246936 121606 246945
rect 121380 246894 121500 246922
rect 121472 246362 121500 246894
rect 121550 246871 121606 246880
rect 121460 246356 121512 246362
rect 121460 246298 121512 246304
rect 121458 246256 121514 246265
rect 121458 246191 121514 246200
rect 121472 245682 121500 246191
rect 121564 245750 121592 246871
rect 121552 245744 121604 245750
rect 121552 245686 121604 245692
rect 121460 245676 121512 245682
rect 121460 245618 121512 245624
rect 121550 245576 121606 245585
rect 121550 245511 121606 245520
rect 121458 244896 121514 244905
rect 121458 244831 121514 244840
rect 121472 244254 121500 244831
rect 121564 244390 121592 245511
rect 121552 244384 121604 244390
rect 121552 244326 121604 244332
rect 121460 244248 121512 244254
rect 121460 244190 121512 244196
rect 121550 244216 121606 244225
rect 121550 244151 121606 244160
rect 121564 243030 121592 244151
rect 121552 243024 121604 243030
rect 121552 242966 121604 242972
rect 121552 242888 121604 242894
rect 121458 242856 121514 242865
rect 121552 242830 121604 242836
rect 121458 242791 121460 242800
rect 121512 242791 121514 242800
rect 121460 242762 121512 242768
rect 121564 242185 121592 242830
rect 121550 242176 121606 242185
rect 121550 242111 121606 242120
rect 121656 241505 121684 248386
rect 122102 243536 122158 243545
rect 122102 243471 122158 243480
rect 122116 242214 122144 243471
rect 122104 242208 122156 242214
rect 122104 242150 122156 242156
rect 121642 241496 121698 241505
rect 121642 241431 121698 241440
rect 121458 240816 121514 240825
rect 121656 240786 121684 241431
rect 122760 240825 122788 249358
rect 122852 247722 122880 249834
rect 122840 247716 122892 247722
rect 122840 247658 122892 247664
rect 122746 240816 122802 240825
rect 121458 240751 121514 240760
rect 121644 240780 121696 240786
rect 121472 240174 121500 240751
rect 122746 240751 122802 240760
rect 121644 240722 121696 240728
rect 121460 240168 121512 240174
rect 121460 240110 121512 240116
rect 122102 240136 122158 240145
rect 122102 240071 122158 240080
rect 122116 205154 122144 240071
rect 123588 237318 123616 274722
rect 123680 271182 123708 294238
rect 124128 291848 124180 291854
rect 124128 291790 124180 291796
rect 124140 275330 124168 291790
rect 124128 275324 124180 275330
rect 124128 275266 124180 275272
rect 123668 271176 123720 271182
rect 123668 271118 123720 271124
rect 124128 263560 124180 263566
rect 124128 263502 124180 263508
rect 124140 260166 124168 263502
rect 124128 260160 124180 260166
rect 124128 260102 124180 260108
rect 124232 249422 124260 331842
rect 124324 321570 124352 393926
rect 124494 379672 124550 379681
rect 124494 379607 124496 379616
rect 124548 379607 124550 379616
rect 124496 379578 124548 379584
rect 124404 368552 124456 368558
rect 124404 368494 124456 368500
rect 124416 334694 124444 368494
rect 125520 360330 125548 466414
rect 125600 463684 125652 463690
rect 125600 463626 125652 463632
rect 125612 463010 125640 463626
rect 125600 463004 125652 463010
rect 125600 462946 125652 462952
rect 125508 360324 125560 360330
rect 125508 360266 125560 360272
rect 125520 360126 125548 360266
rect 125508 360120 125560 360126
rect 125508 360062 125560 360068
rect 125612 354618 125640 462946
rect 125704 377466 125732 483006
rect 125796 437374 125824 534754
rect 125876 493332 125928 493338
rect 125876 493274 125928 493280
rect 125784 437368 125836 437374
rect 125784 437310 125836 437316
rect 125888 399498 125916 493274
rect 125980 463690 126008 555426
rect 126992 489190 127020 579702
rect 127072 539640 127124 539646
rect 127072 539582 127124 539588
rect 126980 489184 127032 489190
rect 126980 489126 127032 489132
rect 125968 463684 126020 463690
rect 125968 463626 126020 463632
rect 127084 447846 127112 539582
rect 128372 496126 128400 583782
rect 128452 581120 128504 581126
rect 128452 581062 128504 581068
rect 128360 496120 128412 496126
rect 127346 496088 127402 496097
rect 128360 496062 128412 496068
rect 127346 496023 127402 496032
rect 127164 493400 127216 493406
rect 127164 493342 127216 493348
rect 127072 447840 127124 447846
rect 127072 447782 127124 447788
rect 125968 399628 126020 399634
rect 125968 399570 126020 399576
rect 125876 399492 125928 399498
rect 125876 399434 125928 399440
rect 125784 395412 125836 395418
rect 125784 395354 125836 395360
rect 125692 377460 125744 377466
rect 125692 377402 125744 377408
rect 125600 354612 125652 354618
rect 125600 354554 125652 354560
rect 125612 353326 125640 354554
rect 125600 353320 125652 353326
rect 125600 353262 125652 353268
rect 124404 334688 124456 334694
rect 124404 334630 124456 334636
rect 125598 328400 125654 328409
rect 125598 328335 125654 328344
rect 125612 327894 125640 328335
rect 125600 327888 125652 327894
rect 125600 327830 125652 327836
rect 124312 321564 124364 321570
rect 124312 321506 124364 321512
rect 125508 321564 125560 321570
rect 125508 321506 125560 321512
rect 125520 320958 125548 321506
rect 125508 320952 125560 320958
rect 125508 320894 125560 320900
rect 124310 301472 124366 301481
rect 124310 301407 124366 301416
rect 124324 264625 124352 301407
rect 124864 298784 124916 298790
rect 124864 298726 124916 298732
rect 124310 264616 124366 264625
rect 124310 264551 124366 264560
rect 124324 262857 124352 264551
rect 124310 262848 124366 262857
rect 124310 262783 124366 262792
rect 124220 249416 124272 249422
rect 124220 249358 124272 249364
rect 124876 242962 124904 298726
rect 125612 255814 125640 327830
rect 125796 306338 125824 395354
rect 125876 377596 125928 377602
rect 125876 377538 125928 377544
rect 125888 376786 125916 377538
rect 125876 376780 125928 376786
rect 125876 376722 125928 376728
rect 125888 313954 125916 376722
rect 125980 329730 126008 399570
rect 126980 353320 127032 353326
rect 126980 353262 127032 353268
rect 125968 329724 126020 329730
rect 125968 329666 126020 329672
rect 126888 329724 126940 329730
rect 126888 329666 126940 329672
rect 126900 329118 126928 329666
rect 126888 329112 126940 329118
rect 126888 329054 126940 329060
rect 125876 313948 125928 313954
rect 125876 313890 125928 313896
rect 125784 306332 125836 306338
rect 125784 306274 125836 306280
rect 125796 305182 125824 306274
rect 125784 305176 125836 305182
rect 125784 305118 125836 305124
rect 126244 304292 126296 304298
rect 126244 304234 126296 304240
rect 125692 297424 125744 297430
rect 125692 297366 125744 297372
rect 125704 286550 125732 297366
rect 125692 286544 125744 286550
rect 125692 286486 125744 286492
rect 125704 284986 125732 286486
rect 125692 284980 125744 284986
rect 125692 284922 125744 284928
rect 125600 255808 125652 255814
rect 125600 255750 125652 255756
rect 125612 253230 125640 255750
rect 125600 253224 125652 253230
rect 125600 253166 125652 253172
rect 126256 244322 126284 304234
rect 126334 295488 126390 295497
rect 126334 295423 126390 295432
rect 126348 278050 126376 295423
rect 126336 278044 126388 278050
rect 126336 277986 126388 277992
rect 126244 244316 126296 244322
rect 126244 244258 126296 244264
rect 124864 242956 124916 242962
rect 124864 242898 124916 242904
rect 124876 239970 124904 242898
rect 126256 242826 126284 244258
rect 126244 242820 126296 242826
rect 126244 242762 126296 242768
rect 124864 239964 124916 239970
rect 124864 239906 124916 239912
rect 123576 237312 123628 237318
rect 123576 237254 123628 237260
rect 126992 230382 127020 353262
rect 127084 337958 127112 447782
rect 127176 391270 127204 493342
rect 127256 399560 127308 399566
rect 127256 399502 127308 399508
rect 127164 391264 127216 391270
rect 127164 391206 127216 391212
rect 127164 390788 127216 390794
rect 127164 390730 127216 390736
rect 127176 358766 127204 390730
rect 127164 358760 127216 358766
rect 127164 358702 127216 358708
rect 127072 337952 127124 337958
rect 127072 337894 127124 337900
rect 127268 333946 127296 399502
rect 127360 387122 127388 496023
rect 128360 494760 128412 494766
rect 128360 494702 128412 494708
rect 128372 397730 128400 494702
rect 128464 488510 128492 581062
rect 128636 581052 128688 581058
rect 128636 580994 128688 581000
rect 128544 541680 128596 541686
rect 128544 541622 128596 541628
rect 128556 541006 128584 541622
rect 128544 541000 128596 541006
rect 128544 540942 128596 540948
rect 128452 488504 128504 488510
rect 128452 488446 128504 488452
rect 128452 476128 128504 476134
rect 128452 476070 128504 476076
rect 128360 397724 128412 397730
rect 128360 397666 128412 397672
rect 128360 397588 128412 397594
rect 128360 397530 128412 397536
rect 128372 396778 128400 397530
rect 128360 396772 128412 396778
rect 128360 396714 128412 396720
rect 127348 387116 127400 387122
rect 127348 387058 127400 387064
rect 127532 387116 127584 387122
rect 127532 387058 127584 387064
rect 127544 387025 127572 387058
rect 127530 387016 127586 387025
rect 127530 386951 127586 386960
rect 128360 379636 128412 379642
rect 128360 379578 128412 379584
rect 127256 333940 127308 333946
rect 127256 333882 127308 333888
rect 127072 297492 127124 297498
rect 127072 297434 127124 297440
rect 127084 238814 127112 297434
rect 128372 242894 128400 379578
rect 128464 368558 128492 476070
rect 128556 445126 128584 540942
rect 128648 500342 128676 580994
rect 130016 571396 130068 571402
rect 130016 571338 130068 571344
rect 129922 554024 129978 554033
rect 129922 553959 129978 553968
rect 129832 537600 129884 537606
rect 129832 537542 129884 537548
rect 128636 500336 128688 500342
rect 128636 500278 128688 500284
rect 129004 496188 129056 496194
rect 129004 496130 129056 496136
rect 128544 445120 128596 445126
rect 128542 445088 128544 445097
rect 128596 445088 128598 445097
rect 128542 445023 128598 445032
rect 128544 398132 128596 398138
rect 128544 398074 128596 398080
rect 128452 368552 128504 368558
rect 128452 368494 128504 368500
rect 128452 360324 128504 360330
rect 128452 360266 128504 360272
rect 128464 286482 128492 360266
rect 128556 307766 128584 398074
rect 128728 397724 128780 397730
rect 128728 397666 128780 397672
rect 128636 396908 128688 396914
rect 128636 396850 128688 396856
rect 128648 324290 128676 396850
rect 128740 394126 128768 397666
rect 129016 397594 129044 496130
rect 129738 493368 129794 493377
rect 129738 493303 129794 493312
rect 129004 397588 129056 397594
rect 129004 397530 129056 397536
rect 129752 394194 129780 493303
rect 129844 441590 129872 537542
rect 129936 462330 129964 553959
rect 130028 480962 130056 571338
rect 130396 537985 130424 630634
rect 136652 596834 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700398 154160 703520
rect 170324 702434 170352 703520
rect 202800 703322 202828 703520
rect 201500 703316 201552 703322
rect 201500 703258 201552 703264
rect 202788 703316 202840 703322
rect 202788 703258 202840 703264
rect 169772 702406 170352 702434
rect 154120 700392 154172 700398
rect 154120 700334 154172 700340
rect 155224 700392 155276 700398
rect 155224 700334 155276 700340
rect 136640 596828 136692 596834
rect 136640 596770 136692 596776
rect 155236 587178 155264 700334
rect 159364 683188 159416 683194
rect 159364 683130 159416 683136
rect 155224 587172 155276 587178
rect 155224 587114 155276 587120
rect 136640 584044 136692 584050
rect 136640 583986 136692 583992
rect 131120 578264 131172 578270
rect 131120 578206 131172 578212
rect 130382 537976 130438 537985
rect 130382 537911 130438 537920
rect 131132 487150 131160 578206
rect 132592 564528 132644 564534
rect 132592 564470 132644 564476
rect 131396 560380 131448 560386
rect 131396 560322 131448 560328
rect 131212 497480 131264 497486
rect 131212 497422 131264 497428
rect 131120 487144 131172 487150
rect 131120 487086 131172 487092
rect 130016 480956 130068 480962
rect 130016 480898 130068 480904
rect 129924 462324 129976 462330
rect 129924 462266 129976 462272
rect 130384 462324 130436 462330
rect 130384 462266 130436 462272
rect 130396 461145 130424 462266
rect 130382 461136 130438 461145
rect 130382 461071 130438 461080
rect 129832 441584 129884 441590
rect 129832 441526 129884 441532
rect 129844 440910 129872 441526
rect 129832 440904 129884 440910
rect 129832 440846 129884 440852
rect 131120 440360 131172 440366
rect 131120 440302 131172 440308
rect 129924 403708 129976 403714
rect 129924 403650 129976 403656
rect 129740 394188 129792 394194
rect 129740 394130 129792 394136
rect 128728 394120 128780 394126
rect 128728 394062 128780 394068
rect 128740 393990 128768 394062
rect 128728 393984 128780 393990
rect 128728 393926 128780 393932
rect 129740 393984 129792 393990
rect 129740 393926 129792 393932
rect 128818 335336 128874 335345
rect 128818 335271 128874 335280
rect 128832 335238 128860 335271
rect 128820 335232 128872 335238
rect 128820 335174 128872 335180
rect 128636 324284 128688 324290
rect 128636 324226 128688 324232
rect 128648 323610 128676 324226
rect 128636 323604 128688 323610
rect 128636 323546 128688 323552
rect 128544 307760 128596 307766
rect 128544 307702 128596 307708
rect 128728 307760 128780 307766
rect 128728 307702 128780 307708
rect 128740 307222 128768 307702
rect 128728 307216 128780 307222
rect 128728 307158 128780 307164
rect 128544 305176 128596 305182
rect 128544 305118 128596 305124
rect 128452 286476 128504 286482
rect 128452 286418 128504 286424
rect 128464 279478 128492 286418
rect 128452 279472 128504 279478
rect 128452 279414 128504 279420
rect 128360 242888 128412 242894
rect 128360 242830 128412 242836
rect 127072 238808 127124 238814
rect 127072 238750 127124 238756
rect 128556 238066 128584 305118
rect 129752 292890 129780 393926
rect 129832 358760 129884 358766
rect 129832 358702 129884 358708
rect 129660 292862 129780 292890
rect 129660 291854 129688 292862
rect 129738 292768 129794 292777
rect 129738 292703 129794 292712
rect 129648 291848 129700 291854
rect 129648 291790 129700 291796
rect 129752 287774 129780 292703
rect 129740 287768 129792 287774
rect 129740 287710 129792 287716
rect 129844 274786 129872 358702
rect 129936 339522 129964 403650
rect 130016 398200 130068 398206
rect 130016 398142 130068 398148
rect 129924 339516 129976 339522
rect 129924 339458 129976 339464
rect 130028 339386 130056 398142
rect 130106 342952 130162 342961
rect 130106 342887 130108 342896
rect 130160 342887 130162 342896
rect 130108 342858 130160 342864
rect 130016 339380 130068 339386
rect 130016 339322 130068 339328
rect 131132 338094 131160 440302
rect 131224 394058 131252 497422
rect 131304 487144 131356 487150
rect 131304 487086 131356 487092
rect 131316 486470 131344 487086
rect 131304 486464 131356 486470
rect 131304 486406 131356 486412
rect 131304 485104 131356 485110
rect 131304 485046 131356 485052
rect 131316 395350 131344 485046
rect 131408 469946 131436 560322
rect 132500 493468 132552 493474
rect 132500 493410 132552 493416
rect 131488 488572 131540 488578
rect 131488 488514 131540 488520
rect 131500 485110 131528 488514
rect 131488 485104 131540 485110
rect 131488 485046 131540 485052
rect 131396 469940 131448 469946
rect 131396 469882 131448 469888
rect 131304 395344 131356 395350
rect 131304 395286 131356 395292
rect 131212 394052 131264 394058
rect 131212 393994 131264 394000
rect 132512 392766 132540 493410
rect 132604 472054 132632 564470
rect 135444 561740 135496 561746
rect 135444 561682 135496 561688
rect 133972 560312 134024 560318
rect 133972 560254 134024 560260
rect 132776 559020 132828 559026
rect 132776 558962 132828 558968
rect 132684 537532 132736 537538
rect 132684 537474 132736 537480
rect 132592 472048 132644 472054
rect 132592 471990 132644 471996
rect 132500 392760 132552 392766
rect 132500 392702 132552 392708
rect 132498 392048 132554 392057
rect 132498 391983 132554 391992
rect 131212 389972 131264 389978
rect 131212 389914 131264 389920
rect 131120 338088 131172 338094
rect 131120 338030 131172 338036
rect 131224 303006 131252 389914
rect 131304 385756 131356 385762
rect 131304 385698 131356 385704
rect 131316 318714 131344 385698
rect 131304 318708 131356 318714
rect 131304 318650 131356 318656
rect 131672 318708 131724 318714
rect 131672 318650 131724 318656
rect 131684 318170 131712 318650
rect 131672 318164 131724 318170
rect 131672 318106 131724 318112
rect 131212 303000 131264 303006
rect 131212 302942 131264 302948
rect 131118 293176 131174 293185
rect 131118 293111 131174 293120
rect 130384 286408 130436 286414
rect 130384 286350 130436 286356
rect 129832 274780 129884 274786
rect 129832 274722 129884 274728
rect 130396 264246 130424 286350
rect 130384 264240 130436 264246
rect 130384 264182 130436 264188
rect 131132 255270 131160 293111
rect 132512 282849 132540 391983
rect 132604 365090 132632 471990
rect 132696 445058 132724 537474
rect 132788 468489 132816 558962
rect 133880 558952 133932 558958
rect 133880 558894 133932 558900
rect 132774 468480 132830 468489
rect 132774 468415 132830 468424
rect 133892 467158 133920 558894
rect 133984 480254 134012 560254
rect 135168 559564 135220 559570
rect 135168 559506 135220 559512
rect 135180 558958 135208 559506
rect 135168 558952 135220 558958
rect 135168 558894 135220 558900
rect 134248 549364 134300 549370
rect 134248 549306 134300 549312
rect 134156 542428 134208 542434
rect 134156 542370 134208 542376
rect 133984 480226 134104 480254
rect 134076 469878 134104 480226
rect 134064 469872 134116 469878
rect 134064 469814 134116 469820
rect 133880 467152 133932 467158
rect 133880 467094 133932 467100
rect 133972 459604 134024 459610
rect 133972 459546 134024 459552
rect 132684 445052 132736 445058
rect 132684 444994 132736 445000
rect 132684 400920 132736 400926
rect 132684 400862 132736 400868
rect 132774 400888 132830 400897
rect 132592 365084 132644 365090
rect 132592 365026 132644 365032
rect 132604 303074 132632 365026
rect 132696 317422 132724 400862
rect 132774 400823 132830 400832
rect 132788 320142 132816 400823
rect 133880 389360 133932 389366
rect 133880 389302 133932 389308
rect 132776 320136 132828 320142
rect 132776 320078 132828 320084
rect 133788 320136 133840 320142
rect 133788 320078 133840 320084
rect 133800 319530 133828 320078
rect 133788 319524 133840 319530
rect 133788 319466 133840 319472
rect 132684 317416 132736 317422
rect 132684 317358 132736 317364
rect 133788 317416 133840 317422
rect 133788 317358 133840 317364
rect 133800 316742 133828 317358
rect 133788 316736 133840 316742
rect 133788 316678 133840 316684
rect 132592 303068 132644 303074
rect 132592 303010 132644 303016
rect 132592 300212 132644 300218
rect 132592 300154 132644 300160
rect 132498 282840 132554 282849
rect 132498 282775 132554 282784
rect 131120 255264 131172 255270
rect 131120 255206 131172 255212
rect 131488 255264 131540 255270
rect 131488 255206 131540 255212
rect 131500 254590 131528 255206
rect 131488 254584 131540 254590
rect 131488 254526 131540 254532
rect 132604 238746 132632 300154
rect 133144 296948 133196 296954
rect 133144 296890 133196 296896
rect 132592 238740 132644 238746
rect 132592 238682 132644 238688
rect 128544 238060 128596 238066
rect 128544 238002 128596 238008
rect 126980 230376 127032 230382
rect 126980 230318 127032 230324
rect 127440 230376 127492 230382
rect 127440 230318 127492 230324
rect 127452 229838 127480 230318
rect 127440 229832 127492 229838
rect 127440 229774 127492 229780
rect 122104 205148 122156 205154
rect 122104 205090 122156 205096
rect 120080 203584 120132 203590
rect 120080 203526 120132 203532
rect 133156 198121 133184 296890
rect 133786 282840 133842 282849
rect 133786 282775 133842 282784
rect 133800 282169 133828 282775
rect 133786 282160 133842 282169
rect 133786 282095 133842 282104
rect 133788 238740 133840 238746
rect 133788 238682 133840 238688
rect 133800 238066 133828 238682
rect 133788 238060 133840 238066
rect 133788 238002 133840 238008
rect 133892 205630 133920 389302
rect 133984 336666 134012 459546
rect 134076 362234 134104 469814
rect 134168 451926 134196 542370
rect 134260 458862 134288 549306
rect 135352 546508 135404 546514
rect 135352 546450 135404 546456
rect 135260 500268 135312 500274
rect 135260 500210 135312 500216
rect 134248 458856 134300 458862
rect 134248 458798 134300 458804
rect 134156 451920 134208 451926
rect 134156 451862 134208 451868
rect 135272 388550 135300 500210
rect 135364 454714 135392 546450
rect 135456 471374 135484 561682
rect 136652 491298 136680 583986
rect 138020 576904 138072 576910
rect 138020 576846 138072 576852
rect 136732 570036 136784 570042
rect 136732 569978 136784 569984
rect 136640 491292 136692 491298
rect 136640 491234 136692 491240
rect 136744 477358 136772 569978
rect 136824 556232 136876 556238
rect 136824 556174 136876 556180
rect 136732 477352 136784 477358
rect 136732 477294 136784 477300
rect 135444 471368 135496 471374
rect 135444 471310 135496 471316
rect 136836 465730 136864 556174
rect 136916 496120 136968 496126
rect 136916 496062 136968 496068
rect 136824 465724 136876 465730
rect 136824 465666 136876 465672
rect 135352 454708 135404 454714
rect 135352 454650 135404 454656
rect 135260 388544 135312 388550
rect 135260 388486 135312 388492
rect 134524 367872 134576 367878
rect 134524 367814 134576 367820
rect 134064 362228 134116 362234
rect 134064 362170 134116 362176
rect 134062 353696 134118 353705
rect 134062 353631 134118 353640
rect 134076 353258 134104 353631
rect 134064 353252 134116 353258
rect 134064 353194 134116 353200
rect 133972 336660 134024 336666
rect 133972 336602 134024 336608
rect 133972 335232 134024 335238
rect 133972 335174 134024 335180
rect 133984 240106 134012 335174
rect 134536 267734 134564 367814
rect 135364 346390 135392 454650
rect 136824 440292 136876 440298
rect 136824 440234 136876 440240
rect 135444 398268 135496 398274
rect 135444 398210 135496 398216
rect 135352 346384 135404 346390
rect 135352 346326 135404 346332
rect 135456 340814 135484 398210
rect 136640 392760 136692 392766
rect 136640 392702 136692 392708
rect 136548 388544 136600 388550
rect 136548 388486 136600 388492
rect 136560 388385 136588 388486
rect 136546 388376 136602 388385
rect 136546 388311 136602 388320
rect 135904 360256 135956 360262
rect 135904 360198 135956 360204
rect 135444 340808 135496 340814
rect 135444 340750 135496 340756
rect 135168 336660 135220 336666
rect 135168 336602 135220 336608
rect 135180 336054 135208 336602
rect 135168 336048 135220 336054
rect 135168 335990 135220 335996
rect 135916 311166 135944 360198
rect 136548 346384 136600 346390
rect 136548 346326 136600 346332
rect 136560 345710 136588 346326
rect 136548 345704 136600 345710
rect 136548 345646 136600 345652
rect 135904 311160 135956 311166
rect 135904 311102 135956 311108
rect 135904 295656 135956 295662
rect 135904 295598 135956 295604
rect 134536 267706 134748 267734
rect 134720 262274 134748 267706
rect 134708 262268 134760 262274
rect 134708 262210 134760 262216
rect 134720 260846 134748 262210
rect 134708 260840 134760 260846
rect 134708 260782 134760 260788
rect 135916 250510 135944 295598
rect 135904 250504 135956 250510
rect 135904 250446 135956 250452
rect 133972 240100 134024 240106
rect 133972 240042 134024 240048
rect 134524 240100 134576 240106
rect 134524 240042 134576 240048
rect 134536 231130 134564 240042
rect 136652 235958 136680 392702
rect 136836 331226 136864 440234
rect 136928 385694 136956 496062
rect 138032 487830 138060 576846
rect 159376 574054 159404 683130
rect 159364 574048 159416 574054
rect 159364 573990 159416 573996
rect 139400 569968 139452 569974
rect 139400 569910 139452 569916
rect 138204 545148 138256 545154
rect 138204 545090 138256 545096
rect 138020 487824 138072 487830
rect 138020 487766 138072 487772
rect 137008 478916 137060 478922
rect 137008 478858 137060 478864
rect 136916 385688 136968 385694
rect 136916 385630 136968 385636
rect 137020 367062 137048 478858
rect 138112 465724 138164 465730
rect 138112 465666 138164 465672
rect 138018 461000 138074 461009
rect 138018 460935 138074 460944
rect 137008 367056 137060 367062
rect 137008 366998 137060 367004
rect 137192 367056 137244 367062
rect 137192 366998 137244 367004
rect 137204 366382 137232 366998
rect 137192 366376 137244 366382
rect 137192 366318 137244 366324
rect 138032 351898 138060 460935
rect 138124 357406 138152 465666
rect 138216 454782 138244 545090
rect 139412 476066 139440 569910
rect 140872 565888 140924 565894
rect 140872 565830 140924 565836
rect 139584 547936 139636 547942
rect 139584 547878 139636 547884
rect 139400 476060 139452 476066
rect 139400 476002 139452 476008
rect 139492 469940 139544 469946
rect 139492 469882 139544 469888
rect 138204 454776 138256 454782
rect 138204 454718 138256 454724
rect 139400 394800 139452 394806
rect 139400 394742 139452 394748
rect 138204 386504 138256 386510
rect 138204 386446 138256 386452
rect 138112 357400 138164 357406
rect 138112 357342 138164 357348
rect 138020 351892 138072 351898
rect 138020 351834 138072 351840
rect 138032 351286 138060 351834
rect 138020 351280 138072 351286
rect 138020 351222 138072 351228
rect 138020 340808 138072 340814
rect 138020 340750 138072 340756
rect 137282 336152 137338 336161
rect 137282 336087 137338 336096
rect 136824 331220 136876 331226
rect 136824 331162 136876 331168
rect 137100 331220 137152 331226
rect 137100 331162 137152 331168
rect 137112 330546 137140 331162
rect 137100 330540 137152 330546
rect 137100 330482 137152 330488
rect 137296 259486 137324 336087
rect 137284 259480 137336 259486
rect 137284 259422 137336 259428
rect 138032 237386 138060 340750
rect 138216 309126 138244 386446
rect 138204 309120 138256 309126
rect 138204 309062 138256 309068
rect 138664 309120 138716 309126
rect 138664 309062 138716 309068
rect 138676 308514 138704 309062
rect 138664 308508 138716 308514
rect 138664 308450 138716 308456
rect 138020 237380 138072 237386
rect 138020 237322 138072 237328
rect 138032 236706 138060 237322
rect 138020 236700 138072 236706
rect 138020 236642 138072 236648
rect 136640 235952 136692 235958
rect 136640 235894 136692 235900
rect 134524 231124 134576 231130
rect 134524 231066 134576 231072
rect 139412 212537 139440 394742
rect 139504 360262 139532 469882
rect 139596 457502 139624 547878
rect 140884 474706 140912 565830
rect 143448 564460 143500 564466
rect 143448 564402 143500 564408
rect 140964 554056 141016 554062
rect 140964 553998 141016 554004
rect 140976 553450 141004 553998
rect 140964 553444 141016 553450
rect 140964 553386 141016 553392
rect 140872 474700 140924 474706
rect 140872 474642 140924 474648
rect 140976 462398 141004 553386
rect 142160 549296 142212 549302
rect 142160 549238 142212 549244
rect 141146 490512 141202 490521
rect 141146 490447 141202 490456
rect 140964 462392 141016 462398
rect 140964 462334 141016 462340
rect 139584 457496 139636 457502
rect 139584 457438 139636 457444
rect 139584 440904 139636 440910
rect 139584 440846 139636 440852
rect 139492 360256 139544 360262
rect 139492 360198 139544 360204
rect 139596 336734 139624 440846
rect 140780 390652 140832 390658
rect 140780 390594 140832 390600
rect 139584 336728 139636 336734
rect 139584 336670 139636 336676
rect 140792 262206 140820 390594
rect 140872 357400 140924 357406
rect 140872 357342 140924 357348
rect 140780 262200 140832 262206
rect 140780 262142 140832 262148
rect 140792 261526 140820 262142
rect 140780 261520 140832 261526
rect 140780 261462 140832 261468
rect 140884 234433 140912 357342
rect 140976 354686 141004 462334
rect 141056 403640 141108 403646
rect 141056 403582 141108 403588
rect 140964 354680 141016 354686
rect 140964 354622 141016 354628
rect 140976 354074 141004 354622
rect 140964 354068 141016 354074
rect 140964 354010 141016 354016
rect 141068 325694 141096 403582
rect 141160 387977 141188 490447
rect 141240 474700 141292 474706
rect 141240 474642 141292 474648
rect 141252 474026 141280 474642
rect 141240 474020 141292 474026
rect 141240 473962 141292 473968
rect 142172 456754 142200 549238
rect 142344 486464 142396 486470
rect 142344 486406 142396 486412
rect 142252 457496 142304 457502
rect 142252 457438 142304 457444
rect 142160 456748 142212 456754
rect 142160 456690 142212 456696
rect 142160 445052 142212 445058
rect 142160 444994 142212 445000
rect 141146 387968 141202 387977
rect 141146 387903 141202 387912
rect 142172 332586 142200 444994
rect 142264 345778 142292 457438
rect 142356 382226 142384 486406
rect 143460 473362 143488 564402
rect 169772 535430 169800 702406
rect 201512 559570 201540 703258
rect 218992 700398 219020 703520
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 235184 700330 235212 703520
rect 267660 703254 267688 703520
rect 267648 703248 267700 703254
rect 267648 703190 267700 703196
rect 283852 700330 283880 703520
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 238024 700324 238076 700330
rect 238024 700266 238076 700272
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 238036 585818 238064 700266
rect 238024 585812 238076 585818
rect 238024 585754 238076 585760
rect 204904 564460 204956 564466
rect 204904 564402 204956 564408
rect 201500 559564 201552 559570
rect 201500 559506 201552 559512
rect 204916 538218 204944 564402
rect 299492 541686 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703186 332548 703520
rect 332508 703180 332560 703186
rect 332508 703122 332560 703128
rect 348804 703118 348832 703520
rect 348792 703112 348844 703118
rect 348792 703054 348844 703060
rect 364996 703050 365024 703520
rect 364984 703044 365036 703050
rect 364984 702986 365036 702992
rect 364996 701729 365024 702986
rect 381544 702840 381596 702846
rect 381544 702782 381596 702788
rect 386420 702840 386472 702846
rect 386420 702782 386472 702788
rect 364982 701720 365038 701729
rect 364982 701655 365038 701664
rect 374644 563712 374696 563718
rect 374644 563654 374696 563660
rect 299480 541680 299532 541686
rect 299480 541622 299532 541628
rect 204904 538212 204956 538218
rect 204904 538154 204956 538160
rect 169760 535424 169812 535430
rect 169760 535366 169812 535372
rect 147680 487824 147732 487830
rect 147680 487766 147732 487772
rect 144920 474020 144972 474026
rect 144920 473962 144972 473968
rect 143460 473334 143580 473362
rect 143552 472666 143580 473334
rect 143540 472660 143592 472666
rect 143540 472602 143592 472608
rect 143448 456748 143500 456754
rect 143448 456690 143500 456696
rect 143460 456074 143488 456690
rect 143448 456068 143500 456074
rect 143448 456010 143500 456016
rect 142436 391264 142488 391270
rect 142436 391206 142488 391212
rect 142344 382220 142396 382226
rect 142344 382162 142396 382168
rect 142252 345772 142304 345778
rect 142252 345714 142304 345720
rect 142252 340944 142304 340950
rect 142252 340886 142304 340892
rect 142160 332580 142212 332586
rect 142160 332522 142212 332528
rect 140976 325666 141096 325694
rect 140976 322930 141004 325666
rect 140964 322924 141016 322930
rect 140964 322866 141016 322872
rect 140976 322318 141004 322866
rect 140964 322312 141016 322318
rect 140964 322254 141016 322260
rect 142264 244254 142292 340886
rect 142448 288386 142476 391206
rect 143448 382220 143500 382226
rect 143448 382162 143500 382168
rect 143460 381546 143488 382162
rect 143448 381540 143500 381546
rect 143448 381482 143500 381488
rect 143552 366450 143580 472602
rect 143632 471368 143684 471374
rect 143632 471310 143684 471316
rect 143540 366444 143592 366450
rect 143540 366386 143592 366392
rect 143448 332580 143500 332586
rect 143448 332522 143500 332528
rect 143460 331906 143488 332522
rect 143448 331900 143500 331906
rect 143448 331842 143500 331848
rect 142804 292868 142856 292874
rect 142804 292810 142856 292816
rect 142436 288380 142488 288386
rect 142436 288322 142488 288328
rect 142252 244248 142304 244254
rect 142252 244190 142304 244196
rect 140870 234424 140926 234433
rect 140870 234359 140926 234368
rect 139398 212528 139454 212537
rect 139398 212463 139454 212472
rect 139412 211857 139440 212463
rect 139398 211848 139454 211857
rect 139398 211783 139454 211792
rect 133880 205624 133932 205630
rect 133880 205566 133932 205572
rect 135168 205624 135220 205630
rect 135168 205566 135220 205572
rect 135180 204950 135208 205566
rect 135168 204944 135220 204950
rect 135168 204886 135220 204892
rect 133142 198112 133198 198121
rect 133142 198047 133198 198056
rect 118700 188488 118752 188494
rect 118700 188430 118752 188436
rect 131028 187740 131080 187746
rect 131028 187682 131080 187688
rect 129648 183592 129700 183598
rect 129648 183534 129700 183540
rect 115940 182980 115992 182986
rect 115940 182922 115992 182928
rect 119528 182232 119580 182238
rect 119528 182174 119580 182180
rect 116952 180872 117004 180878
rect 116952 180814 117004 180820
rect 115848 179580 115900 179586
rect 115848 179522 115900 179528
rect 112260 179444 112312 179450
rect 112260 179386 112312 179392
rect 112272 176905 112300 179386
rect 114376 178288 114428 178294
rect 114376 178230 114428 178236
rect 112258 176896 112314 176905
rect 111064 176860 111116 176866
rect 112258 176831 112314 176840
rect 111064 176802 111116 176808
rect 110696 176792 110748 176798
rect 109774 176760 109830 176769
rect 109774 176695 109830 176704
rect 110694 176760 110696 176769
rect 114388 176769 114416 178230
rect 115860 177177 115888 179522
rect 116964 177721 116992 180814
rect 118424 178016 118476 178022
rect 118424 177958 118476 177964
rect 116950 177712 117006 177721
rect 116950 177647 117006 177656
rect 115846 177168 115902 177177
rect 115846 177103 115902 177112
rect 118436 176769 118464 177958
rect 119540 177721 119568 182174
rect 122012 180940 122064 180946
rect 122012 180882 122064 180888
rect 121000 179648 121052 179654
rect 121000 179590 121052 179596
rect 119526 177712 119582 177721
rect 119526 177647 119582 177656
rect 121012 177177 121040 179590
rect 122024 177721 122052 180882
rect 127072 178152 127124 178158
rect 127072 178094 127124 178100
rect 122010 177712 122066 177721
rect 122010 177647 122066 177656
rect 120998 177168 121054 177177
rect 120998 177103 121054 177112
rect 125784 176928 125836 176934
rect 125784 176870 125836 176876
rect 124496 176860 124548 176866
rect 124496 176802 124548 176808
rect 124508 176769 124536 176802
rect 125796 176769 125824 176870
rect 127084 176769 127112 178094
rect 129660 177721 129688 183534
rect 131040 177721 131068 187682
rect 142816 183054 142844 292810
rect 143448 288380 143500 288386
rect 143448 288322 143500 288328
rect 143460 287706 143488 288322
rect 143448 287700 143500 287706
rect 143448 287642 143500 287648
rect 143448 244248 143500 244254
rect 143448 244190 143500 244196
rect 143460 243574 143488 244190
rect 143448 243568 143500 243574
rect 143448 243510 143500 243516
rect 143552 229094 143580 366386
rect 143644 362914 143672 471310
rect 143724 390720 143776 390726
rect 143724 390662 143776 390668
rect 143632 362908 143684 362914
rect 143632 362850 143684 362856
rect 143736 316034 143764 390662
rect 144932 367810 144960 473962
rect 146300 471300 146352 471306
rect 146300 471242 146352 471248
rect 146312 470626 146340 471242
rect 146300 470620 146352 470626
rect 146300 470562 146352 470568
rect 145012 382288 145064 382294
rect 145012 382230 145064 382236
rect 144920 367804 144972 367810
rect 144920 367746 144972 367752
rect 144828 362908 144880 362914
rect 144828 362850 144880 362856
rect 144840 362234 144868 362850
rect 144828 362228 144880 362234
rect 144828 362170 144880 362176
rect 143644 316006 143764 316034
rect 143644 306338 143672 316006
rect 145024 309874 145052 382230
rect 146312 365022 146340 470562
rect 146392 445800 146444 445806
rect 146392 445742 146444 445748
rect 146300 365016 146352 365022
rect 146300 364958 146352 364964
rect 146300 353320 146352 353326
rect 146300 353262 146352 353268
rect 145012 309868 145064 309874
rect 145012 309810 145064 309816
rect 143632 306332 143684 306338
rect 143632 306274 143684 306280
rect 143644 305726 143672 306274
rect 143632 305720 143684 305726
rect 143632 305662 143684 305668
rect 144184 294228 144236 294234
rect 144184 294170 144236 294176
rect 143552 229066 143672 229094
rect 143644 219337 143672 229066
rect 143630 219328 143686 219337
rect 143630 219263 143686 219272
rect 143644 218657 143672 219263
rect 143630 218648 143686 218657
rect 143630 218583 143686 218592
rect 144196 199578 144224 294170
rect 146312 222154 146340 353262
rect 146404 327078 146432 445742
rect 146576 390584 146628 390590
rect 146576 390526 146628 390532
rect 146484 389292 146536 389298
rect 146484 389234 146536 389240
rect 146392 327072 146444 327078
rect 146392 327014 146444 327020
rect 146496 294642 146524 389234
rect 146588 307086 146616 390526
rect 147692 381614 147720 487766
rect 150624 481704 150676 481710
rect 150624 481646 150676 481652
rect 147864 480956 147916 480962
rect 147864 480898 147916 480904
rect 147772 451920 147824 451926
rect 147772 451862 147824 451868
rect 147680 381608 147732 381614
rect 147680 381550 147732 381556
rect 147692 380934 147720 381550
rect 147680 380928 147732 380934
rect 147680 380870 147732 380876
rect 147680 375352 147732 375358
rect 147680 375294 147732 375300
rect 147692 374678 147720 375294
rect 147680 374672 147732 374678
rect 147680 374614 147732 374620
rect 147680 354068 147732 354074
rect 147680 354010 147732 354016
rect 146760 327072 146812 327078
rect 146760 327014 146812 327020
rect 146772 326398 146800 327014
rect 146760 326392 146812 326398
rect 146760 326334 146812 326340
rect 146576 307080 146628 307086
rect 146576 307022 146628 307028
rect 146484 294636 146536 294642
rect 146484 294578 146536 294584
rect 146942 291952 146998 291961
rect 146942 291887 146998 291896
rect 146300 222148 146352 222154
rect 146300 222090 146352 222096
rect 146760 222148 146812 222154
rect 146760 222090 146812 222096
rect 146772 221542 146800 222090
rect 146760 221536 146812 221542
rect 146760 221478 146812 221484
rect 144184 199572 144236 199578
rect 144184 199514 144236 199520
rect 146956 187134 146984 291887
rect 147692 217462 147720 354010
rect 147784 340882 147812 451862
rect 147876 375358 147904 480898
rect 149244 458856 149296 458862
rect 149244 458798 149296 458804
rect 149150 451344 149206 451353
rect 149150 451279 149206 451288
rect 147956 380928 148008 380934
rect 147956 380870 148008 380876
rect 147864 375352 147916 375358
rect 147864 375294 147916 375300
rect 147772 340876 147824 340882
rect 147772 340818 147824 340824
rect 147784 340202 147812 340818
rect 147772 340196 147824 340202
rect 147772 340138 147824 340144
rect 147968 298353 147996 380870
rect 149060 376712 149112 376718
rect 149060 376654 149112 376660
rect 149072 375426 149100 376654
rect 149060 375420 149112 375426
rect 149060 375362 149112 375368
rect 147954 298344 148010 298353
rect 147954 298279 148010 298288
rect 147968 296714 147996 298279
rect 147968 296686 148364 296714
rect 148336 283626 148364 296686
rect 148324 283620 148376 283626
rect 148324 283562 148376 283568
rect 149072 230450 149100 375362
rect 149164 335306 149192 451279
rect 149256 345030 149284 458798
rect 150532 454776 150584 454782
rect 150532 454718 150584 454724
rect 150440 393984 150492 393990
rect 150440 393926 150492 393932
rect 149244 345024 149296 345030
rect 149244 344966 149296 344972
rect 149256 344350 149284 344966
rect 149244 344344 149296 344350
rect 149244 344286 149296 344292
rect 149152 335300 149204 335306
rect 149152 335242 149204 335248
rect 149164 334665 149192 335242
rect 149150 334656 149206 334665
rect 149150 334591 149206 334600
rect 150452 269074 150480 393926
rect 150544 342242 150572 454718
rect 150636 376718 150664 481646
rect 151818 480312 151874 480321
rect 151818 480247 151874 480256
rect 150624 376712 150676 376718
rect 150624 376654 150676 376660
rect 151832 371210 151860 480247
rect 152002 468480 152058 468489
rect 152002 468415 152058 468424
rect 151912 456068 151964 456074
rect 151912 456010 151964 456016
rect 151820 371204 151872 371210
rect 151820 371146 151872 371152
rect 151820 369912 151872 369918
rect 151820 369854 151872 369860
rect 150532 342236 150584 342242
rect 150532 342178 150584 342184
rect 150992 342236 151044 342242
rect 150992 342178 151044 342184
rect 151004 341562 151032 342178
rect 150992 341556 151044 341562
rect 150992 341498 151044 341504
rect 151084 314016 151136 314022
rect 151084 313958 151136 313964
rect 150440 269068 150492 269074
rect 150440 269010 150492 269016
rect 150452 268394 150480 269010
rect 150440 268388 150492 268394
rect 150440 268330 150492 268336
rect 149060 230444 149112 230450
rect 149060 230386 149112 230392
rect 147680 217456 147732 217462
rect 147680 217398 147732 217404
rect 147692 216730 147720 217398
rect 147600 216702 147720 216730
rect 147600 188329 147628 216702
rect 147586 188320 147642 188329
rect 147586 188255 147642 188264
rect 146944 187128 146996 187134
rect 146944 187070 146996 187076
rect 151096 184482 151124 313958
rect 151832 215286 151860 369854
rect 151924 347750 151952 456010
rect 152016 360194 152044 468415
rect 336002 405784 336058 405793
rect 336002 405719 336058 405728
rect 304264 401668 304316 401674
rect 304264 401610 304316 401616
rect 166262 400344 166318 400353
rect 166262 400279 166318 400288
rect 153108 371204 153160 371210
rect 153108 371146 153160 371152
rect 153120 370569 153148 371146
rect 153106 370560 153162 370569
rect 153106 370495 153162 370504
rect 152004 360188 152056 360194
rect 152004 360130 152056 360136
rect 153108 360188 153160 360194
rect 153108 360130 153160 360136
rect 153120 359514 153148 360130
rect 153108 359508 153160 359514
rect 153108 359450 153160 359456
rect 151912 347744 151964 347750
rect 151912 347686 151964 347692
rect 153108 347744 153160 347750
rect 153108 347686 153160 347692
rect 153120 347070 153148 347686
rect 153108 347064 153160 347070
rect 153108 347006 153160 347012
rect 159364 315308 159416 315314
rect 159364 315250 159416 315256
rect 155316 309188 155368 309194
rect 155316 309130 155368 309136
rect 153844 307828 153896 307834
rect 153844 307770 153896 307776
rect 151820 215280 151872 215286
rect 151820 215222 151872 215228
rect 153108 215280 153160 215286
rect 153108 215222 153160 215228
rect 153120 214606 153148 215222
rect 153108 214600 153160 214606
rect 153108 214542 153160 214548
rect 153856 185910 153884 307770
rect 155224 307216 155276 307222
rect 155224 307158 155276 307164
rect 155236 193866 155264 307158
rect 155328 197985 155356 309130
rect 157984 232756 158036 232762
rect 157984 232698 158036 232704
rect 157996 202298 158024 232698
rect 157984 202292 158036 202298
rect 157984 202234 158036 202240
rect 155314 197976 155370 197985
rect 155314 197911 155370 197920
rect 155224 193860 155276 193866
rect 155224 193802 155276 193808
rect 153844 185904 153896 185910
rect 153844 185846 153896 185852
rect 151084 184476 151136 184482
rect 151084 184418 151136 184424
rect 142804 183048 142856 183054
rect 142804 182990 142856 182996
rect 132408 181008 132460 181014
rect 132408 180950 132460 180956
rect 132420 177721 132448 180950
rect 159376 180198 159404 315250
rect 162124 311228 162176 311234
rect 162124 311170 162176 311176
rect 160744 295588 160796 295594
rect 160744 295530 160796 295536
rect 159456 294160 159508 294166
rect 159456 294102 159508 294108
rect 159468 247790 159496 294102
rect 159456 247784 159508 247790
rect 159456 247726 159508 247732
rect 160756 192574 160784 295530
rect 160744 192568 160796 192574
rect 160744 192510 160796 192516
rect 162136 181762 162164 311170
rect 162214 292632 162270 292641
rect 162214 292567 162270 292576
rect 162228 257378 162256 292567
rect 162216 257372 162268 257378
rect 162216 257314 162268 257320
rect 164884 225752 164936 225758
rect 164884 225694 164936 225700
rect 164896 203590 164924 225694
rect 164884 203584 164936 203590
rect 164884 203526 164936 203532
rect 162124 181756 162176 181762
rect 162124 181698 162176 181704
rect 164884 181008 164936 181014
rect 164884 180950 164936 180956
rect 159364 180192 159416 180198
rect 159364 180134 159416 180140
rect 133144 179716 133196 179722
rect 133144 179658 133196 179664
rect 164424 179716 164476 179722
rect 164424 179658 164476 179664
rect 129646 177712 129702 177721
rect 129646 177647 129702 177656
rect 131026 177712 131082 177721
rect 131026 177647 131082 177656
rect 132406 177712 132462 177721
rect 132406 177647 132462 177656
rect 133156 177177 133184 179658
rect 148232 178356 148284 178362
rect 148232 178298 148284 178304
rect 133142 177168 133198 177177
rect 133142 177103 133198 177112
rect 134432 176996 134484 177002
rect 134432 176938 134484 176944
rect 134444 176769 134472 176938
rect 148244 176769 148272 178298
rect 110748 176760 110750 176769
rect 110694 176695 110750 176704
rect 114374 176760 114430 176769
rect 114374 176695 114430 176704
rect 118422 176760 118478 176769
rect 118422 176695 118478 176704
rect 124494 176760 124550 176769
rect 124494 176695 124550 176704
rect 125782 176760 125838 176769
rect 125782 176695 125838 176704
rect 127070 176760 127126 176769
rect 127070 176695 127126 176704
rect 134430 176760 134486 176769
rect 134430 176695 134486 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 135720 176656 135772 176662
rect 135720 176598 135772 176604
rect 123116 176180 123168 176186
rect 123116 176122 123168 176128
rect 109684 176044 109736 176050
rect 109684 175986 109736 175992
rect 113180 176044 113232 176050
rect 113180 175986 113232 175992
rect 98368 175918 98420 175924
rect 109406 175944 109462 175953
rect 98380 175409 98408 175918
rect 109406 175879 109462 175888
rect 98366 175400 98422 175409
rect 98366 175335 98422 175344
rect 113192 175001 113220 175986
rect 123128 175001 123156 176122
rect 128176 176112 128228 176118
rect 128176 176054 128228 176060
rect 128188 175409 128216 176054
rect 135732 175545 135760 176598
rect 158904 176248 158956 176254
rect 158904 176190 158956 176196
rect 135718 175536 135774 175545
rect 135718 175471 135774 175480
rect 158916 175409 158944 176190
rect 128174 175400 128230 175409
rect 128174 175335 128230 175344
rect 158902 175400 158958 175409
rect 158902 175335 158958 175344
rect 164436 175166 164464 179658
rect 164424 175160 164476 175166
rect 164424 175102 164476 175108
rect 113178 174992 113234 175001
rect 113178 174927 113234 174936
rect 123114 174992 123170 175001
rect 123114 174927 123170 174936
rect 164896 173874 164924 180950
rect 166276 178673 166304 400279
rect 198004 399492 198056 399498
rect 198004 399434 198056 399440
rect 170404 398880 170456 398886
rect 170404 398822 170456 398828
rect 167644 306400 167696 306406
rect 167644 306342 167696 306348
rect 166356 203856 166408 203862
rect 166356 203798 166408 203804
rect 166262 178664 166318 178673
rect 166262 178599 166318 178608
rect 166368 177342 166396 203798
rect 167656 181626 167684 306342
rect 169024 298444 169076 298450
rect 169024 298386 169076 298392
rect 169036 250578 169064 298386
rect 169024 250572 169076 250578
rect 169024 250514 169076 250520
rect 169022 237960 169078 237969
rect 169022 237895 169078 237904
rect 169036 189786 169064 237895
rect 169024 189780 169076 189786
rect 169024 189722 169076 189728
rect 169116 189236 169168 189242
rect 169116 189178 169168 189184
rect 167644 181620 167696 181626
rect 167644 181562 167696 181568
rect 167828 180940 167880 180946
rect 167828 180882 167880 180888
rect 167736 180872 167788 180878
rect 167736 180814 167788 180820
rect 166540 179648 166592 179654
rect 166540 179590 166592 179596
rect 166448 179580 166500 179586
rect 166448 179522 166500 179528
rect 166356 177336 166408 177342
rect 166356 177278 166408 177284
rect 165252 176996 165304 177002
rect 165252 176938 165304 176944
rect 165264 175234 165292 176938
rect 166264 176180 166316 176186
rect 166264 176122 166316 176128
rect 165252 175228 165304 175234
rect 165252 175170 165304 175176
rect 164884 173868 164936 173874
rect 164884 173810 164936 173816
rect 166276 169726 166304 176122
rect 166264 169720 166316 169726
rect 166264 169662 166316 169668
rect 166460 165578 166488 179522
rect 166552 168366 166580 179590
rect 166632 176928 166684 176934
rect 166632 176870 166684 176876
rect 166644 171086 166672 176870
rect 167644 176248 167696 176254
rect 167644 176190 167696 176196
rect 167090 171592 167146 171601
rect 167090 171527 167146 171536
rect 167104 171358 167132 171527
rect 167092 171352 167144 171358
rect 167092 171294 167144 171300
rect 166632 171080 166684 171086
rect 166632 171022 166684 171028
rect 166540 168360 166592 168366
rect 166540 168302 166592 168308
rect 166448 165572 166500 165578
rect 166448 165514 166500 165520
rect 167656 149054 167684 176190
rect 167748 167006 167776 180814
rect 167840 168298 167868 180882
rect 169024 178356 169076 178362
rect 169024 178298 169076 178304
rect 167920 178288 167972 178294
rect 167920 178230 167972 178236
rect 167828 168292 167880 168298
rect 167828 168234 167880 168240
rect 167736 167000 167788 167006
rect 167736 166942 167788 166948
rect 167932 165510 167960 178230
rect 167920 165504 167972 165510
rect 167920 165446 167972 165452
rect 169036 150414 169064 178298
rect 169128 160070 169156 189178
rect 169208 184952 169260 184958
rect 169208 184894 169260 184900
rect 169116 160064 169168 160070
rect 169116 160006 169168 160012
rect 169220 157350 169248 184894
rect 169300 171352 169352 171358
rect 169300 171294 169352 171300
rect 169312 160750 169340 171294
rect 169300 160744 169352 160750
rect 169300 160686 169352 160692
rect 169208 157344 169260 157350
rect 169208 157286 169260 157292
rect 169024 150408 169076 150414
rect 169024 150350 169076 150356
rect 167644 149048 167696 149054
rect 167644 148990 167696 148996
rect 167644 146328 167696 146334
rect 167644 146270 167696 146276
rect 66166 129296 66222 129305
rect 66166 129231 66222 129240
rect 66074 128072 66130 128081
rect 66074 128007 66130 128016
rect 65154 126304 65210 126313
rect 65154 126239 65210 126248
rect 65168 125662 65196 126239
rect 65156 125656 65208 125662
rect 65156 125598 65208 125604
rect 65982 102368 66038 102377
rect 65982 102303 66038 102312
rect 65996 89690 66024 102303
rect 66088 94897 66116 128007
rect 66074 94888 66130 94897
rect 66074 94823 66130 94832
rect 66180 93809 66208 129231
rect 67638 125216 67694 125225
rect 67638 125151 67694 125160
rect 67546 123584 67602 123593
rect 67546 123519 67602 123528
rect 67362 122632 67418 122641
rect 67362 122567 67418 122576
rect 66166 93800 66222 93809
rect 66166 93735 66222 93744
rect 67376 91089 67404 122567
rect 67454 120864 67510 120873
rect 67454 120799 67510 120808
rect 67362 91080 67418 91089
rect 67362 91015 67418 91024
rect 65984 89684 66036 89690
rect 65984 89626 66036 89632
rect 67468 84182 67496 120799
rect 67560 85542 67588 123519
rect 67652 93838 67680 125151
rect 166356 117360 166408 117366
rect 166356 117302 166408 117308
rect 166264 110492 166316 110498
rect 166264 110434 166316 110440
rect 67730 100736 67786 100745
rect 67730 100671 67786 100680
rect 67640 93832 67692 93838
rect 67640 93774 67692 93780
rect 67744 86970 67772 100671
rect 164884 99408 164936 99414
rect 164884 99350 164936 99356
rect 93858 94752 93914 94761
rect 93858 94687 93914 94696
rect 106646 94752 106702 94761
rect 106646 94687 106702 94696
rect 118238 94752 118294 94761
rect 118238 94687 118294 94696
rect 120630 94752 120686 94761
rect 120630 94687 120686 94696
rect 93872 93906 93900 94687
rect 106660 93974 106688 94687
rect 118252 94042 118280 94687
rect 120644 94110 120672 94687
rect 130384 94512 130436 94518
rect 130384 94454 130436 94460
rect 120632 94104 120684 94110
rect 120632 94046 120684 94052
rect 118240 94036 118292 94042
rect 118240 93978 118292 93984
rect 106648 93968 106700 93974
rect 106648 93910 106700 93916
rect 93860 93900 93912 93906
rect 93860 93842 93912 93848
rect 114374 93664 114430 93673
rect 114374 93599 114430 93608
rect 113822 93528 113878 93537
rect 113822 93463 113878 93472
rect 103426 93256 103482 93265
rect 103426 93191 103482 93200
rect 110142 93256 110198 93265
rect 113836 93226 113864 93463
rect 114388 93362 114416 93599
rect 129462 93528 129518 93537
rect 129462 93463 129518 93472
rect 114376 93356 114428 93362
rect 114376 93298 114428 93304
rect 129476 93294 129504 93463
rect 129464 93288 129516 93294
rect 129464 93230 129516 93236
rect 110142 93191 110198 93200
rect 113824 93220 113876 93226
rect 88984 92472 89036 92478
rect 74814 92440 74870 92449
rect 74814 92375 74870 92384
rect 84382 92440 84438 92449
rect 84382 92375 84438 92384
rect 88982 92440 88984 92449
rect 89036 92440 89038 92449
rect 88982 92375 89038 92384
rect 98182 92440 98238 92449
rect 98182 92375 98238 92384
rect 74828 91118 74856 92375
rect 84396 92070 84424 92375
rect 98196 92342 98224 92375
rect 98184 92336 98236 92342
rect 98184 92278 98236 92284
rect 84384 92064 84436 92070
rect 84384 92006 84436 92012
rect 100574 91760 100630 91769
rect 100574 91695 100630 91704
rect 102874 91760 102930 91769
rect 102874 91695 102930 91704
rect 97814 91352 97870 91361
rect 97814 91287 97870 91296
rect 99194 91352 99250 91361
rect 99194 91287 99250 91296
rect 85854 91216 85910 91225
rect 85854 91151 85910 91160
rect 86866 91216 86922 91225
rect 86866 91151 86922 91160
rect 88062 91216 88118 91225
rect 88062 91151 88118 91160
rect 90638 91216 90694 91225
rect 90638 91151 90694 91160
rect 92294 91216 92350 91225
rect 92294 91151 92350 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 74816 91112 74868 91118
rect 74816 91054 74868 91060
rect 85868 88262 85896 91151
rect 85856 88256 85908 88262
rect 85856 88198 85908 88204
rect 67732 86964 67784 86970
rect 67732 86906 67784 86912
rect 67548 85536 67600 85542
rect 67548 85478 67600 85484
rect 67456 84176 67508 84182
rect 67456 84118 67508 84124
rect 86880 78538 86908 91151
rect 88076 86766 88104 91151
rect 88064 86760 88116 86766
rect 88064 86702 88116 86708
rect 90652 85474 90680 91151
rect 90640 85468 90692 85474
rect 90640 85410 90692 85416
rect 92308 85338 92336 91151
rect 92296 85332 92348 85338
rect 92296 85274 92348 85280
rect 93780 81326 93808 91151
rect 93768 81320 93820 81326
rect 93768 81262 93820 81268
rect 95160 78606 95188 91151
rect 96540 82686 96568 91151
rect 96528 82680 96580 82686
rect 96528 82622 96580 82628
rect 97828 81433 97856 91287
rect 97906 91216 97962 91225
rect 97906 91151 97962 91160
rect 97814 81424 97870 81433
rect 97814 81359 97870 81368
rect 97920 80034 97948 91151
rect 99208 83978 99236 91287
rect 99286 91216 99342 91225
rect 99286 91151 99342 91160
rect 99196 83972 99248 83978
rect 99196 83914 99248 83920
rect 97908 80028 97960 80034
rect 97908 79970 97960 79976
rect 99300 78674 99328 91151
rect 100588 89622 100616 91695
rect 101954 91488 102010 91497
rect 101954 91423 102010 91432
rect 101862 91352 101918 91361
rect 101862 91287 101918 91296
rect 100666 91216 100722 91225
rect 100666 91151 100722 91160
rect 100576 89616 100628 89622
rect 100576 89558 100628 89564
rect 100680 86902 100708 91151
rect 101876 88330 101904 91287
rect 101864 88324 101916 88330
rect 101864 88266 101916 88272
rect 100668 86896 100720 86902
rect 100668 86838 100720 86844
rect 101968 85513 101996 91423
rect 102046 91216 102102 91225
rect 102046 91151 102102 91160
rect 101954 85504 102010 85513
rect 101954 85439 102010 85448
rect 102060 79898 102088 91151
rect 102888 89554 102916 91695
rect 102876 89548 102928 89554
rect 102876 89490 102928 89496
rect 103440 82793 103468 93191
rect 105910 92440 105966 92449
rect 105910 92375 105966 92384
rect 104714 91352 104770 91361
rect 104714 91287 104770 91296
rect 104728 83910 104756 91287
rect 104806 91216 104862 91225
rect 104806 91151 104862 91160
rect 104716 83904 104768 83910
rect 104716 83846 104768 83852
rect 103426 82784 103482 82793
rect 103426 82719 103482 82728
rect 104820 81297 104848 91151
rect 105924 91050 105952 92375
rect 108946 91352 109002 91361
rect 108946 91287 109002 91296
rect 106094 91216 106150 91225
rect 106094 91151 106150 91160
rect 107198 91216 107254 91225
rect 107198 91151 107254 91160
rect 108854 91216 108910 91225
rect 108854 91151 108910 91160
rect 105912 91044 105964 91050
rect 105912 90986 105964 90992
rect 106108 82822 106136 91151
rect 107212 88194 107240 91151
rect 107200 88188 107252 88194
rect 107200 88130 107252 88136
rect 108868 84046 108896 91151
rect 108856 84040 108908 84046
rect 108856 83982 108908 83988
rect 106096 82816 106148 82822
rect 106096 82758 106148 82764
rect 104806 81288 104862 81297
rect 104806 81223 104862 81232
rect 102048 79892 102100 79898
rect 102048 79834 102100 79840
rect 108960 79830 108988 91287
rect 110156 86698 110184 93191
rect 113824 93162 113876 93168
rect 118700 93152 118752 93158
rect 118700 93094 118752 93100
rect 111614 92440 111670 92449
rect 111614 92375 111670 92384
rect 115846 92440 115902 92449
rect 115846 92375 115902 92384
rect 110326 91352 110382 91361
rect 110326 91287 110382 91296
rect 110234 91216 110290 91225
rect 110234 91151 110290 91160
rect 110144 86692 110196 86698
rect 110144 86634 110196 86640
rect 108948 79824 109000 79830
rect 108948 79766 109000 79772
rect 99288 78668 99340 78674
rect 99288 78610 99340 78616
rect 95148 78600 95200 78606
rect 95148 78542 95200 78548
rect 86868 78532 86920 78538
rect 86868 78474 86920 78480
rect 110248 77246 110276 91151
rect 110236 77240 110288 77246
rect 110236 77182 110288 77188
rect 110340 77178 110368 91287
rect 110786 91216 110842 91225
rect 110786 91151 110842 91160
rect 110800 88233 110828 91151
rect 111628 90982 111656 92375
rect 115860 92206 115888 92375
rect 118712 92342 118740 93094
rect 124586 92440 124642 92449
rect 124586 92375 124642 92384
rect 125966 92440 126022 92449
rect 125966 92375 126022 92384
rect 126518 92440 126574 92449
rect 126518 92375 126574 92384
rect 118700 92336 118752 92342
rect 118700 92278 118752 92284
rect 115848 92200 115900 92206
rect 115848 92142 115900 92148
rect 121090 91896 121146 91905
rect 121090 91831 121146 91840
rect 115846 91624 115902 91633
rect 115846 91559 115902 91568
rect 113086 91352 113142 91361
rect 113086 91287 113142 91296
rect 112994 91216 113050 91225
rect 112994 91151 113050 91160
rect 111616 90976 111668 90982
rect 111616 90918 111668 90924
rect 110786 88224 110842 88233
rect 110786 88159 110842 88168
rect 113008 81394 113036 91151
rect 112996 81388 113048 81394
rect 112996 81330 113048 81336
rect 113100 78470 113128 91287
rect 115754 91216 115810 91225
rect 115754 91151 115810 91160
rect 115768 86630 115796 91151
rect 115860 89486 115888 91559
rect 117134 91352 117190 91361
rect 117134 91287 117190 91296
rect 115848 89480 115900 89486
rect 115848 89422 115900 89428
rect 117148 88126 117176 91287
rect 117226 91216 117282 91225
rect 117226 91151 117282 91160
rect 118238 91216 118294 91225
rect 118238 91151 118294 91160
rect 119986 91216 120042 91225
rect 119986 91151 120042 91160
rect 117136 88120 117188 88126
rect 117136 88062 117188 88068
rect 115756 86624 115808 86630
rect 115756 86566 115808 86572
rect 117240 82657 117268 91151
rect 118252 85406 118280 91151
rect 118240 85400 118292 85406
rect 118240 85342 118292 85348
rect 120000 83842 120028 91151
rect 121104 89729 121132 91831
rect 122746 91352 122802 91361
rect 122746 91287 122802 91296
rect 124034 91352 124090 91361
rect 124034 91287 124090 91296
rect 122654 91216 122710 91225
rect 122654 91151 122710 91160
rect 121090 89720 121146 89729
rect 121090 89655 121146 89664
rect 122668 84114 122696 91151
rect 122656 84108 122708 84114
rect 122656 84050 122708 84056
rect 119988 83836 120040 83842
rect 119988 83778 120040 83784
rect 117226 82648 117282 82657
rect 122760 82618 122788 91287
rect 122838 91216 122894 91225
rect 122838 91151 122894 91160
rect 122852 90846 122880 91151
rect 122840 90840 122892 90846
rect 122840 90782 122892 90788
rect 124048 82754 124076 91287
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 124036 82748 124088 82754
rect 124036 82690 124088 82696
rect 117226 82583 117282 82592
rect 122748 82612 122800 82618
rect 122748 82554 122800 82560
rect 124140 79762 124168 91151
rect 124600 90778 124628 92375
rect 125980 92274 126008 92375
rect 125968 92268 126020 92274
rect 125968 92210 126020 92216
rect 125414 91216 125470 91225
rect 125414 91151 125470 91160
rect 124588 90772 124640 90778
rect 124588 90714 124640 90720
rect 125428 85270 125456 91151
rect 126532 90914 126560 92375
rect 130396 92206 130424 94454
rect 151726 93664 151782 93673
rect 151726 93599 151782 93608
rect 151740 93430 151768 93599
rect 151728 93424 151780 93430
rect 151728 93366 151780 93372
rect 164896 92478 164924 99350
rect 164884 92472 164936 92478
rect 133142 92440 133198 92449
rect 133142 92375 133198 92384
rect 136086 92440 136142 92449
rect 136086 92375 136142 92384
rect 151542 92440 151598 92449
rect 151542 92375 151598 92384
rect 152094 92440 152150 92449
rect 164884 92414 164936 92420
rect 152094 92375 152150 92384
rect 133156 92342 133184 92375
rect 133144 92336 133196 92342
rect 133144 92278 133196 92284
rect 136100 92206 136128 92375
rect 130384 92200 130436 92206
rect 130384 92142 130436 92148
rect 136088 92200 136140 92206
rect 136088 92142 136140 92148
rect 132406 91624 132462 91633
rect 132406 91559 132462 91568
rect 126886 91216 126942 91225
rect 126886 91151 126942 91160
rect 128174 91216 128230 91225
rect 128174 91151 128230 91160
rect 131026 91216 131082 91225
rect 131026 91151 131082 91160
rect 126520 90908 126572 90914
rect 126520 90850 126572 90856
rect 125416 85264 125468 85270
rect 125416 85206 125468 85212
rect 126900 79966 126928 91151
rect 128188 86834 128216 91151
rect 128176 86828 128228 86834
rect 128176 86770 128228 86776
rect 131040 81258 131068 91151
rect 132420 89418 132448 91559
rect 135074 91216 135130 91225
rect 135074 91151 135130 91160
rect 132408 89412 132460 89418
rect 132408 89354 132460 89360
rect 135088 87990 135116 91151
rect 135904 91112 135956 91118
rect 135904 91054 135956 91060
rect 135076 87984 135128 87990
rect 135076 87926 135128 87932
rect 131028 81252 131080 81258
rect 131028 81194 131080 81200
rect 126888 79960 126940 79966
rect 126888 79902 126940 79908
rect 124128 79756 124180 79762
rect 124128 79698 124180 79704
rect 113088 78464 113140 78470
rect 113088 78406 113140 78412
rect 135916 78402 135944 91054
rect 151556 90710 151584 92375
rect 152108 92138 152136 92375
rect 152096 92132 152148 92138
rect 152096 92074 152148 92080
rect 151634 91216 151690 91225
rect 151634 91151 151690 91160
rect 151544 90704 151596 90710
rect 151544 90646 151596 90652
rect 151648 88058 151676 91151
rect 151636 88052 151688 88058
rect 151636 87994 151688 88000
rect 166276 83978 166304 110434
rect 166368 90982 166396 117302
rect 166448 98048 166500 98054
rect 166448 97990 166500 97996
rect 166356 90976 166408 90982
rect 166356 90918 166408 90924
rect 166460 88262 166488 97990
rect 166540 97300 166592 97306
rect 166540 97242 166592 97248
rect 166552 92313 166580 97242
rect 166538 92304 166594 92313
rect 166538 92239 166594 92248
rect 166448 88256 166500 88262
rect 166448 88198 166500 88204
rect 167656 87990 167684 146270
rect 169024 142860 169076 142866
rect 169024 142802 169076 142808
rect 167828 122868 167880 122874
rect 167828 122810 167880 122816
rect 167736 113212 167788 113218
rect 167736 113154 167788 113160
rect 167644 87984 167696 87990
rect 167644 87926 167696 87932
rect 166264 83972 166316 83978
rect 166264 83914 166316 83920
rect 167748 83910 167776 113154
rect 167840 94110 167868 122810
rect 167920 111784 167972 111790
rect 167918 111752 167920 111761
rect 167972 111752 167974 111761
rect 167918 111687 167974 111696
rect 168104 110424 168156 110430
rect 168104 110366 168156 110372
rect 168116 110129 168144 110366
rect 168102 110120 168158 110129
rect 168102 110055 168158 110064
rect 167920 108996 167972 109002
rect 167920 108938 167972 108944
rect 167932 108769 167960 108938
rect 167918 108760 167974 108769
rect 167918 108695 167974 108704
rect 167920 98116 167972 98122
rect 167920 98058 167972 98064
rect 167828 94104 167880 94110
rect 167828 94046 167880 94052
rect 167736 83904 167788 83910
rect 167736 83846 167788 83852
rect 167932 78538 167960 98058
rect 169036 92342 169064 142802
rect 169116 124228 169168 124234
rect 169116 124170 169168 124176
rect 169024 92336 169076 92342
rect 169024 92278 169076 92284
rect 169128 79762 169156 124170
rect 170416 120766 170444 398822
rect 195244 396092 195296 396098
rect 195244 396034 195296 396040
rect 191104 374672 191156 374678
rect 191104 374614 191156 374620
rect 188344 359508 188396 359514
rect 188344 359450 188396 359456
rect 184204 347064 184256 347070
rect 184204 347006 184256 347012
rect 177304 325100 177356 325106
rect 177304 325042 177356 325048
rect 173164 303068 173216 303074
rect 173164 303010 173216 303016
rect 173176 249082 173204 303010
rect 173900 271924 173952 271930
rect 173900 271866 173952 271872
rect 173164 249076 173216 249082
rect 173164 249018 173216 249024
rect 173164 229832 173216 229838
rect 173164 229774 173216 229780
rect 171784 187808 171836 187814
rect 171784 187750 171836 187756
rect 170496 178220 170548 178226
rect 170496 178162 170548 178168
rect 170508 162858 170536 178162
rect 170588 176860 170640 176866
rect 170588 176802 170640 176808
rect 170600 169658 170628 176802
rect 170588 169652 170640 169658
rect 170588 169594 170640 169600
rect 170496 162852 170548 162858
rect 170496 162794 170548 162800
rect 171796 158710 171824 187750
rect 173176 180130 173204 229774
rect 173256 189168 173308 189174
rect 173256 189110 173308 189116
rect 173164 180124 173216 180130
rect 173164 180066 173216 180072
rect 173268 160002 173296 189110
rect 173348 179512 173400 179518
rect 173348 179454 173400 179460
rect 173256 159996 173308 160002
rect 173256 159938 173308 159944
rect 171784 158704 171836 158710
rect 171784 158646 171836 158652
rect 173360 155922 173388 179454
rect 173348 155916 173400 155922
rect 173348 155858 173400 155864
rect 171784 144968 171836 144974
rect 171784 144910 171836 144916
rect 170588 132524 170640 132530
rect 170588 132466 170640 132472
rect 170496 121508 170548 121514
rect 170496 121450 170548 121456
rect 170404 120760 170456 120766
rect 170404 120702 170456 120708
rect 169208 114572 169260 114578
rect 169208 114514 169260 114520
rect 169220 88194 169248 114514
rect 170404 106344 170456 106350
rect 170404 106286 170456 106292
rect 169300 99476 169352 99482
rect 169300 99418 169352 99424
rect 169208 88188 169260 88194
rect 169208 88130 169260 88136
rect 169312 86766 169340 99418
rect 169300 86760 169352 86766
rect 169300 86702 169352 86708
rect 170416 85338 170444 106286
rect 170404 85332 170456 85338
rect 170404 85274 170456 85280
rect 170508 83842 170536 121450
rect 170600 93974 170628 132466
rect 170680 124296 170732 124302
rect 170680 124238 170732 124244
rect 170588 93968 170640 93974
rect 170588 93910 170640 93916
rect 170692 90846 170720 124238
rect 170680 90840 170732 90846
rect 170680 90782 170732 90788
rect 171796 89418 171824 144910
rect 171876 140820 171928 140826
rect 171876 140762 171928 140768
rect 171888 90778 171916 140762
rect 173256 135312 173308 135318
rect 173256 135254 173308 135260
rect 173164 128376 173216 128382
rect 173164 128318 173216 128324
rect 172060 121576 172112 121582
rect 172060 121518 172112 121524
rect 171968 109064 172020 109070
rect 171968 109006 172020 109012
rect 171876 90772 171928 90778
rect 171876 90714 171928 90720
rect 171784 89412 171836 89418
rect 171784 89354 171836 89360
rect 170496 83836 170548 83842
rect 170496 83778 170548 83784
rect 171980 82686 172008 109006
rect 172072 94042 172100 121518
rect 172060 94036 172112 94042
rect 172060 93978 172112 93984
rect 171968 82680 172020 82686
rect 171968 82622 172020 82628
rect 173176 79898 173204 128318
rect 173268 93362 173296 135254
rect 173440 120148 173492 120154
rect 173440 120090 173492 120096
rect 173348 116000 173400 116006
rect 173348 115942 173400 115948
rect 173256 93356 173308 93362
rect 173256 93298 173308 93304
rect 173164 79892 173216 79898
rect 173164 79834 173216 79840
rect 169116 79756 169168 79762
rect 169116 79698 169168 79704
rect 167920 78532 167972 78538
rect 167920 78474 167972 78480
rect 135904 78396 135956 78402
rect 135904 78338 135956 78344
rect 173360 77178 173388 115942
rect 173452 86630 173480 120090
rect 173440 86624 173492 86630
rect 173440 86566 173492 86572
rect 110328 77172 110380 77178
rect 110328 77114 110380 77120
rect 173348 77172 173400 77178
rect 173348 77114 173400 77120
rect 122840 76628 122892 76634
rect 122840 76570 122892 76576
rect 104900 75268 104952 75274
rect 104900 75210 104952 75216
rect 75920 73840 75972 73846
rect 75920 73782 75972 73788
rect 64420 72480 64472 72486
rect 64420 72422 64472 72428
rect 74540 68332 74592 68338
rect 74540 68274 74592 68280
rect 64880 61396 64932 61402
rect 64880 61338 64932 61344
rect 64892 16574 64920 61338
rect 69020 60104 69072 60110
rect 69020 60046 69072 60052
rect 67640 21412 67692 21418
rect 67640 21354 67692 21360
rect 64892 16546 65104 16574
rect 63408 11756 63460 11762
rect 63408 11698 63460 11704
rect 63224 4820 63276 4826
rect 63224 4762 63276 4768
rect 63236 480 63264 4762
rect 64328 3528 64380 3534
rect 64328 3470 64380 3476
rect 64340 480 64368 3470
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66718 2000 66774 2009
rect 66718 1935 66774 1944
rect 66732 480 66760 1935
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 21354
rect 69032 16574 69060 60046
rect 71780 58676 71832 58682
rect 71780 58618 71832 58624
rect 70400 18624 70452 18630
rect 70400 18566 70452 18572
rect 70412 16574 70440 18566
rect 71792 16574 71820 58618
rect 73160 28348 73212 28354
rect 73160 28290 73212 28296
rect 73172 16574 73200 28290
rect 74552 16574 74580 68274
rect 69032 16546 69152 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69124 480 69152 16546
rect 70308 7676 70360 7682
rect 70308 7618 70360 7624
rect 70320 480 70348 7618
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 73782
rect 98000 69692 98052 69698
rect 98000 69634 98052 69640
rect 81440 66972 81492 66978
rect 81440 66914 81492 66920
rect 78678 50280 78734 50289
rect 78678 50215 78734 50224
rect 77300 19984 77352 19990
rect 77300 19926 77352 19932
rect 77312 16574 77340 19926
rect 78692 16574 78720 50215
rect 81452 16574 81480 66914
rect 85580 65544 85632 65550
rect 85580 65486 85632 65492
rect 84200 20052 84252 20058
rect 84200 19994 84252 20000
rect 82820 18692 82872 18698
rect 82820 18634 82872 18640
rect 82832 16574 82860 18634
rect 77312 16546 77432 16574
rect 78692 16546 79272 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77404 480 77432 16546
rect 78128 10328 78180 10334
rect 78128 10270 78180 10276
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 10270
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80888 13184 80940 13190
rect 80888 13126 80940 13132
rect 80900 480 80928 13126
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 19994
rect 85592 6914 85620 65486
rect 87604 64252 87656 64258
rect 87604 64194 87656 64200
rect 85672 57316 85724 57322
rect 85672 57258 85724 57264
rect 85684 16574 85712 57258
rect 85684 16546 86448 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 87512 14544 87564 14550
rect 87512 14486 87564 14492
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 14486
rect 87616 3534 87644 64194
rect 88340 62892 88392 62898
rect 88340 62834 88392 62840
rect 88352 16574 88380 62834
rect 92480 61464 92532 61470
rect 92480 61406 92532 61412
rect 89720 21480 89772 21486
rect 89720 21422 89772 21428
rect 89732 16574 89760 21422
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 87604 3528 87656 3534
rect 87604 3470 87656 3476
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 4888 91612 4894
rect 91560 4830 91612 4836
rect 91572 480 91600 4830
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 61406
rect 96620 49088 96672 49094
rect 96620 49030 96672 49036
rect 93860 47660 93912 47666
rect 93860 47602 93912 47608
rect 93872 16574 93900 47602
rect 95240 31204 95292 31210
rect 95240 31146 95292 31152
rect 95252 16574 95280 31146
rect 96632 16574 96660 49030
rect 98012 16574 98040 69634
rect 100760 40792 100812 40798
rect 100760 40734 100812 40740
rect 93872 16546 93992 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 93964 480 93992 16546
rect 94688 13116 94740 13122
rect 94688 13058 94740 13064
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 13058
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99840 3392 99892 3398
rect 99840 3334 99892 3340
rect 99852 480 99880 3334
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 40734
rect 103520 35284 103572 35290
rect 103520 35226 103572 35232
rect 103532 16574 103560 35226
rect 104912 16574 104940 75210
rect 110420 69760 110472 69766
rect 110420 69702 110472 69708
rect 107660 53168 107712 53174
rect 107660 53110 107712 53116
rect 106280 46300 106332 46306
rect 106280 46242 106332 46248
rect 106292 16574 106320 46242
rect 107672 16574 107700 53110
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102140 15972 102192 15978
rect 102140 15914 102192 15920
rect 102152 3534 102180 15914
rect 102232 9036 102284 9042
rect 102232 8978 102284 8984
rect 102140 3528 102192 3534
rect 102140 3470 102192 3476
rect 102244 480 102272 8978
rect 103336 3528 103388 3534
rect 103336 3470 103388 3476
rect 103428 3528 103480 3534
rect 103428 3470 103480 3476
rect 103348 480 103376 3470
rect 103440 3398 103468 3470
rect 103428 3392 103480 3398
rect 103428 3334 103480 3340
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 110432 6914 110460 69702
rect 113180 60172 113232 60178
rect 113180 60114 113232 60120
rect 111800 58744 111852 58750
rect 111800 58686 111852 58692
rect 110512 39432 110564 39438
rect 110512 39374 110564 39380
rect 110524 16574 110552 39374
rect 111812 16574 111840 58686
rect 113192 16574 113220 60114
rect 118700 51808 118752 51814
rect 118700 51750 118752 51756
rect 117320 46368 117372 46374
rect 117320 46310 117372 46316
rect 114560 29708 114612 29714
rect 114560 29650 114612 29656
rect 114572 16574 114600 29650
rect 115940 22840 115992 22846
rect 115940 22782 115992 22788
rect 115952 16574 115980 22782
rect 110524 16546 111656 16574
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 110432 6886 110552 6914
rect 109316 2100 109368 2106
rect 109316 2042 109368 2048
rect 109328 480 109356 2042
rect 110524 480 110552 6886
rect 111628 480 111656 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 46310
rect 118712 16574 118740 51750
rect 121460 31136 121512 31142
rect 121460 31078 121512 31084
rect 120078 25528 120134 25537
rect 120078 25463 120134 25472
rect 120092 16574 120120 25463
rect 121472 16574 121500 31078
rect 122852 16574 122880 76570
rect 124220 56024 124272 56030
rect 124220 55966 124272 55972
rect 124232 16574 124260 55966
rect 118712 16546 118832 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 118804 480 118832 16546
rect 119894 14512 119950 14521
rect 119894 14447 119950 14456
rect 119908 480 119936 14447
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 164424 14476 164476 14482
rect 164424 14418 164476 14424
rect 136456 6316 136508 6322
rect 136456 6258 136508 6264
rect 132960 6248 133012 6254
rect 132960 6190 133012 6196
rect 125876 3664 125928 3670
rect 125876 3606 125928 3612
rect 125888 480 125916 3606
rect 129372 3596 129424 3602
rect 129372 3538 129424 3544
rect 129384 480 129412 3538
rect 132972 480 133000 6190
rect 136468 480 136496 6258
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 14418
rect 173912 3670 173940 271866
rect 175924 187128 175976 187134
rect 175924 187070 175976 187076
rect 174544 184476 174596 184482
rect 174544 184418 174596 184424
rect 174556 32502 174584 184418
rect 174636 137284 174688 137290
rect 174636 137226 174688 137232
rect 174648 92177 174676 137226
rect 174728 107704 174780 107710
rect 174728 107646 174780 107652
rect 174740 93906 174768 107646
rect 175936 102814 175964 187070
rect 176016 143608 176068 143614
rect 176016 143550 176068 143556
rect 175924 102808 175976 102814
rect 175924 102750 175976 102756
rect 174728 93900 174780 93906
rect 174728 93842 174780 93848
rect 176028 93294 176056 143550
rect 176108 125656 176160 125662
rect 176108 125598 176160 125604
rect 176016 93288 176068 93294
rect 176016 93230 176068 93236
rect 174634 92168 174690 92177
rect 174634 92103 174690 92112
rect 176120 85270 176148 125598
rect 176200 116068 176252 116074
rect 176200 116010 176252 116016
rect 176108 85264 176160 85270
rect 176108 85206 176160 85212
rect 176212 79830 176240 116010
rect 176200 79824 176252 79830
rect 176200 79766 176252 79772
rect 177316 53242 177344 325042
rect 180064 303952 180116 303958
rect 180064 303894 180116 303900
rect 178682 299568 178738 299577
rect 178682 299503 178738 299512
rect 178696 251938 178724 299503
rect 178776 291372 178828 291378
rect 178776 291314 178828 291320
rect 178684 251932 178736 251938
rect 178684 251874 178736 251880
rect 178684 238332 178736 238338
rect 178684 238274 178736 238280
rect 177488 148368 177540 148374
rect 177488 148310 177540 148316
rect 177396 122936 177448 122942
rect 177396 122878 177448 122884
rect 177408 82618 177436 122878
rect 177500 111790 177528 148310
rect 177580 117428 177632 117434
rect 177580 117370 177632 117376
rect 177488 111784 177540 111790
rect 177488 111726 177540 111732
rect 177488 106412 177540 106418
rect 177488 106354 177540 106360
rect 177396 82612 177448 82618
rect 177396 82554 177448 82560
rect 177500 81326 177528 106354
rect 177592 86698 177620 117370
rect 178696 92342 178724 238274
rect 178788 178906 178816 291314
rect 180076 229838 180104 303894
rect 182180 240780 182232 240786
rect 182180 240722 182232 240728
rect 180064 229832 180116 229838
rect 180064 229774 180116 229780
rect 178776 178900 178828 178906
rect 178776 178842 178828 178848
rect 180062 178664 180118 178673
rect 180062 178599 180118 178608
rect 178868 140072 178920 140078
rect 178868 140014 178920 140020
rect 178776 120216 178828 120222
rect 178776 120158 178828 120164
rect 178684 92336 178736 92342
rect 178684 92278 178736 92284
rect 178788 88126 178816 120158
rect 178880 110430 178908 140014
rect 178960 118720 179012 118726
rect 178960 118662 179012 118668
rect 178868 110424 178920 110430
rect 178868 110366 178920 110372
rect 178868 107772 178920 107778
rect 178868 107714 178920 107720
rect 178776 88120 178828 88126
rect 178776 88062 178828 88068
rect 177580 86692 177632 86698
rect 177580 86634 177632 86640
rect 177488 81320 177540 81326
rect 177488 81262 177540 81268
rect 178880 78606 178908 107714
rect 178972 89486 179000 118662
rect 178960 89480 179012 89486
rect 178960 89422 179012 89428
rect 178868 78600 178920 78606
rect 178868 78542 178920 78548
rect 177304 53236 177356 53242
rect 177304 53178 177356 53184
rect 174544 32496 174596 32502
rect 174544 32438 174596 32444
rect 180076 17270 180104 178599
rect 180248 151836 180300 151842
rect 180248 151778 180300 151784
rect 180156 132592 180208 132598
rect 180156 132534 180208 132540
rect 180168 84046 180196 132534
rect 180260 109002 180288 151778
rect 181444 133952 181496 133958
rect 181444 133894 181496 133900
rect 180340 125724 180392 125730
rect 180340 125666 180392 125672
rect 180248 108996 180300 109002
rect 180248 108938 180300 108944
rect 180352 90914 180380 125666
rect 180340 90908 180392 90914
rect 180340 90850 180392 90856
rect 180156 84040 180208 84046
rect 180156 83982 180208 83988
rect 181456 77246 181484 133894
rect 181536 111852 181588 111858
rect 181536 111794 181588 111800
rect 181548 88330 181576 111794
rect 181536 88324 181588 88330
rect 181536 88266 181588 88272
rect 181444 77240 181496 77246
rect 181444 77182 181496 77188
rect 182192 69601 182220 240722
rect 182914 70272 182970 70281
rect 182914 70207 182970 70216
rect 182928 69601 182956 70207
rect 182178 69592 182234 69601
rect 182178 69527 182234 69536
rect 182914 69592 182970 69601
rect 182914 69527 182970 69536
rect 180064 17264 180116 17270
rect 180064 17206 180116 17212
rect 184216 4962 184244 347006
rect 186964 345704 187016 345710
rect 186964 345646 187016 345652
rect 184296 135380 184348 135386
rect 184296 135322 184348 135328
rect 184308 78470 184336 135322
rect 185584 118788 185636 118794
rect 185584 118730 185636 118736
rect 185596 93226 185624 118730
rect 185584 93220 185636 93226
rect 185584 93162 185636 93168
rect 184296 78464 184348 78470
rect 184296 78406 184348 78412
rect 186976 9654 187004 345646
rect 187056 224324 187108 224330
rect 187056 224266 187108 224272
rect 187068 183122 187096 224266
rect 187056 183116 187108 183122
rect 187056 183058 187108 183064
rect 187056 153264 187108 153270
rect 187056 153206 187108 153212
rect 187068 93430 187096 153206
rect 187056 93424 187108 93430
rect 187056 93366 187108 93372
rect 188356 13258 188384 359450
rect 188434 295352 188490 295361
rect 188434 295287 188490 295296
rect 188448 96422 188476 295287
rect 189724 151904 189776 151910
rect 189724 151846 189776 151852
rect 188528 111920 188580 111926
rect 188528 111862 188580 111868
rect 188436 96416 188488 96422
rect 188436 96358 188488 96364
rect 188540 86902 188568 111862
rect 189736 92138 189764 151846
rect 189724 92132 189776 92138
rect 189724 92074 189776 92080
rect 188528 86896 188580 86902
rect 188528 86838 188580 86844
rect 191116 20670 191144 374614
rect 192484 180192 192536 180198
rect 192484 180134 192536 180140
rect 191196 147688 191248 147694
rect 191196 147630 191248 147636
rect 191208 92206 191236 147630
rect 192496 92478 192524 180134
rect 193864 131164 193916 131170
rect 193864 131106 193916 131112
rect 192576 105052 192628 105058
rect 192576 104994 192628 105000
rect 192588 93809 192616 104994
rect 192574 93800 192630 93809
rect 192574 93735 192630 93744
rect 192484 92472 192536 92478
rect 192484 92414 192536 92420
rect 191196 92200 191248 92206
rect 191196 92142 191248 92148
rect 193876 91050 193904 131106
rect 193864 91044 193916 91050
rect 193864 90986 193916 90992
rect 191104 20664 191156 20670
rect 191104 20606 191156 20612
rect 195256 19242 195284 396034
rect 196624 351280 196676 351286
rect 196624 351222 196676 351228
rect 195336 265056 195388 265062
rect 195336 264998 195388 265004
rect 195348 93770 195376 264998
rect 195428 142180 195480 142186
rect 195428 142122 195480 142128
rect 195336 93764 195388 93770
rect 195336 93706 195388 93712
rect 195440 92274 195468 142122
rect 195428 92268 195480 92274
rect 195428 92210 195480 92216
rect 196636 28966 196664 351222
rect 196716 248464 196768 248470
rect 196716 248406 196768 248412
rect 196728 95130 196756 248406
rect 196808 145036 196860 145042
rect 196808 144978 196860 144984
rect 196716 95124 196768 95130
rect 196716 95066 196768 95072
rect 196820 81258 196848 144978
rect 198016 87650 198044 399434
rect 215944 397588 215996 397594
rect 215944 397530 215996 397536
rect 206284 394732 206336 394738
rect 206284 394674 206336 394680
rect 204904 381540 204956 381546
rect 204904 381482 204956 381488
rect 202144 362228 202196 362234
rect 202144 362170 202196 362176
rect 199384 292800 199436 292806
rect 199384 292742 199436 292748
rect 198096 289196 198148 289202
rect 198096 289138 198148 289144
rect 198108 180198 198136 289138
rect 199396 181694 199424 292742
rect 200856 273284 200908 273290
rect 200856 273226 200908 273232
rect 200868 181762 200896 273226
rect 200764 181756 200816 181762
rect 200764 181698 200816 181704
rect 200856 181756 200908 181762
rect 200856 181698 200908 181704
rect 199384 181688 199436 181694
rect 199384 181630 199436 181636
rect 199474 181384 199530 181393
rect 199474 181319 199530 181328
rect 198096 180192 198148 180198
rect 198096 180134 198148 180140
rect 198188 179444 198240 179450
rect 198188 179386 198240 179392
rect 198200 164218 198228 179386
rect 198188 164212 198240 164218
rect 198188 164154 198240 164160
rect 198096 153332 198148 153338
rect 198096 153274 198148 153280
rect 198108 90710 198136 153274
rect 198188 113280 198240 113286
rect 198188 113222 198240 113228
rect 198096 90704 198148 90710
rect 198096 90646 198148 90652
rect 198200 89554 198228 113222
rect 199384 103556 199436 103562
rect 199384 103498 199436 103504
rect 199396 93838 199424 103498
rect 199384 93832 199436 93838
rect 199488 93809 199516 181319
rect 199384 93774 199436 93780
rect 199474 93800 199530 93809
rect 199474 93735 199530 93744
rect 198188 89548 198240 89554
rect 198188 89490 198240 89496
rect 198096 89004 198148 89010
rect 198096 88946 198148 88952
rect 198004 87644 198056 87650
rect 198004 87586 198056 87592
rect 196808 81252 196860 81258
rect 196808 81194 196860 81200
rect 196624 28960 196676 28966
rect 196624 28902 196676 28908
rect 195244 19236 195296 19242
rect 195244 19178 195296 19184
rect 188344 13252 188396 13258
rect 188344 13194 188396 13200
rect 186964 9648 187016 9654
rect 186964 9590 187016 9596
rect 184204 4956 184256 4962
rect 184204 4898 184256 4904
rect 173900 3664 173952 3670
rect 173900 3606 173952 3612
rect 198108 3534 198136 88946
rect 200776 29782 200804 181698
rect 200856 102196 200908 102202
rect 200856 102138 200908 102144
rect 200868 85542 200896 102138
rect 200856 85536 200908 85542
rect 200856 85478 200908 85484
rect 200764 29776 200816 29782
rect 200764 29718 200816 29724
rect 202156 7750 202184 362170
rect 203524 298308 203576 298314
rect 203524 298250 203576 298256
rect 203536 191418 203564 298250
rect 203524 191412 203576 191418
rect 203524 191354 203576 191360
rect 202236 181552 202288 181558
rect 202236 181494 202288 181500
rect 202248 92410 202276 181494
rect 203614 180160 203670 180169
rect 203614 180095 203670 180104
rect 203524 120760 203576 120766
rect 203524 120702 203576 120708
rect 202328 103624 202380 103630
rect 202328 103566 202380 103572
rect 202236 92404 202288 92410
rect 202236 92346 202288 92352
rect 202340 75886 202368 103566
rect 202328 75880 202380 75886
rect 202328 75822 202380 75828
rect 203536 21554 203564 120702
rect 203628 95062 203656 180095
rect 203708 100768 203760 100774
rect 203708 100710 203760 100716
rect 203616 95056 203668 95062
rect 203616 94998 203668 95004
rect 203720 92070 203748 100710
rect 203708 92064 203760 92070
rect 203708 92006 203760 92012
rect 204916 29850 204944 381482
rect 205088 104984 205140 104990
rect 205088 104926 205140 104932
rect 204996 95260 205048 95266
rect 204996 95202 205048 95208
rect 205008 78402 205036 95202
rect 205100 94897 205128 104926
rect 205086 94888 205142 94897
rect 205086 94823 205142 94832
rect 204996 78396 205048 78402
rect 204996 78338 205048 78344
rect 204904 29844 204956 29850
rect 204904 29786 204956 29792
rect 206296 26994 206324 394674
rect 214564 326460 214616 326466
rect 214564 326402 214616 326408
rect 210424 303884 210476 303890
rect 210424 303826 210476 303832
rect 209134 301472 209190 301481
rect 209134 301407 209190 301416
rect 206376 278860 206428 278866
rect 206376 278802 206428 278808
rect 206388 177410 206416 278802
rect 209044 214668 209096 214674
rect 209044 214610 209096 214616
rect 206376 177404 206428 177410
rect 206376 177346 206428 177352
rect 206376 175976 206428 175982
rect 206376 175918 206428 175924
rect 206388 155854 206416 175918
rect 206376 155848 206428 155854
rect 206376 155790 206428 155796
rect 206376 140888 206428 140894
rect 206376 140830 206428 140836
rect 206388 82754 206416 140830
rect 207664 128444 207716 128450
rect 207664 128386 207716 128392
rect 206468 109132 206520 109138
rect 206468 109074 206520 109080
rect 206376 82748 206428 82754
rect 206376 82690 206428 82696
rect 206480 80034 206508 109074
rect 206468 80028 206520 80034
rect 206468 79970 206520 79976
rect 207676 78674 207704 128386
rect 207756 110560 207808 110566
rect 207756 110502 207808 110508
rect 207768 89622 207796 110502
rect 209056 95198 209084 214610
rect 209148 195430 209176 301407
rect 209136 195424 209188 195430
rect 209136 195366 209188 195372
rect 209136 187740 209188 187746
rect 209136 187682 209188 187688
rect 209148 173806 209176 187682
rect 210436 184482 210464 303826
rect 211804 298376 211856 298382
rect 211804 298318 211856 298324
rect 211816 186969 211844 298318
rect 213276 295520 213328 295526
rect 213276 295462 213328 295468
rect 213182 294400 213238 294409
rect 213182 294335 213238 294344
rect 211896 195492 211948 195498
rect 211896 195434 211948 195440
rect 211802 186960 211858 186969
rect 211802 186895 211858 186904
rect 210424 184476 210476 184482
rect 210424 184418 210476 184424
rect 209320 183592 209372 183598
rect 209320 183534 209372 183540
rect 209228 176044 209280 176050
rect 209228 175986 209280 175992
rect 209136 173800 209188 173806
rect 209136 173742 209188 173748
rect 209240 164150 209268 175986
rect 209332 172514 209360 183534
rect 211804 182232 211856 182238
rect 211804 182174 211856 182180
rect 209320 172508 209372 172514
rect 209320 172450 209372 172456
rect 211816 166938 211844 182174
rect 211908 177478 211936 195434
rect 211988 178152 212040 178158
rect 211988 178094 212040 178100
rect 211896 177472 211948 177478
rect 211896 177414 211948 177420
rect 212000 171018 212028 178094
rect 211988 171012 212040 171018
rect 211988 170954 212040 170960
rect 211804 166932 211856 166938
rect 211804 166874 211856 166880
rect 209228 164144 209280 164150
rect 209228 164086 209280 164092
rect 211804 152448 211856 152454
rect 211804 152390 211856 152396
rect 210424 143676 210476 143682
rect 210424 143618 210476 143624
rect 209136 139460 209188 139466
rect 209136 139402 209188 139408
rect 209044 95192 209096 95198
rect 209044 95134 209096 95140
rect 207756 89616 207808 89622
rect 207756 89558 207808 89564
rect 209148 84114 209176 139402
rect 209228 114640 209280 114646
rect 209228 114582 209280 114588
rect 209136 84108 209188 84114
rect 209136 84050 209188 84056
rect 209240 82822 209268 114582
rect 210436 86834 210464 143618
rect 210516 118856 210568 118862
rect 210516 118798 210568 118804
rect 210424 86828 210476 86834
rect 210424 86770 210476 86776
rect 209228 82816 209280 82822
rect 209228 82758 209280 82764
rect 210528 81394 210556 118798
rect 210608 96688 210660 96694
rect 210608 96630 210660 96636
rect 210620 89690 210648 96630
rect 210608 89684 210660 89690
rect 210608 89626 210660 89632
rect 211816 88058 211844 152390
rect 213196 95033 213224 294335
rect 213288 177313 213316 295462
rect 214576 178838 214604 326402
rect 214656 305108 214708 305114
rect 214656 305050 214708 305056
rect 214668 181558 214696 305050
rect 214748 190528 214800 190534
rect 214748 190470 214800 190476
rect 214656 181552 214708 181558
rect 214656 181494 214708 181500
rect 214564 178832 214616 178838
rect 214564 178774 214616 178780
rect 214656 178084 214708 178090
rect 214656 178026 214708 178032
rect 213274 177304 213330 177313
rect 213274 177239 213330 177248
rect 214564 176792 214616 176798
rect 214564 176734 214616 176740
rect 213368 176724 213420 176730
rect 213368 176666 213420 176672
rect 213380 158137 213408 176666
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175817 213960 176598
rect 214104 176112 214156 176118
rect 214104 176054 214156 176060
rect 213918 175808 213974 175817
rect 213918 175743 213974 175752
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175137 213960 175170
rect 214012 175160 214064 175166
rect 213918 175128 213974 175137
rect 214012 175102 214064 175108
rect 213918 175063 213974 175072
rect 214024 174729 214052 175102
rect 214010 174720 214066 174729
rect 214010 174655 214066 174664
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173777 213960 173810
rect 214012 173800 214064 173806
rect 213918 173768 213974 173777
rect 214012 173742 214064 173748
rect 213918 173703 213974 173712
rect 214024 173369 214052 173742
rect 214010 173360 214066 173369
rect 214010 173295 214066 173304
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172417 213960 172450
rect 213918 172408 213974 172417
rect 213918 172343 213974 172352
rect 214116 172009 214144 176054
rect 214102 172000 214158 172009
rect 214102 171935 214158 171944
rect 213920 171080 213972 171086
rect 213920 171022 213972 171028
rect 213932 170785 213960 171022
rect 214012 171012 214064 171018
rect 214012 170954 214064 170960
rect 214024 170921 214052 170954
rect 214010 170912 214066 170921
rect 214010 170847 214066 170856
rect 213918 170776 213974 170785
rect 213918 170711 213974 170720
rect 214012 169720 214064 169726
rect 213918 169688 213974 169697
rect 214012 169662 214064 169668
rect 213918 169623 213920 169632
rect 213972 169623 213974 169632
rect 213920 169594 213972 169600
rect 214024 169425 214052 169662
rect 214010 169416 214066 169425
rect 214010 169351 214066 169360
rect 214012 168360 214064 168366
rect 213918 168328 213974 168337
rect 214012 168302 214064 168308
rect 213918 168263 213920 168272
rect 213972 168263 213974 168272
rect 213920 168234 213972 168240
rect 214024 168065 214052 168302
rect 214010 168056 214066 168065
rect 214010 167991 214066 168000
rect 213920 167000 213972 167006
rect 213920 166942 213972 166948
rect 214102 166968 214158 166977
rect 213932 166161 213960 166942
rect 214102 166903 214104 166912
rect 214156 166903 214158 166912
rect 214104 166874 214156 166880
rect 213918 166152 213974 166161
rect 213918 166087 213974 166096
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165345 213960 165514
rect 214012 165504 214064 165510
rect 214012 165446 214064 165452
rect 213918 165336 213974 165345
rect 213918 165271 213974 165280
rect 214024 164801 214052 165446
rect 214010 164792 214066 164801
rect 214010 164727 214066 164736
rect 214012 164212 214064 164218
rect 214012 164154 214064 164160
rect 213920 164144 213972 164150
rect 213918 164112 213920 164121
rect 213972 164112 213974 164121
rect 213918 164047 213974 164056
rect 214024 163441 214052 164154
rect 214010 163432 214066 163441
rect 214010 163367 214066 163376
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162081 213960 162794
rect 214576 162761 214604 176734
rect 214668 166705 214696 178026
rect 214760 173894 214788 190470
rect 214760 173866 214880 173894
rect 214654 166696 214710 166705
rect 214654 166631 214710 166640
rect 214852 164234 214880 173866
rect 214760 164206 214880 164234
rect 214562 162752 214618 162761
rect 214562 162687 214618 162696
rect 213918 162072 213974 162081
rect 213918 162007 213974 162016
rect 214760 161265 214788 164206
rect 214746 161256 214802 161265
rect 214746 161191 214802 161200
rect 214564 160744 214616 160750
rect 214564 160686 214616 160692
rect 213920 160064 213972 160070
rect 213918 160032 213920 160041
rect 213972 160032 213974 160041
rect 213918 159967 213974 159976
rect 214012 159996 214064 160002
rect 214012 159938 214064 159944
rect 214024 159497 214052 159938
rect 214010 159488 214066 159497
rect 214010 159423 214066 159432
rect 213920 158704 213972 158710
rect 213918 158672 213920 158681
rect 213972 158672 213974 158681
rect 213918 158607 213974 158616
rect 213366 158128 213422 158137
rect 213366 158063 213422 158072
rect 214010 157992 214066 158001
rect 214010 157927 214066 157936
rect 213920 157344 213972 157350
rect 214024 157321 214052 157927
rect 213920 157286 213972 157292
rect 214010 157312 214066 157321
rect 213932 156913 213960 157286
rect 214010 157247 214066 157256
rect 213918 156904 213974 156913
rect 213918 156839 213974 156848
rect 213918 155952 213974 155961
rect 213918 155887 213974 155896
rect 214012 155916 214064 155922
rect 213932 155854 213960 155887
rect 214012 155858 214064 155864
rect 213920 155848 213972 155854
rect 213920 155790 213972 155796
rect 214024 155553 214052 155858
rect 214010 155544 214066 155553
rect 214010 155479 214066 155488
rect 214010 153912 214066 153921
rect 214010 153847 214066 153856
rect 213918 153504 213974 153513
rect 213918 153439 213974 153448
rect 213932 153270 213960 153439
rect 214024 153338 214052 153847
rect 214012 153332 214064 153338
rect 214012 153274 214064 153280
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 213918 152688 213974 152697
rect 213918 152623 213974 152632
rect 213932 152454 213960 152623
rect 213920 152448 213972 152454
rect 213920 152390 213972 152396
rect 214010 152280 214066 152289
rect 214010 152215 214066 152224
rect 213918 152008 213974 152017
rect 213918 151943 213974 151952
rect 213932 151842 213960 151943
rect 214024 151910 214052 152215
rect 214012 151904 214064 151910
rect 214012 151846 214064 151852
rect 213920 151836 213972 151842
rect 213920 151778 213972 151784
rect 214010 150648 214066 150657
rect 214010 150583 214066 150592
rect 213920 150408 213972 150414
rect 213920 150350 213972 150356
rect 213932 150113 213960 150350
rect 213918 150104 213974 150113
rect 213918 150039 213974 150048
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148753 213960 148990
rect 213918 148744 213974 148753
rect 213918 148679 213974 148688
rect 214024 148374 214052 150583
rect 214576 149569 214604 160686
rect 214654 150784 214710 150793
rect 214654 150719 214710 150728
rect 214562 149560 214618 149569
rect 214562 149495 214618 149504
rect 214012 148368 214064 148374
rect 214012 148310 214064 148316
rect 213918 148064 213974 148073
rect 213918 147999 213974 148008
rect 213932 147694 213960 147999
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 213918 146704 213974 146713
rect 213918 146639 213974 146648
rect 213932 146334 213960 146639
rect 214102 146432 214158 146441
rect 214102 146367 214158 146376
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 214010 145344 214066 145353
rect 214010 145279 214066 145288
rect 213920 145036 213972 145042
rect 213920 144978 213972 144984
rect 213932 144945 213960 144978
rect 214024 144974 214052 145279
rect 214012 144968 214064 144974
rect 213918 144936 213974 144945
rect 214012 144910 214064 144916
rect 213918 144871 213974 144880
rect 213918 143984 213974 143993
rect 213918 143919 213974 143928
rect 213932 143614 213960 143919
rect 214012 143676 214064 143682
rect 214012 143618 214064 143624
rect 213920 143608 213972 143614
rect 214024 143585 214052 143618
rect 213920 143550 213972 143556
rect 214010 143576 214066 143585
rect 214010 143511 214066 143520
rect 214116 142866 214144 146367
rect 214104 142860 214156 142866
rect 214104 142802 214156 142808
rect 213274 142760 213330 142769
rect 213274 142695 213330 142704
rect 213182 95024 213238 95033
rect 213182 94959 213238 94968
rect 211804 88052 211856 88058
rect 211804 87994 211856 88000
rect 210516 81388 210568 81394
rect 210516 81330 210568 81336
rect 213288 79966 213316 142695
rect 213918 142216 213974 142225
rect 213918 142151 213920 142160
rect 213972 142151 213974 142160
rect 213920 142122 213972 142128
rect 214010 141400 214066 141409
rect 214010 141335 214066 141344
rect 213918 140992 213974 141001
rect 213918 140927 213974 140936
rect 213932 140894 213960 140927
rect 213920 140888 213972 140894
rect 213920 140830 213972 140836
rect 214024 140826 214052 141335
rect 214012 140820 214064 140826
rect 214012 140762 214064 140768
rect 214668 140078 214696 150719
rect 214656 140072 214708 140078
rect 213918 140040 213974 140049
rect 214656 140014 214708 140020
rect 213918 139975 213974 139984
rect 213932 139466 213960 139975
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 213918 138816 213974 138825
rect 213918 138751 213974 138760
rect 213366 138136 213422 138145
rect 213366 138071 213422 138080
rect 213380 85406 213408 138071
rect 213932 137290 213960 138751
rect 213920 137284 213972 137290
rect 213920 137226 213972 137232
rect 214562 136776 214618 136785
rect 214562 136711 214618 136720
rect 214010 136096 214066 136105
rect 214010 136031 214066 136040
rect 213918 135416 213974 135425
rect 213918 135351 213920 135360
rect 213972 135351 213974 135360
rect 213920 135322 213972 135328
rect 214024 135318 214052 136031
rect 214012 135312 214064 135318
rect 214012 135254 214064 135260
rect 213918 134056 213974 134065
rect 213918 133991 213974 134000
rect 213932 133958 213960 133991
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 214010 132832 214066 132841
rect 214010 132767 214066 132776
rect 214024 132598 214052 132767
rect 214012 132592 214064 132598
rect 213918 132560 213974 132569
rect 214012 132534 214064 132540
rect 213918 132495 213920 132504
rect 213972 132495 213974 132504
rect 213920 132466 213972 132472
rect 213918 131472 213974 131481
rect 213918 131407 213974 131416
rect 213932 131170 213960 131407
rect 213920 131164 213972 131170
rect 213920 131106 213972 131112
rect 214010 128888 214066 128897
rect 214010 128823 214066 128832
rect 213918 128480 213974 128489
rect 213918 128415 213920 128424
rect 213972 128415 213974 128424
rect 213920 128386 213972 128392
rect 214024 128382 214052 128823
rect 214012 128376 214064 128382
rect 214012 128318 214064 128324
rect 214010 126168 214066 126177
rect 214010 126103 214066 126112
rect 213918 125760 213974 125769
rect 214024 125730 214052 126103
rect 213918 125695 213974 125704
rect 214012 125724 214064 125730
rect 213932 125662 213960 125695
rect 214012 125666 214064 125672
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214010 124808 214066 124817
rect 214010 124743 214066 124752
rect 213918 124400 213974 124409
rect 213918 124335 213974 124344
rect 213932 124302 213960 124335
rect 213920 124296 213972 124302
rect 213920 124238 213972 124244
rect 214024 124234 214052 124743
rect 214012 124228 214064 124234
rect 214012 124170 214064 124176
rect 214010 123584 214066 123593
rect 214010 123519 214066 123528
rect 214024 122942 214052 123519
rect 214012 122936 214064 122942
rect 213918 122904 213974 122913
rect 214012 122878 214064 122884
rect 213918 122839 213920 122848
rect 213972 122839 213974 122848
rect 213920 122810 213972 122816
rect 214010 122224 214066 122233
rect 214010 122159 214066 122168
rect 213918 121816 213974 121825
rect 213918 121751 213974 121760
rect 213932 121582 213960 121751
rect 213920 121576 213972 121582
rect 213920 121518 213972 121524
rect 214024 121514 214052 122159
rect 214012 121508 214064 121514
rect 214012 121450 214064 121456
rect 214010 120864 214066 120873
rect 214010 120799 214066 120808
rect 214024 120222 214052 120799
rect 214012 120216 214064 120222
rect 213918 120184 213974 120193
rect 214012 120158 214064 120164
rect 213918 120119 213920 120128
rect 213972 120119 213974 120128
rect 213920 120090 213972 120096
rect 214010 119640 214066 119649
rect 214010 119575 214066 119584
rect 213918 118960 213974 118969
rect 213918 118895 213974 118904
rect 213932 118794 213960 118895
rect 213920 118788 213972 118794
rect 213920 118730 213972 118736
rect 214024 118726 214052 119575
rect 214104 118856 214156 118862
rect 214102 118824 214104 118833
rect 214156 118824 214158 118833
rect 214102 118759 214158 118768
rect 214012 118720 214064 118726
rect 214012 118662 214064 118668
rect 214010 117600 214066 117609
rect 214010 117535 214066 117544
rect 213920 117428 213972 117434
rect 213920 117370 213972 117376
rect 213932 117337 213960 117370
rect 214024 117366 214052 117535
rect 214012 117360 214064 117366
rect 213918 117328 213974 117337
rect 214012 117302 214064 117308
rect 213918 117263 213974 117272
rect 214010 116240 214066 116249
rect 214010 116175 214066 116184
rect 213920 116068 213972 116074
rect 213920 116010 213972 116016
rect 213932 115977 213960 116010
rect 214024 116006 214052 116175
rect 214012 116000 214064 116006
rect 213918 115968 213974 115977
rect 214012 115942 214064 115948
rect 213918 115903 213974 115912
rect 214010 115016 214066 115025
rect 214010 114951 214066 114960
rect 213920 114640 213972 114646
rect 213918 114608 213920 114617
rect 213972 114608 213974 114617
rect 214024 114578 214052 114951
rect 213918 114543 213974 114552
rect 214012 114572 214064 114578
rect 214012 114514 214064 114520
rect 214010 113656 214066 113665
rect 214010 113591 214066 113600
rect 213920 113280 213972 113286
rect 213918 113248 213920 113257
rect 213972 113248 213974 113257
rect 214024 113218 214052 113591
rect 213918 113183 213974 113192
rect 214012 113212 214064 113218
rect 214012 113154 214064 113160
rect 214010 112296 214066 112305
rect 214010 112231 214066 112240
rect 213920 111920 213972 111926
rect 213918 111888 213920 111897
rect 213972 111888 213974 111897
rect 214024 111858 214052 112231
rect 213918 111823 213974 111832
rect 214012 111852 214064 111858
rect 214012 111794 214064 111800
rect 214010 110936 214066 110945
rect 214010 110871 214066 110880
rect 214024 110566 214052 110871
rect 214012 110560 214064 110566
rect 213918 110528 213974 110537
rect 214012 110502 214064 110508
rect 213918 110463 213920 110472
rect 213972 110463 213974 110472
rect 213920 110434 213972 110440
rect 214010 109712 214066 109721
rect 214010 109647 214066 109656
rect 213918 109304 213974 109313
rect 213918 109239 213974 109248
rect 213932 109070 213960 109239
rect 214024 109138 214052 109647
rect 214012 109132 214064 109138
rect 214012 109074 214064 109080
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108352 214066 108361
rect 214010 108287 214066 108296
rect 213918 107944 213974 107953
rect 213918 107879 213974 107888
rect 213932 107710 213960 107879
rect 214024 107778 214052 108287
rect 214012 107772 214064 107778
rect 214012 107714 214064 107720
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 214010 106992 214066 107001
rect 214010 106927 214066 106936
rect 213918 106584 213974 106593
rect 213918 106519 213974 106528
rect 213932 106350 213960 106519
rect 214024 106418 214052 106927
rect 214012 106412 214064 106418
rect 214012 106354 214064 106360
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 213458 105768 213514 105777
rect 213458 105703 213514 105712
rect 213472 85474 213500 105703
rect 214010 105360 214066 105369
rect 214010 105295 214066 105304
rect 213918 105088 213974 105097
rect 214024 105058 214052 105295
rect 213918 105023 213974 105032
rect 214012 105052 214064 105058
rect 213932 104990 213960 105023
rect 214012 104994 214064 105000
rect 213920 104984 213972 104990
rect 213920 104926 213972 104932
rect 214010 104000 214066 104009
rect 214010 103935 214066 103944
rect 213918 103728 213974 103737
rect 213918 103663 213974 103672
rect 213932 103562 213960 103663
rect 214024 103630 214052 103935
rect 214012 103624 214064 103630
rect 214012 103566 214064 103572
rect 213920 103556 213972 103562
rect 213920 103498 213972 103504
rect 213918 102640 213974 102649
rect 213918 102575 213974 102584
rect 213932 102202 213960 102575
rect 213920 102196 213972 102202
rect 213920 102138 213972 102144
rect 213918 100872 213974 100881
rect 213918 100807 213974 100816
rect 213932 100774 213960 100807
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214010 99784 214066 99793
rect 214010 99719 214066 99728
rect 213918 99512 213974 99521
rect 213918 99447 213920 99456
rect 213972 99447 213974 99456
rect 213920 99418 213972 99424
rect 214024 99414 214052 99719
rect 214012 99408 214064 99414
rect 214012 99350 214064 99356
rect 214010 98424 214066 98433
rect 214010 98359 214066 98368
rect 214024 98122 214052 98359
rect 214012 98116 214064 98122
rect 214012 98058 214064 98064
rect 213920 98048 213972 98054
rect 213918 98016 213920 98025
rect 213972 98016 213974 98025
rect 213918 97951 213974 97960
rect 213918 97064 213974 97073
rect 213918 96999 213974 97008
rect 213932 96694 213960 96999
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 213918 95840 213974 95849
rect 213918 95775 213974 95784
rect 213932 95266 213960 95775
rect 213920 95260 213972 95266
rect 213920 95202 213972 95208
rect 214576 94518 214604 136711
rect 214654 135552 214710 135561
rect 214654 135487 214710 135496
rect 214668 97306 214696 135487
rect 214746 127528 214802 127537
rect 214746 127463 214802 127472
rect 214656 97300 214708 97306
rect 214656 97242 214708 97248
rect 214564 94512 214616 94518
rect 214564 94454 214616 94460
rect 214760 93158 214788 127463
rect 214838 101144 214894 101153
rect 214838 101079 214894 101088
rect 214748 93152 214800 93158
rect 214748 93094 214800 93100
rect 214562 90400 214618 90409
rect 214562 90335 214618 90344
rect 213460 85468 213512 85474
rect 213460 85410 213512 85416
rect 213368 85400 213420 85406
rect 213368 85342 213420 85348
rect 213276 79960 213328 79966
rect 213276 79902 213328 79908
rect 207664 78668 207716 78674
rect 207664 78610 207716 78616
rect 206284 26988 206336 26994
rect 206284 26930 206336 26936
rect 203524 21548 203576 21554
rect 203524 21490 203576 21496
rect 202144 7744 202196 7750
rect 202144 7686 202196 7692
rect 198096 3528 198148 3534
rect 198096 3470 198148 3476
rect 214576 3466 214604 90335
rect 214852 84182 214880 101079
rect 214930 96656 214986 96665
rect 214930 96591 214986 96600
rect 214944 86970 214972 96591
rect 214932 86964 214984 86970
rect 214932 86906 214984 86912
rect 214840 84176 214892 84182
rect 214840 84118 214892 84124
rect 215956 64326 215984 397530
rect 291844 397520 291896 397526
rect 291844 397462 291896 397468
rect 260104 393372 260156 393378
rect 260104 393314 260156 393320
rect 249064 384328 249116 384334
rect 249064 384270 249116 384276
rect 244924 343664 244976 343670
rect 244924 343606 244976 343612
rect 220084 337476 220136 337482
rect 220084 337418 220136 337424
rect 216036 328500 216088 328506
rect 216036 328442 216088 328448
rect 215944 64320 215996 64326
rect 215944 64262 215996 64268
rect 216048 4078 216076 328442
rect 216128 319524 216180 319530
rect 216128 319466 216180 319472
rect 216036 4072 216088 4078
rect 216036 4014 216088 4020
rect 216140 3466 216168 319466
rect 218704 292732 218756 292738
rect 218704 292674 218756 292680
rect 217324 198144 217376 198150
rect 217324 198086 217376 198092
rect 217336 178974 217364 198086
rect 217324 178968 217376 178974
rect 217324 178910 217376 178916
rect 218716 178673 218744 292674
rect 220096 178702 220124 337418
rect 231124 314696 231176 314702
rect 231124 314638 231176 314644
rect 226984 313336 227036 313342
rect 226984 313278 227036 313284
rect 220176 301232 220228 301238
rect 220176 301174 220228 301180
rect 220188 180266 220216 301174
rect 222844 294092 222896 294098
rect 222844 294034 222896 294040
rect 221464 270564 221516 270570
rect 221464 270506 221516 270512
rect 220268 252680 220320 252686
rect 220268 252622 220320 252628
rect 220280 181830 220308 252622
rect 220268 181824 220320 181830
rect 220268 181766 220320 181772
rect 220176 180260 220228 180266
rect 220176 180202 220228 180208
rect 220084 178696 220136 178702
rect 218702 178664 218758 178673
rect 220084 178638 220136 178644
rect 218702 178599 218758 178608
rect 221476 176050 221504 270506
rect 221556 249824 221608 249830
rect 221556 249766 221608 249772
rect 221568 177857 221596 249766
rect 222856 195498 222884 294034
rect 225604 289944 225656 289950
rect 225604 289886 225656 289892
rect 224224 281580 224276 281586
rect 224224 281522 224276 281528
rect 222936 232688 222988 232694
rect 222936 232630 222988 232636
rect 222844 195492 222896 195498
rect 222844 195434 222896 195440
rect 221648 192636 221700 192642
rect 221648 192578 221700 192584
rect 221554 177848 221610 177857
rect 221554 177783 221610 177792
rect 221660 177614 221688 192578
rect 222948 180402 222976 232630
rect 223028 199572 223080 199578
rect 223028 199514 223080 199520
rect 223040 180470 223068 199514
rect 223028 180464 223080 180470
rect 223028 180406 223080 180412
rect 222936 180396 222988 180402
rect 222936 180338 222988 180344
rect 221648 177608 221700 177614
rect 221648 177550 221700 177556
rect 221464 176044 221516 176050
rect 221464 175986 221516 175992
rect 224236 175982 224264 281522
rect 224316 278044 224368 278050
rect 224316 277986 224368 277992
rect 224328 189689 224356 277986
rect 224314 189680 224370 189689
rect 224314 189615 224370 189624
rect 225616 180334 225644 289886
rect 225696 206372 225748 206378
rect 225696 206314 225748 206320
rect 225604 180328 225656 180334
rect 225604 180270 225656 180276
rect 224960 178900 225012 178906
rect 224960 178842 225012 178848
rect 224224 175976 224276 175982
rect 224224 175918 224276 175924
rect 224972 175846 225000 178842
rect 225708 176118 225736 206314
rect 226996 177449 227024 313278
rect 228456 303816 228508 303822
rect 228456 303758 228508 303764
rect 227076 299736 227128 299742
rect 227076 299678 227128 299684
rect 226982 177440 227038 177449
rect 226982 177375 227038 177384
rect 227088 176361 227116 299678
rect 228364 278792 228416 278798
rect 228364 278734 228416 278740
rect 227168 256760 227220 256766
rect 227168 256702 227220 256708
rect 227180 177546 227208 256702
rect 227168 177540 227220 177546
rect 227168 177482 227220 177488
rect 228376 176662 228404 278734
rect 228468 201142 228496 303758
rect 231136 235346 231164 314638
rect 240784 302320 240836 302326
rect 240784 302262 240836 302268
rect 234620 295452 234672 295458
rect 234620 295394 234672 295400
rect 233884 288448 233936 288454
rect 233884 288390 233936 288396
rect 231952 269204 232004 269210
rect 231952 269146 232004 269152
rect 231216 268388 231268 268394
rect 231216 268330 231268 268336
rect 231228 239426 231256 268330
rect 231216 239420 231268 239426
rect 231216 239362 231268 239368
rect 231124 235340 231176 235346
rect 231124 235282 231176 235288
rect 229284 231192 229336 231198
rect 229284 231134 229336 231140
rect 228456 201136 228508 201142
rect 228456 201078 228508 201084
rect 229192 189916 229244 189922
rect 229192 189858 229244 189864
rect 228364 176656 228416 176662
rect 228364 176598 228416 176604
rect 227074 176352 227130 176361
rect 227074 176287 227130 176296
rect 229098 176352 229154 176361
rect 229098 176287 229154 176296
rect 225696 176112 225748 176118
rect 225696 176054 225748 176060
rect 224960 175840 225012 175846
rect 227720 175840 227772 175846
rect 224960 175782 225012 175788
rect 227718 175808 227720 175817
rect 227772 175808 227774 175817
rect 227718 175743 227774 175752
rect 229112 174321 229140 176287
rect 229098 174312 229154 174321
rect 229098 174247 229154 174256
rect 229204 161537 229232 189858
rect 229190 161528 229246 161537
rect 229190 161463 229246 161472
rect 229296 146849 229324 231134
rect 230480 229900 230532 229906
rect 230480 229842 230532 229848
rect 229560 177608 229612 177614
rect 229560 177550 229612 177556
rect 229468 176656 229520 176662
rect 229468 176598 229520 176604
rect 229376 176044 229428 176050
rect 229376 175986 229428 175992
rect 229388 171873 229416 175986
rect 229480 172825 229508 176598
rect 229572 173777 229600 177550
rect 229558 173768 229614 173777
rect 229558 173703 229614 173712
rect 229466 172816 229522 172825
rect 229466 172751 229522 172760
rect 229374 171864 229430 171873
rect 229374 171799 229430 171808
rect 229928 163736 229980 163742
rect 229928 163678 229980 163684
rect 229744 163532 229796 163538
rect 229744 163474 229796 163480
rect 229282 146840 229338 146849
rect 229282 146775 229338 146784
rect 229756 142497 229784 163474
rect 229940 143449 229968 163678
rect 230492 158681 230520 229842
rect 230572 224256 230624 224262
rect 230572 224198 230624 224204
rect 230584 166326 230612 224198
rect 230664 194132 230716 194138
rect 230664 194074 230716 194080
rect 230572 166320 230624 166326
rect 230572 166262 230624 166268
rect 230478 158672 230534 158681
rect 230478 158607 230534 158616
rect 230110 157448 230166 157457
rect 230110 157383 230166 157392
rect 229926 143440 229982 143449
rect 229926 143375 229982 143384
rect 230020 142860 230072 142866
rect 230020 142802 230072 142808
rect 229742 142488 229798 142497
rect 229742 142423 229798 142432
rect 229928 139460 229980 139466
rect 229928 139402 229980 139408
rect 229836 136672 229888 136678
rect 229836 136614 229888 136620
rect 229744 113212 229796 113218
rect 229744 113154 229796 113160
rect 216220 102808 216272 102814
rect 216220 102750 216272 102756
rect 216232 92274 216260 102750
rect 226984 95940 227036 95946
rect 226984 95882 227036 95888
rect 222844 94580 222896 94586
rect 222844 94522 222896 94528
rect 216220 92268 216272 92274
rect 216220 92210 216272 92216
rect 222856 65618 222884 94522
rect 224224 94512 224276 94518
rect 224224 94454 224276 94460
rect 222844 65612 222896 65618
rect 222844 65554 222896 65560
rect 224236 22846 224264 94454
rect 226996 66910 227024 95882
rect 228364 95260 228416 95266
rect 228364 95202 228416 95208
rect 226984 66904 227036 66910
rect 226984 66846 227036 66852
rect 228376 60042 228404 95202
rect 228364 60036 228416 60042
rect 228364 59978 228416 59984
rect 224224 22840 224276 22846
rect 224224 22782 224276 22788
rect 229756 8974 229784 113154
rect 229848 46306 229876 136614
rect 229940 55894 229968 139402
rect 230032 98977 230060 142802
rect 230124 137873 230152 157383
rect 230480 152584 230532 152590
rect 230480 152526 230532 152532
rect 230492 150657 230520 152526
rect 230478 150648 230534 150657
rect 230478 150583 230534 150592
rect 230676 140729 230704 194074
rect 230756 182912 230808 182918
rect 230756 182854 230808 182860
rect 230768 147801 230796 182854
rect 231400 173868 231452 173874
rect 231400 173810 231452 173816
rect 231412 173369 231440 173810
rect 231398 173360 231454 173369
rect 231398 173295 231454 173304
rect 231676 172440 231728 172446
rect 231676 172382 231728 172388
rect 231766 172408 231822 172417
rect 231688 171465 231716 172382
rect 231766 172343 231768 172352
rect 231820 172343 231822 172352
rect 231768 172314 231820 172320
rect 231674 171456 231730 171465
rect 231674 171391 231730 171400
rect 231768 171080 231820 171086
rect 231768 171022 231820 171028
rect 231676 170944 231728 170950
rect 231674 170912 231676 170921
rect 231728 170912 231730 170921
rect 231674 170847 231730 170856
rect 231780 170513 231808 171022
rect 231766 170504 231822 170513
rect 231766 170439 231822 170448
rect 231768 170196 231820 170202
rect 231768 170138 231820 170144
rect 231780 169969 231808 170138
rect 231766 169960 231822 169969
rect 231766 169895 231822 169904
rect 231676 169720 231728 169726
rect 231676 169662 231728 169668
rect 231400 169652 231452 169658
rect 231400 169594 231452 169600
rect 231412 168609 231440 169594
rect 231688 169017 231716 169662
rect 231768 169584 231820 169590
rect 231766 169552 231768 169561
rect 231820 169552 231822 169561
rect 231766 169487 231822 169496
rect 231674 169008 231730 169017
rect 231674 168943 231730 168952
rect 231398 168600 231454 168609
rect 231398 168535 231454 168544
rect 231768 168360 231820 168366
rect 231768 168302 231820 168308
rect 231780 168065 231808 168302
rect 231766 168056 231822 168065
rect 231216 168020 231268 168026
rect 231766 167991 231822 168000
rect 231216 167962 231268 167968
rect 231228 167113 231256 167962
rect 231214 167104 231270 167113
rect 231214 167039 231270 167048
rect 231768 167000 231820 167006
rect 231768 166942 231820 166948
rect 231492 166932 231544 166938
rect 231492 166874 231544 166880
rect 230940 166320 230992 166326
rect 230940 166262 230992 166268
rect 230952 156233 230980 166262
rect 231504 166161 231532 166874
rect 231780 166705 231808 166942
rect 231766 166696 231822 166705
rect 231766 166631 231822 166640
rect 231584 166320 231636 166326
rect 231584 166262 231636 166268
rect 231490 166152 231546 166161
rect 231490 166087 231546 166096
rect 231596 165753 231624 166262
rect 231582 165744 231638 165753
rect 231582 165679 231638 165688
rect 231032 165572 231084 165578
rect 231032 165514 231084 165520
rect 231044 165209 231072 165514
rect 231124 165504 231176 165510
rect 231124 165446 231176 165452
rect 231030 165200 231086 165209
rect 231030 165135 231086 165144
rect 231136 164393 231164 165446
rect 231122 164384 231178 164393
rect 231122 164319 231178 164328
rect 231768 164212 231820 164218
rect 231768 164154 231820 164160
rect 231676 164144 231728 164150
rect 231676 164086 231728 164092
rect 231492 164076 231544 164082
rect 231492 164018 231544 164024
rect 231504 162897 231532 164018
rect 231688 163441 231716 164086
rect 231780 163849 231808 164154
rect 231766 163840 231822 163849
rect 231766 163775 231822 163784
rect 231674 163432 231730 163441
rect 231674 163367 231730 163376
rect 231490 162888 231546 162897
rect 231490 162823 231546 162832
rect 231768 162784 231820 162790
rect 231768 162726 231820 162732
rect 231780 161945 231808 162726
rect 231964 162489 231992 269146
rect 232136 269136 232188 269142
rect 232136 269078 232188 269084
rect 232044 176112 232096 176118
rect 232044 176054 232096 176060
rect 231950 162480 232006 162489
rect 231950 162415 232006 162424
rect 231766 161936 231822 161945
rect 231766 161871 231822 161880
rect 231768 161424 231820 161430
rect 231768 161366 231820 161372
rect 231308 161356 231360 161362
rect 231308 161298 231360 161304
rect 231320 160993 231348 161298
rect 231306 160984 231362 160993
rect 231306 160919 231362 160928
rect 231780 160585 231808 161366
rect 231766 160576 231822 160585
rect 231766 160511 231822 160520
rect 231768 160064 231820 160070
rect 231582 160032 231638 160041
rect 231032 159996 231084 160002
rect 231768 160006 231820 160012
rect 231582 159967 231638 159976
rect 231032 159938 231084 159944
rect 231044 159633 231072 159938
rect 231596 159934 231624 159967
rect 231584 159928 231636 159934
rect 231584 159870 231636 159876
rect 231030 159624 231086 159633
rect 231030 159559 231086 159568
rect 231780 159089 231808 160006
rect 231766 159080 231822 159089
rect 231766 159015 231822 159024
rect 231768 158704 231820 158710
rect 231768 158646 231820 158652
rect 231216 158636 231268 158642
rect 231216 158578 231268 158584
rect 231228 158137 231256 158578
rect 231214 158128 231270 158137
rect 231214 158063 231270 158072
rect 231780 157729 231808 158646
rect 231766 157720 231822 157729
rect 231766 157655 231822 157664
rect 231768 157344 231820 157350
rect 231768 157286 231820 157292
rect 231124 157276 231176 157282
rect 231124 157218 231176 157224
rect 231136 156777 231164 157218
rect 231780 157185 231808 157286
rect 231766 157176 231822 157185
rect 231766 157111 231822 157120
rect 231584 156800 231636 156806
rect 231122 156768 231178 156777
rect 231584 156742 231636 156748
rect 231122 156703 231178 156712
rect 230938 156224 230994 156233
rect 230938 156159 230994 156168
rect 231492 155916 231544 155922
rect 231492 155858 231544 155864
rect 231504 154873 231532 155858
rect 231490 154864 231546 154873
rect 231490 154799 231546 154808
rect 231124 153808 231176 153814
rect 231124 153750 231176 153756
rect 230754 147792 230810 147801
rect 230754 147727 230810 147736
rect 230848 146056 230900 146062
rect 230848 145998 230900 146004
rect 230860 145897 230888 145998
rect 230846 145888 230902 145897
rect 230846 145823 230902 145832
rect 230662 140720 230718 140729
rect 230662 140655 230718 140664
rect 230110 137864 230166 137873
rect 230110 137799 230166 137808
rect 230756 136536 230808 136542
rect 230756 136478 230808 136484
rect 230768 135425 230796 136478
rect 230754 135416 230810 135425
rect 230754 135351 230810 135360
rect 230572 135108 230624 135114
rect 230572 135050 230624 135056
rect 230584 134065 230612 135050
rect 230570 134056 230626 134065
rect 230570 133991 230626 134000
rect 230664 132388 230716 132394
rect 230664 132330 230716 132336
rect 230676 132161 230704 132330
rect 230662 132152 230718 132161
rect 230662 132087 230718 132096
rect 231136 126041 231164 153750
rect 231596 152017 231624 156742
rect 231768 155848 231820 155854
rect 232056 155825 232084 176054
rect 231768 155790 231820 155796
rect 232042 155816 232098 155825
rect 231780 155281 231808 155790
rect 232042 155751 232098 155760
rect 231766 155272 231822 155281
rect 231766 155207 231822 155216
rect 231768 154556 231820 154562
rect 231768 154498 231820 154504
rect 231676 154488 231728 154494
rect 231676 154430 231728 154436
rect 231688 153921 231716 154430
rect 231780 154329 231808 154498
rect 231766 154320 231822 154329
rect 231766 154255 231822 154264
rect 231674 153912 231730 153921
rect 231674 153847 231730 153856
rect 231768 153196 231820 153202
rect 231768 153138 231820 153144
rect 231780 152969 231808 153138
rect 231766 152960 231822 152969
rect 231766 152895 231822 152904
rect 231582 152008 231638 152017
rect 231582 151943 231638 151952
rect 232148 151814 232176 269078
rect 233240 238264 233292 238270
rect 233240 238206 233292 238212
rect 232688 156732 232740 156738
rect 232688 156674 232740 156680
rect 231872 151786 232176 151814
rect 231676 151768 231728 151774
rect 231676 151710 231728 151716
rect 231688 151065 231716 151710
rect 231768 151700 231820 151706
rect 231768 151642 231820 151648
rect 231780 151609 231808 151642
rect 231766 151600 231822 151609
rect 231766 151535 231822 151544
rect 231674 151056 231730 151065
rect 231674 150991 231730 151000
rect 231676 150408 231728 150414
rect 231676 150350 231728 150356
rect 231688 149161 231716 150350
rect 231768 149864 231820 149870
rect 231768 149806 231820 149812
rect 231780 149705 231808 149806
rect 231766 149696 231822 149705
rect 231766 149631 231822 149640
rect 231674 149152 231730 149161
rect 231674 149087 231730 149096
rect 231308 148980 231360 148986
rect 231308 148922 231360 148928
rect 231320 148209 231348 148922
rect 231306 148200 231362 148209
rect 231306 148135 231362 148144
rect 231216 147756 231268 147762
rect 231216 147698 231268 147704
rect 231228 127401 231256 147698
rect 231766 146296 231822 146305
rect 231766 146231 231822 146240
rect 231780 146198 231808 146231
rect 231768 146192 231820 146198
rect 231768 146134 231820 146140
rect 231400 146124 231452 146130
rect 231400 146066 231452 146072
rect 231412 145353 231440 146066
rect 231398 145344 231454 145353
rect 231398 145279 231454 145288
rect 231766 144392 231822 144401
rect 231872 144378 231900 151786
rect 232700 146062 232728 156674
rect 233252 152590 233280 238206
rect 233896 220182 233924 288390
rect 233884 220176 233936 220182
rect 233884 220118 233936 220124
rect 233424 218816 233476 218822
rect 233424 218758 233476 218764
rect 233332 196852 233384 196858
rect 233332 196794 233384 196800
rect 233240 152584 233292 152590
rect 233240 152526 233292 152532
rect 232688 146056 232740 146062
rect 232688 145998 232740 146004
rect 232596 145580 232648 145586
rect 232596 145522 232648 145528
rect 232504 145104 232556 145110
rect 232504 145046 232556 145052
rect 231822 144350 231900 144378
rect 231766 144327 231822 144336
rect 231768 144016 231820 144022
rect 231766 143984 231768 143993
rect 231820 143984 231822 143993
rect 231766 143919 231822 143928
rect 231768 143540 231820 143546
rect 231768 143482 231820 143488
rect 231780 143041 231808 143482
rect 231766 143032 231822 143041
rect 231766 142967 231822 142976
rect 231492 142112 231544 142118
rect 231492 142054 231544 142060
rect 231504 141137 231532 142054
rect 231768 142044 231820 142050
rect 231768 141986 231820 141992
rect 231780 141681 231808 141986
rect 231766 141672 231822 141681
rect 231766 141607 231822 141616
rect 231490 141128 231546 141137
rect 231490 141063 231546 141072
rect 231400 140072 231452 140078
rect 231400 140014 231452 140020
rect 231308 139800 231360 139806
rect 231306 139768 231308 139777
rect 231360 139768 231362 139777
rect 231306 139703 231362 139712
rect 231308 139324 231360 139330
rect 231308 139266 231360 139272
rect 231320 139233 231348 139266
rect 231306 139224 231362 139233
rect 231306 139159 231362 139168
rect 231412 138122 231440 140014
rect 231768 139256 231820 139262
rect 231768 139198 231820 139204
rect 231780 138825 231808 139198
rect 231766 138816 231822 138825
rect 231766 138751 231822 138760
rect 231584 138712 231636 138718
rect 231584 138654 231636 138660
rect 231492 138304 231544 138310
rect 231490 138272 231492 138281
rect 231544 138272 231546 138281
rect 231490 138207 231546 138216
rect 231320 138094 231440 138122
rect 231320 129849 231348 138094
rect 231400 137964 231452 137970
rect 231400 137906 231452 137912
rect 231412 137329 231440 137906
rect 231398 137320 231454 137329
rect 231398 137255 231454 137264
rect 231400 136604 231452 136610
rect 231400 136546 231452 136552
rect 231412 135969 231440 136546
rect 231398 135960 231454 135969
rect 231398 135895 231454 135904
rect 231596 132569 231624 138654
rect 231768 137896 231820 137902
rect 231768 137838 231820 137844
rect 231780 136921 231808 137838
rect 231766 136912 231822 136921
rect 231766 136847 231822 136856
rect 231768 135244 231820 135250
rect 231768 135186 231820 135192
rect 231676 135176 231728 135182
rect 231676 135118 231728 135124
rect 231688 134473 231716 135118
rect 231780 135017 231808 135186
rect 231766 135008 231822 135017
rect 231766 134943 231822 134952
rect 231674 134464 231730 134473
rect 231674 134399 231730 134408
rect 231768 133884 231820 133890
rect 231768 133826 231820 133832
rect 231676 133816 231728 133822
rect 231676 133758 231728 133764
rect 231688 133113 231716 133758
rect 231780 133521 231808 133826
rect 231766 133512 231822 133521
rect 231766 133447 231822 133456
rect 231674 133104 231730 133113
rect 231674 133039 231730 133048
rect 231582 132560 231638 132569
rect 231582 132495 231638 132504
rect 231676 132456 231728 132462
rect 231676 132398 231728 132404
rect 231688 131617 231716 132398
rect 231768 132320 231820 132326
rect 231768 132262 231820 132268
rect 231674 131608 231730 131617
rect 231674 131543 231730 131552
rect 231780 131209 231808 132262
rect 231766 131200 231822 131209
rect 231766 131135 231822 131144
rect 231768 131096 231820 131102
rect 231768 131038 231820 131044
rect 231400 131028 231452 131034
rect 231400 130970 231452 130976
rect 231412 130257 231440 130970
rect 231780 130665 231808 131038
rect 231766 130656 231822 130665
rect 231766 130591 231822 130600
rect 231584 130416 231636 130422
rect 231584 130358 231636 130364
rect 231398 130248 231454 130257
rect 231398 130183 231454 130192
rect 231306 129840 231362 129849
rect 231306 129775 231362 129784
rect 231400 129668 231452 129674
rect 231400 129610 231452 129616
rect 231412 128897 231440 129610
rect 231398 128888 231454 128897
rect 231398 128823 231454 128832
rect 231492 127628 231544 127634
rect 231492 127570 231544 127576
rect 231214 127392 231270 127401
rect 231214 127327 231270 127336
rect 231122 126032 231178 126041
rect 231122 125967 231178 125976
rect 231308 125588 231360 125594
rect 231308 125530 231360 125536
rect 231320 125089 231348 125530
rect 231306 125080 231362 125089
rect 231306 125015 231362 125024
rect 231504 124386 231532 127570
rect 231596 125497 231624 130358
rect 231768 129736 231820 129742
rect 231768 129678 231820 129684
rect 231780 129305 231808 129678
rect 231766 129296 231822 129305
rect 231766 129231 231822 129240
rect 231766 128344 231822 128353
rect 231676 128308 231728 128314
rect 231766 128279 231822 128288
rect 231676 128250 231728 128256
rect 231688 127945 231716 128250
rect 231780 128246 231808 128279
rect 231768 128240 231820 128246
rect 231768 128182 231820 128188
rect 231674 127936 231730 127945
rect 231674 127871 231730 127880
rect 231766 126984 231822 126993
rect 231676 126948 231728 126954
rect 231766 126919 231822 126928
rect 231676 126890 231728 126896
rect 231688 126449 231716 126890
rect 231780 126886 231808 126919
rect 231768 126880 231820 126886
rect 231768 126822 231820 126828
rect 231674 126440 231730 126449
rect 231674 126375 231730 126384
rect 231676 125520 231728 125526
rect 231582 125488 231638 125497
rect 231676 125462 231728 125468
rect 231582 125423 231638 125432
rect 231688 124545 231716 125462
rect 231766 124808 231822 124817
rect 231766 124743 231822 124752
rect 231674 124536 231730 124545
rect 231674 124471 231730 124480
rect 231504 124358 231716 124386
rect 231492 124160 231544 124166
rect 231492 124102 231544 124108
rect 231308 124092 231360 124098
rect 231308 124034 231360 124040
rect 231320 123593 231348 124034
rect 231306 123584 231362 123593
rect 231306 123519 231362 123528
rect 231308 123480 231360 123486
rect 231308 123422 231360 123428
rect 231124 120964 231176 120970
rect 231124 120906 231176 120912
rect 231136 120737 231164 120906
rect 231122 120728 231178 120737
rect 231122 120663 231178 120672
rect 231320 119785 231348 123422
rect 231504 123185 231532 124102
rect 231490 123176 231546 123185
rect 231490 123111 231546 123120
rect 231492 122732 231544 122738
rect 231492 122674 231544 122680
rect 231504 121689 231532 122674
rect 231584 122664 231636 122670
rect 231582 122632 231584 122641
rect 231636 122632 231638 122641
rect 231582 122567 231638 122576
rect 231490 121680 231546 121689
rect 231490 121615 231546 121624
rect 231492 121372 231544 121378
rect 231492 121314 231544 121320
rect 231504 120329 231532 121314
rect 231490 120320 231546 120329
rect 231490 120255 231546 120264
rect 231400 120012 231452 120018
rect 231400 119954 231452 119960
rect 231306 119776 231362 119785
rect 231306 119711 231362 119720
rect 231308 119400 231360 119406
rect 231412 119377 231440 119954
rect 231308 119342 231360 119348
rect 231398 119368 231454 119377
rect 231124 118516 231176 118522
rect 231124 118458 231176 118464
rect 231136 118017 231164 118458
rect 231122 118008 231178 118017
rect 231122 117943 231178 117952
rect 231216 116816 231268 116822
rect 231216 116758 231268 116764
rect 231124 116612 231176 116618
rect 231124 116554 231176 116560
rect 230664 115796 230716 115802
rect 230664 115738 230716 115744
rect 230676 115569 230704 115738
rect 230662 115560 230718 115569
rect 230662 115495 230718 115504
rect 230572 114844 230624 114850
rect 230572 114786 230624 114792
rect 230584 114617 230612 114786
rect 230570 114608 230626 114617
rect 230570 114543 230626 114552
rect 230572 114436 230624 114442
rect 230572 114378 230624 114384
rect 230584 113257 230612 114378
rect 231136 114209 231164 116554
rect 231122 114200 231178 114209
rect 231122 114135 231178 114144
rect 230664 113824 230716 113830
rect 230664 113766 230716 113772
rect 230570 113248 230626 113257
rect 230570 113183 230626 113192
rect 230572 112532 230624 112538
rect 230572 112474 230624 112480
rect 230584 107953 230612 112474
rect 230676 109449 230704 113766
rect 231124 112464 231176 112470
rect 231124 112406 231176 112412
rect 230662 109440 230718 109449
rect 230662 109375 230718 109384
rect 230570 107944 230626 107953
rect 230570 107879 230626 107888
rect 231136 103329 231164 112406
rect 231228 112305 231256 116758
rect 231214 112296 231270 112305
rect 231214 112231 231270 112240
rect 231122 103320 231178 103329
rect 231122 103255 231178 103264
rect 230572 103012 230624 103018
rect 230572 102954 230624 102960
rect 230584 102785 230612 102954
rect 230570 102776 230626 102785
rect 230570 102711 230626 102720
rect 231124 102196 231176 102202
rect 231124 102138 231176 102144
rect 230940 99612 230992 99618
rect 230940 99554 230992 99560
rect 230018 98968 230074 98977
rect 230018 98903 230074 98912
rect 230480 98252 230532 98258
rect 230480 98194 230532 98200
rect 230492 98025 230520 98194
rect 230478 98016 230534 98025
rect 230478 97951 230534 97960
rect 230952 97617 230980 99554
rect 230938 97608 230994 97617
rect 230938 97543 230994 97552
rect 230478 97064 230534 97073
rect 230478 96999 230534 97008
rect 230492 96694 230520 96999
rect 230480 96688 230532 96694
rect 230480 96630 230532 96636
rect 229928 55888 229980 55894
rect 229928 55830 229980 55836
rect 229836 46300 229888 46306
rect 229836 46242 229888 46248
rect 230492 11014 230520 96630
rect 230570 95704 230626 95713
rect 230570 95639 230626 95648
rect 230584 88330 230612 95639
rect 230572 88324 230624 88330
rect 230572 88266 230624 88272
rect 231136 28286 231164 102138
rect 231320 98569 231348 119342
rect 231398 119303 231454 119312
rect 231492 118652 231544 118658
rect 231492 118594 231544 118600
rect 231504 117473 231532 118594
rect 231490 117464 231546 117473
rect 231490 117399 231546 117408
rect 231492 117292 231544 117298
rect 231492 117234 231544 117240
rect 231504 116521 231532 117234
rect 231490 116512 231546 116521
rect 231490 116447 231546 116456
rect 231688 116113 231716 124358
rect 231780 124137 231808 124743
rect 231766 124128 231822 124137
rect 231766 124063 231822 124072
rect 231768 122800 231820 122806
rect 231768 122742 231820 122748
rect 231780 122233 231808 122742
rect 231766 122224 231822 122233
rect 231766 122159 231822 122168
rect 231768 121440 231820 121446
rect 231768 121382 231820 121388
rect 231780 121281 231808 121382
rect 231766 121272 231822 121281
rect 231766 121207 231822 121216
rect 231768 120080 231820 120086
rect 231768 120022 231820 120028
rect 231780 118969 231808 120022
rect 231766 118960 231822 118969
rect 231766 118895 231822 118904
rect 231768 118584 231820 118590
rect 231768 118526 231820 118532
rect 231780 118425 231808 118526
rect 231766 118416 231822 118425
rect 231766 118351 231822 118360
rect 231674 116104 231730 116113
rect 231674 116039 231730 116048
rect 231676 115524 231728 115530
rect 231676 115466 231728 115472
rect 231688 115161 231716 115466
rect 231674 115152 231730 115161
rect 231674 115087 231730 115096
rect 231768 114504 231820 114510
rect 231768 114446 231820 114452
rect 231780 113665 231808 114446
rect 231766 113656 231822 113665
rect 231766 113591 231822 113600
rect 231768 112872 231820 112878
rect 231768 112814 231820 112820
rect 231780 112713 231808 112814
rect 231766 112704 231822 112713
rect 231766 112639 231822 112648
rect 231768 111784 231820 111790
rect 231768 111726 231820 111732
rect 231492 111716 231544 111722
rect 231492 111658 231544 111664
rect 231504 110809 231532 111658
rect 231780 111353 231808 111726
rect 231766 111344 231822 111353
rect 231766 111279 231822 111288
rect 231490 110800 231546 110809
rect 231490 110735 231546 110744
rect 231768 110424 231820 110430
rect 231766 110392 231768 110401
rect 231820 110392 231822 110401
rect 231766 110327 231822 110336
rect 231768 110016 231820 110022
rect 231768 109958 231820 109964
rect 231780 109857 231808 109958
rect 231766 109848 231822 109857
rect 231766 109783 231822 109792
rect 231768 108996 231820 109002
rect 231768 108938 231820 108944
rect 231676 108928 231728 108934
rect 231780 108905 231808 108938
rect 231676 108870 231728 108876
rect 231766 108896 231822 108905
rect 231688 108497 231716 108870
rect 231766 108831 231822 108840
rect 231674 108488 231730 108497
rect 231674 108423 231730 108432
rect 231400 108316 231452 108322
rect 231400 108258 231452 108264
rect 231412 99929 231440 108258
rect 231768 107636 231820 107642
rect 231768 107578 231820 107584
rect 231676 107568 231728 107574
rect 231780 107545 231808 107578
rect 231676 107510 231728 107516
rect 231766 107536 231822 107545
rect 231688 107137 231716 107510
rect 231766 107471 231822 107480
rect 231674 107128 231730 107137
rect 231674 107063 231730 107072
rect 231768 107092 231820 107098
rect 231768 107034 231820 107040
rect 231780 106593 231808 107034
rect 231766 106584 231822 106593
rect 231766 106519 231822 106528
rect 231768 106276 231820 106282
rect 231768 106218 231820 106224
rect 231780 106185 231808 106218
rect 231766 106176 231822 106185
rect 231766 106111 231822 106120
rect 231676 105392 231728 105398
rect 231676 105334 231728 105340
rect 231688 105233 231716 105334
rect 231674 105224 231730 105233
rect 231674 105159 231730 105168
rect 231768 104848 231820 104854
rect 231768 104790 231820 104796
rect 231492 104780 231544 104786
rect 231492 104722 231544 104728
rect 231504 103737 231532 104722
rect 231676 104712 231728 104718
rect 231674 104680 231676 104689
rect 231728 104680 231730 104689
rect 231674 104615 231730 104624
rect 231780 104281 231808 104790
rect 231766 104272 231822 104281
rect 231766 104207 231822 104216
rect 231490 103728 231546 103737
rect 231490 103663 231546 103672
rect 232516 103018 232544 145046
rect 232608 114850 232636 145522
rect 232688 140888 232740 140894
rect 232688 140830 232740 140836
rect 232596 114844 232648 114850
rect 232596 114786 232648 114792
rect 232504 103012 232556 103018
rect 232504 102954 232556 102960
rect 232596 102264 232648 102270
rect 232596 102206 232648 102212
rect 231492 102128 231544 102134
rect 231492 102070 231544 102076
rect 231504 101833 231532 102070
rect 231768 101992 231820 101998
rect 231768 101934 231820 101940
rect 231490 101824 231546 101833
rect 231490 101759 231546 101768
rect 231584 101516 231636 101522
rect 231584 101458 231636 101464
rect 231596 101425 231624 101458
rect 231676 101448 231728 101454
rect 231582 101416 231638 101425
rect 231676 101390 231728 101396
rect 231582 101351 231638 101360
rect 231688 100473 231716 101390
rect 231780 100881 231808 101934
rect 231766 100872 231822 100881
rect 231766 100807 231822 100816
rect 231768 100700 231820 100706
rect 231768 100642 231820 100648
rect 231674 100464 231730 100473
rect 231674 100399 231730 100408
rect 231398 99920 231454 99929
rect 231398 99855 231454 99864
rect 231780 99521 231808 100642
rect 231766 99512 231822 99521
rect 231766 99447 231822 99456
rect 231306 98560 231362 98569
rect 231306 98495 231362 98504
rect 232504 98116 232556 98122
rect 232504 98058 232556 98064
rect 231216 98048 231268 98054
rect 231216 97990 231268 97996
rect 231228 37942 231256 97990
rect 231768 96756 231820 96762
rect 231768 96698 231820 96704
rect 231780 96665 231808 96698
rect 231766 96656 231822 96665
rect 231766 96591 231822 96600
rect 231216 37936 231268 37942
rect 231216 37878 231268 37884
rect 231124 28280 231176 28286
rect 231124 28222 231176 28228
rect 232516 11830 232544 98058
rect 232608 38010 232636 102206
rect 232700 98258 232728 140830
rect 232780 140820 232832 140826
rect 232780 140762 232832 140768
rect 232792 99618 232820 140762
rect 233344 139330 233372 196794
rect 233436 165510 233464 218758
rect 233424 165504 233476 165510
rect 233424 165446 233476 165452
rect 234160 162920 234212 162926
rect 234160 162862 234212 162868
rect 234068 161832 234120 161838
rect 234068 161774 234120 161780
rect 234080 159934 234108 161774
rect 234068 159928 234120 159934
rect 234068 159870 234120 159876
rect 234172 156618 234200 162862
rect 234080 156590 234200 156618
rect 233976 142928 234028 142934
rect 233976 142870 234028 142876
rect 233332 139324 233384 139330
rect 233332 139266 233384 139272
rect 233884 121508 233936 121514
rect 233884 121450 233936 121456
rect 233608 102332 233660 102338
rect 233608 102274 233660 102280
rect 232780 99612 232832 99618
rect 232780 99554 232832 99560
rect 232688 98252 232740 98258
rect 232688 98194 232740 98200
rect 233620 94586 233648 102274
rect 233608 94580 233660 94586
rect 233608 94522 233660 94528
rect 232596 38004 232648 38010
rect 232596 37946 232648 37952
rect 233896 20058 233924 121450
rect 233988 102134 234016 142870
rect 234080 122670 234108 156590
rect 234160 152516 234212 152522
rect 234160 152458 234212 152464
rect 234068 122664 234120 122670
rect 234068 122606 234120 122612
rect 234172 114442 234200 152458
rect 234632 148986 234660 295394
rect 234712 274712 234764 274718
rect 234712 274654 234764 274660
rect 234724 156806 234752 274654
rect 239036 263628 239088 263634
rect 239036 263570 239088 263576
rect 238852 250504 238904 250510
rect 238852 250446 238904 250452
rect 234804 245744 234856 245750
rect 234804 245686 234856 245692
rect 234712 156800 234764 156806
rect 234712 156742 234764 156748
rect 234620 148980 234672 148986
rect 234620 148922 234672 148928
rect 234816 144022 234844 245686
rect 236000 227044 236052 227050
rect 236000 226986 236052 226992
rect 234896 177540 234948 177546
rect 234896 177482 234948 177488
rect 234908 163742 234936 177482
rect 234896 163736 234948 163742
rect 234896 163678 234948 163684
rect 235448 150476 235500 150482
rect 235448 150418 235500 150424
rect 235264 149728 235316 149734
rect 235264 149670 235316 149676
rect 234804 144016 234856 144022
rect 234804 143958 234856 143964
rect 234252 137284 234304 137290
rect 234252 137226 234304 137232
rect 234160 114436 234212 114442
rect 234160 114378 234212 114384
rect 234068 109064 234120 109070
rect 234068 109006 234120 109012
rect 233976 102128 234028 102134
rect 233976 102070 234028 102076
rect 233976 96688 234028 96694
rect 233976 96630 234028 96636
rect 233988 93702 234016 96630
rect 233976 93696 234028 93702
rect 233976 93638 234028 93644
rect 233976 88324 234028 88330
rect 233976 88266 234028 88272
rect 233884 20052 233936 20058
rect 233884 19994 233936 20000
rect 232504 11824 232556 11830
rect 232504 11766 232556 11772
rect 230480 11008 230532 11014
rect 230480 10950 230532 10956
rect 229744 8968 229796 8974
rect 229744 8910 229796 8916
rect 214564 3460 214616 3466
rect 214564 3402 214616 3408
rect 216128 3460 216180 3466
rect 216128 3402 216180 3408
rect 233988 3058 234016 88266
rect 234080 49094 234108 109006
rect 234264 104718 234292 137226
rect 235276 111722 235304 149670
rect 235356 143608 235408 143614
rect 235356 143550 235408 143556
rect 235264 111716 235316 111722
rect 235264 111658 235316 111664
rect 235264 109132 235316 109138
rect 235264 109074 235316 109080
rect 234252 104712 234304 104718
rect 234252 104654 234304 104660
rect 234068 49088 234120 49094
rect 234068 49030 234120 49036
rect 235276 40798 235304 109074
rect 235368 101522 235396 143550
rect 235460 110022 235488 150418
rect 236012 149870 236040 226986
rect 237380 200932 237432 200938
rect 237380 200874 237432 200880
rect 236184 180464 236236 180470
rect 236184 180406 236236 180412
rect 236092 180396 236144 180402
rect 236092 180338 236144 180344
rect 236000 149864 236052 149870
rect 236000 149806 236052 149812
rect 235540 146328 235592 146334
rect 235540 146270 235592 146276
rect 235448 110016 235500 110022
rect 235448 109958 235500 109964
rect 235552 105398 235580 146270
rect 236104 138310 236132 180338
rect 236196 139806 236224 180406
rect 237392 170202 237420 200874
rect 238760 183048 238812 183054
rect 238760 182990 238812 182996
rect 237472 181824 237524 181830
rect 237472 181766 237524 181772
rect 237380 170196 237432 170202
rect 237380 170138 237432 170144
rect 237484 168026 237512 181766
rect 237564 181552 237616 181558
rect 237564 181494 237616 181500
rect 237576 170950 237604 181494
rect 237656 177472 237708 177478
rect 237656 177414 237708 177420
rect 237564 170944 237616 170950
rect 237564 170886 237616 170892
rect 237472 168020 237524 168026
rect 237472 167962 237524 167968
rect 237668 166326 237696 177414
rect 238772 173874 238800 182990
rect 238760 173868 238812 173874
rect 238760 173810 238812 173816
rect 238864 168366 238892 250446
rect 238944 178968 238996 178974
rect 238944 178910 238996 178916
rect 238852 168360 238904 168366
rect 238758 168328 238814 168337
rect 238852 168302 238904 168308
rect 238758 168263 238814 168272
rect 238024 167068 238076 167074
rect 238024 167010 238076 167016
rect 237656 166320 237708 166326
rect 237656 166262 237708 166268
rect 237380 157412 237432 157418
rect 237380 157354 237432 157360
rect 237392 154601 237420 157354
rect 237378 154592 237434 154601
rect 237378 154527 237434 154536
rect 236736 153264 236788 153270
rect 236736 153206 236788 153212
rect 236184 139800 236236 139806
rect 236184 139742 236236 139748
rect 236092 138304 236144 138310
rect 236092 138246 236144 138252
rect 236644 135312 236696 135318
rect 236644 135254 236696 135260
rect 235540 105392 235592 105398
rect 235540 105334 235592 105340
rect 235356 101516 235408 101522
rect 235356 101458 235408 101464
rect 235356 96688 235408 96694
rect 235356 96630 235408 96636
rect 235368 54534 235396 96630
rect 235356 54528 235408 54534
rect 235356 54470 235408 54476
rect 235264 40792 235316 40798
rect 235264 40734 235316 40740
rect 236656 31210 236684 135254
rect 236748 112878 236776 153206
rect 238036 147762 238064 167010
rect 238392 165640 238444 165646
rect 238392 165582 238444 165588
rect 238116 161492 238168 161498
rect 238116 161434 238168 161440
rect 238024 147756 238076 147762
rect 238024 147698 238076 147704
rect 236920 147688 236972 147694
rect 236920 147630 236972 147636
rect 236828 133952 236880 133958
rect 236828 133894 236880 133900
rect 236736 112872 236788 112878
rect 236736 112814 236788 112820
rect 236736 99408 236788 99414
rect 236736 99350 236788 99356
rect 236644 31204 236696 31210
rect 236644 31146 236696 31152
rect 236748 7614 236776 99350
rect 236840 66978 236868 133894
rect 236932 107098 236960 147630
rect 238024 138032 238076 138038
rect 238024 137974 238076 137980
rect 236920 107092 236972 107098
rect 236920 107034 236972 107040
rect 236828 66972 236880 66978
rect 236828 66914 236880 66920
rect 238036 46374 238064 137974
rect 238128 120970 238156 161434
rect 238208 155236 238260 155242
rect 238208 155178 238260 155184
rect 238116 120964 238168 120970
rect 238116 120906 238168 120912
rect 238220 115530 238248 155178
rect 238404 153814 238432 165582
rect 238772 161474 238800 168263
rect 238956 166938 238984 178910
rect 238944 166932 238996 166938
rect 238944 166874 238996 166880
rect 239048 164082 239076 263570
rect 240140 247104 240192 247110
rect 240140 247046 240192 247052
rect 240152 172666 240180 247046
rect 240232 196784 240284 196790
rect 240232 196726 240284 196732
rect 240060 172638 240180 172666
rect 239404 172576 239456 172582
rect 239404 172518 239456 172524
rect 239036 164076 239088 164082
rect 239036 164018 239088 164024
rect 238772 161446 238892 161474
rect 238864 161362 238892 161446
rect 238852 161356 238904 161362
rect 238852 161298 238904 161304
rect 238392 153808 238444 153814
rect 238392 153750 238444 153756
rect 238300 153332 238352 153338
rect 238300 153274 238352 153280
rect 238312 116822 238340 153274
rect 239416 135114 239444 172518
rect 240060 172446 240088 172638
rect 240140 172508 240192 172514
rect 240140 172450 240192 172456
rect 240048 172440 240100 172446
rect 240048 172382 240100 172388
rect 240152 169658 240180 172450
rect 240140 169652 240192 169658
rect 240140 169594 240192 169600
rect 240244 169590 240272 196726
rect 240324 181756 240376 181762
rect 240324 181698 240376 181704
rect 240336 172378 240364 181698
rect 240796 176730 240824 302262
rect 242900 245676 242952 245682
rect 242900 245618 242952 245624
rect 241796 240168 241848 240174
rect 241796 240110 241848 240116
rect 241612 201068 241664 201074
rect 241612 201010 241664 201016
rect 240784 176724 240836 176730
rect 240784 176666 240836 176672
rect 241520 176724 241572 176730
rect 241520 176666 241572 176672
rect 240416 175976 240468 175982
rect 240416 175918 240468 175924
rect 240324 172372 240376 172378
rect 240324 172314 240376 172320
rect 240232 169584 240284 169590
rect 240232 169526 240284 169532
rect 240140 163192 240192 163198
rect 240140 163134 240192 163140
rect 239496 160132 239548 160138
rect 239496 160074 239548 160080
rect 239404 135108 239456 135114
rect 239404 135050 239456 135056
rect 239404 120148 239456 120154
rect 239404 120090 239456 120096
rect 238300 116816 238352 116822
rect 238300 116758 238352 116764
rect 238208 115524 238260 115530
rect 238208 115466 238260 115472
rect 238300 114572 238352 114578
rect 238300 114514 238352 114520
rect 238208 110628 238260 110634
rect 238208 110570 238260 110576
rect 238116 99476 238168 99482
rect 238116 99418 238168 99424
rect 238024 46368 238076 46374
rect 238024 46310 238076 46316
rect 238128 15910 238156 99418
rect 238220 29714 238248 110570
rect 238312 35222 238340 114514
rect 238300 35216 238352 35222
rect 238300 35158 238352 35164
rect 238208 29708 238260 29714
rect 238208 29650 238260 29656
rect 238116 15904 238168 15910
rect 238116 15846 238168 15852
rect 239416 13190 239444 120090
rect 239508 120018 239536 160074
rect 240152 160002 240180 163134
rect 240428 161838 240456 175918
rect 241532 172514 241560 176666
rect 241520 172508 241572 172514
rect 241520 172450 241572 172456
rect 241624 169726 241652 201010
rect 241704 182980 241756 182986
rect 241704 182922 241756 182928
rect 241612 169720 241664 169726
rect 241612 169662 241664 169668
rect 240968 168496 241020 168502
rect 240968 168438 241020 168444
rect 240876 168428 240928 168434
rect 240876 168370 240928 168376
rect 240416 161832 240468 161838
rect 240416 161774 240468 161780
rect 240784 160200 240836 160206
rect 240784 160142 240836 160148
rect 240140 159996 240192 160002
rect 240140 159938 240192 159944
rect 239680 158772 239732 158778
rect 239680 158714 239732 158720
rect 239588 149116 239640 149122
rect 239588 149058 239640 149064
rect 239496 120012 239548 120018
rect 239496 119954 239548 119960
rect 239496 117360 239548 117366
rect 239496 117302 239548 117308
rect 239508 32434 239536 117302
rect 239600 108934 239628 149058
rect 239692 118522 239720 158714
rect 240796 121378 240824 160142
rect 240888 158642 240916 168370
rect 240876 158636 240928 158642
rect 240876 158578 240928 158584
rect 240876 155984 240928 155990
rect 240876 155926 240928 155932
rect 240784 121372 240836 121378
rect 240784 121314 240836 121320
rect 239680 118516 239732 118522
rect 239680 118458 239732 118464
rect 240888 115802 240916 155926
rect 240980 140078 241008 168438
rect 241716 161430 241744 182922
rect 241808 167006 241836 240110
rect 242256 171148 242308 171154
rect 242256 171090 242308 171096
rect 242164 167136 242216 167142
rect 242164 167078 242216 167084
rect 241796 167000 241848 167006
rect 241796 166942 241848 166948
rect 241704 161424 241756 161430
rect 241704 161366 241756 161372
rect 241152 154624 241204 154630
rect 241152 154566 241204 154572
rect 240968 140072 241020 140078
rect 240968 140014 241020 140020
rect 241060 140072 241112 140078
rect 241060 140014 241112 140020
rect 240968 116000 241020 116006
rect 240968 115942 241020 115948
rect 240876 115796 240928 115802
rect 240876 115738 240928 115744
rect 240784 114640 240836 114646
rect 240784 114582 240836 114588
rect 239588 108928 239640 108934
rect 239588 108870 239640 108876
rect 239588 104916 239640 104922
rect 239588 104858 239640 104864
rect 239600 61402 239628 104858
rect 239680 96756 239732 96762
rect 239680 96698 239732 96704
rect 239692 93838 239720 96698
rect 239680 93832 239732 93838
rect 239680 93774 239732 93780
rect 239588 61396 239640 61402
rect 239588 61338 239640 61344
rect 240414 43616 240470 43625
rect 240414 43551 240416 43560
rect 240468 43551 240470 43560
rect 240416 43522 240468 43528
rect 240796 39370 240824 114582
rect 240876 107908 240928 107914
rect 240876 107850 240928 107856
rect 240888 57322 240916 107850
rect 240980 76566 241008 115942
rect 241072 100706 241100 140014
rect 241164 116618 241192 154566
rect 242176 131034 242204 167078
rect 242268 138718 242296 171090
rect 242912 163538 242940 245618
rect 242992 202224 243044 202230
rect 242992 202166 243044 202172
rect 242900 163532 242952 163538
rect 242900 163474 242952 163480
rect 242440 156664 242492 156670
rect 242440 156606 242492 156612
rect 242348 145036 242400 145042
rect 242348 144978 242400 144984
rect 242256 138712 242308 138718
rect 242256 138654 242308 138660
rect 242164 131028 242216 131034
rect 242164 130970 242216 130976
rect 242164 124228 242216 124234
rect 242164 124170 242216 124176
rect 241152 116612 241204 116618
rect 241152 116554 241204 116560
rect 241060 100700 241112 100706
rect 241060 100642 241112 100648
rect 240968 76560 241020 76566
rect 240968 76502 241020 76508
rect 240876 57316 240928 57322
rect 240876 57258 240928 57264
rect 240784 39364 240836 39370
rect 240784 39306 240836 39312
rect 241888 35216 241940 35222
rect 241886 35184 241888 35193
rect 241940 35184 241942 35193
rect 241886 35119 241942 35128
rect 239496 32428 239548 32434
rect 239496 32370 239548 32376
rect 239404 13184 239456 13190
rect 239404 13126 239456 13132
rect 241334 11792 241390 11801
rect 241334 11727 241390 11736
rect 236736 7608 236788 7614
rect 236736 7550 236788 7556
rect 239128 4956 239180 4962
rect 239128 4898 239180 4904
rect 239140 4146 239168 4898
rect 239128 4140 239180 4146
rect 239128 4082 239180 4088
rect 239312 4140 239364 4146
rect 239312 4082 239364 4088
rect 233976 3052 234028 3058
rect 233976 2994 234028 3000
rect 235816 3052 235868 3058
rect 235816 2994 235868 3000
rect 235828 480 235856 2994
rect 239324 480 239352 4082
rect 241348 3505 241376 11727
rect 240506 3496 240562 3505
rect 240506 3431 240562 3440
rect 241334 3496 241390 3505
rect 241334 3431 241390 3440
rect 241702 3496 241758 3505
rect 241702 3431 241758 3440
rect 240520 480 240548 3431
rect 241716 480 241744 3431
rect 242176 2106 242204 124170
rect 242256 116068 242308 116074
rect 242256 116010 242308 116016
rect 242268 47598 242296 116010
rect 242360 104786 242388 144978
rect 242452 117298 242480 156606
rect 243004 155854 243032 202166
rect 244936 191418 244964 343606
rect 245016 305040 245068 305046
rect 245016 304982 245068 304988
rect 244280 191412 244332 191418
rect 244280 191354 244332 191360
rect 244924 191412 244976 191418
rect 244924 191354 244976 191360
rect 243084 184476 243136 184482
rect 243084 184418 243136 184424
rect 243096 168434 243124 184418
rect 243820 172644 243872 172650
rect 243820 172586 243872 172592
rect 243084 168428 243136 168434
rect 243084 168370 243136 168376
rect 243728 167680 243780 167686
rect 243728 167622 243780 167628
rect 242992 155848 243044 155854
rect 242992 155790 243044 155796
rect 243636 138100 243688 138106
rect 243636 138042 243688 138048
rect 243544 132524 243596 132530
rect 243544 132466 243596 132472
rect 242440 117292 242492 117298
rect 242440 117234 242492 117240
rect 242348 104780 242400 104786
rect 242348 104722 242400 104728
rect 242440 103692 242492 103698
rect 242440 103634 242492 103640
rect 242452 64190 242480 103634
rect 242440 64184 242492 64190
rect 242440 64126 242492 64132
rect 242256 47592 242308 47598
rect 242256 47534 242308 47540
rect 243556 21418 243584 132466
rect 243648 60178 243676 138042
rect 243740 128246 243768 167622
rect 243832 133822 243860 172586
rect 244292 164150 244320 191354
rect 244372 183116 244424 183122
rect 244372 183058 244424 183064
rect 244280 164144 244332 164150
rect 244280 164086 244332 164092
rect 244384 162790 244412 183058
rect 244464 181620 244516 181626
rect 244464 181562 244516 181568
rect 244476 164218 244504 181562
rect 245028 181558 245056 304982
rect 248420 259548 248472 259554
rect 248420 259490 248472 259496
rect 245660 235408 245712 235414
rect 245660 235350 245712 235356
rect 245016 181552 245068 181558
rect 245016 181494 245068 181500
rect 244924 173936 244976 173942
rect 244924 173878 244976 173884
rect 244464 164212 244516 164218
rect 244464 164154 244516 164160
rect 244372 162784 244424 162790
rect 244372 162726 244424 162732
rect 244936 135182 244964 173878
rect 245672 171086 245700 235350
rect 247040 209092 247092 209098
rect 247040 209034 247092 209040
rect 245752 191208 245804 191214
rect 245752 191150 245804 191156
rect 245660 171080 245712 171086
rect 245660 171022 245712 171028
rect 245016 163532 245068 163538
rect 245016 163474 245068 163480
rect 244924 135176 244976 135182
rect 244924 135118 244976 135124
rect 243820 133816 243872 133822
rect 243820 133758 243872 133764
rect 243728 128240 243780 128246
rect 243728 128182 243780 128188
rect 245028 126886 245056 163474
rect 245764 163198 245792 191150
rect 245844 180328 245896 180334
rect 245844 180270 245896 180276
rect 245752 163192 245804 163198
rect 245752 163134 245804 163140
rect 245856 160070 245884 180270
rect 246396 171828 246448 171834
rect 246396 171770 246448 171776
rect 246304 161560 246356 161566
rect 246304 161502 246356 161508
rect 245844 160064 245896 160070
rect 245844 160006 245896 160012
rect 245200 158840 245252 158846
rect 245200 158782 245252 158788
rect 245108 134020 245160 134026
rect 245108 133962 245160 133968
rect 245016 126880 245068 126886
rect 245016 126822 245068 126828
rect 244924 117496 244976 117502
rect 244924 117438 244976 117444
rect 243636 60172 243688 60178
rect 243636 60114 243688 60120
rect 244278 46336 244334 46345
rect 244278 46271 244280 46280
rect 244332 46271 244334 46280
rect 244280 46242 244332 46248
rect 244280 32496 244332 32502
rect 244280 32438 244332 32444
rect 243544 21412 243596 21418
rect 243544 21354 243596 21360
rect 244292 16574 244320 32438
rect 244936 29646 244964 117438
rect 245016 117428 245068 117434
rect 245016 117370 245068 117376
rect 245028 43518 245056 117370
rect 245120 68338 245148 133962
rect 245212 118590 245240 158782
rect 245292 157480 245344 157486
rect 245292 157422 245344 157428
rect 245304 118658 245332 157422
rect 246316 122738 246344 161502
rect 246408 136542 246436 171770
rect 246672 168496 246724 168502
rect 246672 168438 246724 168444
rect 246488 147756 246540 147762
rect 246488 147698 246540 147704
rect 246396 136536 246448 136542
rect 246396 136478 246448 136484
rect 246396 128376 246448 128382
rect 246396 128318 246448 128324
rect 246304 122732 246356 122738
rect 246304 122674 246356 122680
rect 246304 118720 246356 118726
rect 246304 118662 246356 118668
rect 245292 118652 245344 118658
rect 245292 118594 245344 118600
rect 245200 118584 245252 118590
rect 245200 118526 245252 118532
rect 245200 106344 245252 106350
rect 245200 106286 245252 106292
rect 245108 68332 245160 68338
rect 245108 68274 245160 68280
rect 245212 58682 245240 106286
rect 245200 58676 245252 58682
rect 245200 58618 245252 58624
rect 245016 43512 245068 43518
rect 245016 43454 245068 43460
rect 244924 29640 244976 29646
rect 244924 29582 244976 29588
rect 245752 22704 245804 22710
rect 245750 22672 245752 22681
rect 245804 22672 245806 22681
rect 245750 22607 245806 22616
rect 244292 16546 245056 16574
rect 243544 15904 243596 15910
rect 243544 15846 243596 15852
rect 242806 11792 242862 11801
rect 242806 11727 242862 11736
rect 242820 3505 242848 11727
rect 243556 4078 243584 15846
rect 242900 4072 242952 4078
rect 242900 4014 242952 4020
rect 243544 4072 243596 4078
rect 243544 4014 243596 4020
rect 242806 3496 242862 3505
rect 242806 3431 242862 3440
rect 242164 2100 242216 2106
rect 242164 2042 242216 2048
rect 242912 480 242940 4014
rect 244096 3596 244148 3602
rect 244096 3538 244148 3544
rect 244108 480 244136 3538
rect 245028 3482 245056 16546
rect 245106 11792 245162 11801
rect 245106 11727 245162 11736
rect 245120 3602 245148 11727
rect 246316 7682 246344 118662
rect 246408 43450 246436 128318
rect 246500 107574 246528 147698
rect 246580 135380 246632 135386
rect 246580 135322 246632 135328
rect 246488 107568 246540 107574
rect 246488 107510 246540 107516
rect 246488 100768 246540 100774
rect 246488 100710 246540 100716
rect 246396 43444 246448 43450
rect 246396 43386 246448 43392
rect 246500 22778 246528 100710
rect 246592 61470 246620 135322
rect 246684 129674 246712 168438
rect 247052 146198 247080 209034
rect 247132 184340 247184 184346
rect 247132 184282 247184 184288
rect 247040 146192 247092 146198
rect 247040 146134 247092 146140
rect 247144 139262 247172 184282
rect 247224 180260 247276 180266
rect 247224 180202 247276 180208
rect 247236 155922 247264 180202
rect 247868 164892 247920 164898
rect 247868 164834 247920 164840
rect 247224 155916 247276 155922
rect 247224 155858 247276 155864
rect 247132 139256 247184 139262
rect 247132 139198 247184 139204
rect 247776 138168 247828 138174
rect 247776 138110 247828 138116
rect 246672 129668 246724 129674
rect 246672 129610 246724 129616
rect 247684 128444 247736 128450
rect 247684 128386 247736 128392
rect 246580 61464 246632 61470
rect 246580 61406 246632 61412
rect 247696 44878 247724 128386
rect 247788 69766 247816 138110
rect 247880 129742 247908 164834
rect 248432 157282 248460 259490
rect 248512 205080 248564 205086
rect 248512 205022 248564 205028
rect 248420 157276 248472 157282
rect 248420 157218 248472 157224
rect 248524 154494 248552 205022
rect 249076 181694 249104 384270
rect 254584 326392 254636 326398
rect 254584 326334 254636 326340
rect 251824 301164 251876 301170
rect 251824 301106 251876 301112
rect 249800 296880 249852 296886
rect 249800 296822 249852 296828
rect 248604 181688 248656 181694
rect 248604 181630 248656 181636
rect 249064 181688 249116 181694
rect 249064 181630 249116 181636
rect 248512 154488 248564 154494
rect 248512 154430 248564 154436
rect 248616 142050 248644 181630
rect 249708 169788 249760 169794
rect 249708 169730 249760 169736
rect 249064 167204 249116 167210
rect 249064 167146 249116 167152
rect 248604 142044 248656 142050
rect 248604 141986 248656 141992
rect 247868 129736 247920 129742
rect 247868 129678 247920 129684
rect 249076 128314 249104 167146
rect 249720 167142 249748 169730
rect 249708 167136 249760 167142
rect 249708 167078 249760 167084
rect 249812 165578 249840 296822
rect 251180 280220 251232 280226
rect 251180 280162 251232 280168
rect 250444 254040 250496 254046
rect 250444 253982 250496 253988
rect 249892 207732 249944 207738
rect 249892 207674 249944 207680
rect 249800 165572 249852 165578
rect 249800 165514 249852 165520
rect 249904 151706 249932 207674
rect 250456 177546 250484 253982
rect 250444 177540 250496 177546
rect 250444 177482 250496 177488
rect 250444 174004 250496 174010
rect 250444 173946 250496 173952
rect 249892 151700 249944 151706
rect 249892 151642 249944 151648
rect 249156 150544 249208 150550
rect 249156 150486 249208 150492
rect 249064 128308 249116 128314
rect 249064 128250 249116 128256
rect 249064 121576 249116 121582
rect 249064 121518 249116 121524
rect 247868 114708 247920 114714
rect 247868 114650 247920 114656
rect 247776 69760 247828 69766
rect 247776 69702 247828 69708
rect 247880 53106 247908 114650
rect 248972 98184 249024 98190
rect 248972 98126 249024 98132
rect 248984 95946 249012 98126
rect 248972 95940 249024 95946
rect 248972 95882 249024 95888
rect 247868 53100 247920 53106
rect 247868 53042 247920 53048
rect 248512 51740 248564 51746
rect 248512 51682 248564 51688
rect 248524 48385 248552 51682
rect 248510 48376 248566 48385
rect 248510 48311 248566 48320
rect 247684 44872 247736 44878
rect 247684 44814 247736 44820
rect 248512 37936 248564 37942
rect 248510 37904 248512 37913
rect 248564 37904 248566 37913
rect 248510 37839 248566 37848
rect 246488 22772 246540 22778
rect 246488 22714 246540 22720
rect 246946 11792 247002 11801
rect 246946 11727 247002 11736
rect 246304 7676 246356 7682
rect 246304 7618 246356 7624
rect 245108 3596 245160 3602
rect 245108 3538 245160 3544
rect 246960 3505 246988 11727
rect 249076 4894 249104 121518
rect 249168 113830 249196 150486
rect 249248 149184 249300 149190
rect 249248 149126 249300 149132
rect 249156 113824 249208 113830
rect 249156 113766 249208 113772
rect 249260 112538 249288 149126
rect 250456 136610 250484 173946
rect 250536 169856 250588 169862
rect 250536 169798 250588 169804
rect 250444 136604 250496 136610
rect 250444 136546 250496 136552
rect 250444 132592 250496 132598
rect 250444 132534 250496 132540
rect 249248 112532 249300 112538
rect 249248 112474 249300 112480
rect 249156 111852 249208 111858
rect 249156 111794 249208 111800
rect 249168 51814 249196 111794
rect 249248 106412 249300 106418
rect 249248 106354 249300 106360
rect 249260 73846 249288 106354
rect 249248 73840 249300 73846
rect 249248 73782 249300 73788
rect 249156 51808 249208 51814
rect 249156 51750 249208 51756
rect 250456 18630 250484 132534
rect 250548 132326 250576 169798
rect 250628 159384 250680 159390
rect 250628 159326 250680 159332
rect 250536 132320 250588 132326
rect 250536 132262 250588 132268
rect 250536 127016 250588 127022
rect 250536 126958 250588 126964
rect 250548 50386 250576 126958
rect 250640 124098 250668 159326
rect 251192 142118 251220 280162
rect 251272 203788 251324 203794
rect 251272 203730 251324 203736
rect 251284 154562 251312 203730
rect 251364 185768 251416 185774
rect 251364 185710 251416 185716
rect 251376 156738 251404 185710
rect 251836 181762 251864 301106
rect 253940 289876 253992 289882
rect 253940 289818 253992 289824
rect 252560 225684 252612 225690
rect 252560 225626 252612 225632
rect 251824 181756 251876 181762
rect 251824 181698 251876 181704
rect 251916 169924 251968 169930
rect 251916 169866 251968 169872
rect 251364 156732 251416 156738
rect 251364 156674 251416 156680
rect 251272 154556 251324 154562
rect 251272 154498 251324 154504
rect 251180 142112 251232 142118
rect 251180 142054 251232 142060
rect 251928 131102 251956 169866
rect 252572 158710 252600 225626
rect 252652 194200 252704 194206
rect 252652 194142 252704 194148
rect 252560 158704 252612 158710
rect 252560 158646 252612 158652
rect 252100 156052 252152 156058
rect 252100 155994 252152 156000
rect 251916 131096 251968 131102
rect 251916 131038 251968 131044
rect 251824 129804 251876 129810
rect 251824 129746 251876 129752
rect 250628 124092 250680 124098
rect 250628 124034 250680 124040
rect 251180 53236 251232 53242
rect 251180 53178 251232 53184
rect 250536 50380 250588 50386
rect 250536 50322 250588 50328
rect 250444 18624 250496 18630
rect 250444 18566 250496 18572
rect 249800 17264 249852 17270
rect 249800 17206 249852 17212
rect 249812 16574 249840 17206
rect 249812 16546 250024 16574
rect 249706 15600 249762 15609
rect 249706 15535 249762 15544
rect 249064 4888 249116 4894
rect 249064 4830 249116 4836
rect 249720 3505 249748 15535
rect 246394 3496 246450 3505
rect 245028 3454 245240 3482
rect 245212 480 245240 3454
rect 246394 3431 246450 3440
rect 246946 3496 247002 3505
rect 246946 3431 247002 3440
rect 247590 3496 247646 3505
rect 247590 3431 247646 3440
rect 248786 3496 248842 3505
rect 248786 3431 248842 3440
rect 249706 3496 249762 3505
rect 249706 3431 249762 3440
rect 246408 480 246436 3431
rect 247604 480 247632 3431
rect 248800 480 248828 3431
rect 249996 480 250024 16546
rect 251192 480 251220 53178
rect 251836 33794 251864 129746
rect 252112 127634 252140 155994
rect 252192 153876 252244 153882
rect 252192 153818 252244 153824
rect 252100 127628 252152 127634
rect 252100 127570 252152 127576
rect 252008 127084 252060 127090
rect 252008 127026 252060 127032
rect 251916 113280 251968 113286
rect 251916 113222 251968 113228
rect 251824 33788 251876 33794
rect 251824 33730 251876 33736
rect 251928 31074 251956 113222
rect 252020 57254 252048 127026
rect 252204 114510 252232 153818
rect 252664 151774 252692 194142
rect 253204 165708 253256 165714
rect 253204 165650 253256 165656
rect 252652 151768 252704 151774
rect 252652 151710 252704 151716
rect 253112 143676 253164 143682
rect 253112 143618 253164 143624
rect 253124 142769 253152 143618
rect 253110 142760 253166 142769
rect 253110 142695 253166 142704
rect 253216 126954 253244 165650
rect 253296 161628 253348 161634
rect 253296 161570 253348 161576
rect 253204 126948 253256 126954
rect 253204 126890 253256 126896
rect 253308 121446 253336 161570
rect 253952 143546 253980 289818
rect 254032 178764 254084 178770
rect 254032 178706 254084 178712
rect 253940 143540 253992 143546
rect 253940 143482 253992 143488
rect 253480 142180 253532 142186
rect 253480 142122 253532 142128
rect 253388 131164 253440 131170
rect 253388 131106 253440 131112
rect 253296 121440 253348 121446
rect 253296 121382 253348 121388
rect 253204 120216 253256 120222
rect 253204 120158 253256 120164
rect 252192 114504 252244 114510
rect 252192 114446 252244 114452
rect 252100 113348 252152 113354
rect 252100 113290 252152 113296
rect 252008 57248 252060 57254
rect 252008 57190 252060 57196
rect 252112 51678 252140 113290
rect 252100 51672 252152 51678
rect 252100 51614 252152 51620
rect 251916 31068 251968 31074
rect 251916 31010 251968 31016
rect 253216 28354 253244 120158
rect 253296 107772 253348 107778
rect 253296 107714 253348 107720
rect 253204 28348 253256 28354
rect 253204 28290 253256 28296
rect 252926 24304 252982 24313
rect 252926 24239 252928 24248
rect 252980 24239 252982 24248
rect 252928 24210 252980 24216
rect 253308 18698 253336 107714
rect 253400 71058 253428 131106
rect 253492 108322 253520 142122
rect 254044 137902 254072 178706
rect 254032 137896 254084 137902
rect 254032 137838 254084 137844
rect 253480 108316 253532 108322
rect 253480 108258 253532 108264
rect 253480 102400 253532 102406
rect 253480 102342 253532 102348
rect 253388 71052 253440 71058
rect 253388 70994 253440 71000
rect 253492 46238 253520 102342
rect 254596 54534 254624 326334
rect 256700 299668 256752 299674
rect 256700 299610 256752 299616
rect 255964 266484 256016 266490
rect 255964 266426 256016 266432
rect 255976 183122 256004 266426
rect 255964 183116 256016 183122
rect 255964 183058 256016 183064
rect 256056 174072 256108 174078
rect 256056 174014 256108 174020
rect 254676 142248 254728 142254
rect 254676 142190 254728 142196
rect 254688 101454 254716 142190
rect 254768 135448 254820 135454
rect 254768 135390 254820 135396
rect 254676 101448 254728 101454
rect 254676 101390 254728 101396
rect 254676 99544 254728 99550
rect 254676 99486 254728 99492
rect 254584 54528 254636 54534
rect 254584 54470 254636 54476
rect 253480 46232 253532 46238
rect 253480 46174 253532 46180
rect 253296 18692 253348 18698
rect 253296 18634 253348 18640
rect 254596 16574 254624 54470
rect 254688 24138 254716 99486
rect 254780 62898 254808 135390
rect 256068 135250 256096 174014
rect 256712 157350 256740 299610
rect 258080 296812 258132 296818
rect 258080 296754 258132 296760
rect 257344 267776 257396 267782
rect 257344 267718 257396 267724
rect 256792 191276 256844 191282
rect 256792 191218 256844 191224
rect 256700 157344 256752 157350
rect 256700 157286 256752 157292
rect 256332 155304 256384 155310
rect 256332 155246 256384 155252
rect 256240 148368 256292 148374
rect 256240 148310 256292 148316
rect 256056 135244 256108 135250
rect 256056 135186 256108 135192
rect 255964 134088 256016 134094
rect 255964 134030 256016 134036
rect 254860 125656 254912 125662
rect 254860 125598 254912 125604
rect 254872 76634 254900 125598
rect 254860 76628 254912 76634
rect 254860 76570 254912 76576
rect 254768 62892 254820 62898
rect 254768 62834 254820 62840
rect 255318 39400 255374 39409
rect 255318 39335 255320 39344
rect 255372 39335 255374 39344
rect 255320 39306 255372 39312
rect 254676 24132 254728 24138
rect 254676 24074 254728 24080
rect 254596 16546 254716 16574
rect 253846 11792 253902 11801
rect 253846 11727 253902 11736
rect 251270 8256 251326 8265
rect 251270 8191 251272 8200
rect 251324 8191 251326 8200
rect 252376 8220 252428 8226
rect 251272 8162 251324 8168
rect 252376 8162 252428 8168
rect 252388 7614 252416 8162
rect 252376 7608 252428 7614
rect 252376 7550 252428 7556
rect 252388 480 252416 7550
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 354 253562 480
rect 253860 354 253888 11727
rect 254688 480 254716 16546
rect 255976 10334 256004 134030
rect 256148 122868 256200 122874
rect 256148 122810 256200 122816
rect 256056 116136 256108 116142
rect 256056 116078 256108 116084
rect 256068 44946 256096 116078
rect 256160 75274 256188 122810
rect 256252 107642 256280 148310
rect 256344 122806 256372 155246
rect 256804 146130 256832 191218
rect 257356 178906 257384 267718
rect 257344 178900 257396 178906
rect 257344 178842 257396 178848
rect 257344 160268 257396 160274
rect 257344 160210 257396 160216
rect 256792 146124 256844 146130
rect 256792 146066 256844 146072
rect 257356 123486 257384 160210
rect 257528 151836 257580 151842
rect 257528 151778 257580 151784
rect 257436 139528 257488 139534
rect 257436 139470 257488 139476
rect 257344 123480 257396 123486
rect 257344 123422 257396 123428
rect 256332 122800 256384 122806
rect 256332 122742 256384 122748
rect 257344 121644 257396 121650
rect 257344 121586 257396 121592
rect 256240 107636 256292 107642
rect 256240 107578 256292 107584
rect 256240 104984 256292 104990
rect 256240 104926 256292 104932
rect 256148 75268 256200 75274
rect 256148 75210 256200 75216
rect 256252 54602 256280 104926
rect 256240 54596 256292 54602
rect 256240 54538 256292 54544
rect 256056 44940 256108 44946
rect 256056 44882 256108 44888
rect 257356 14550 257384 121586
rect 257448 56030 257476 139470
rect 257540 110430 257568 151778
rect 258092 137970 258120 296754
rect 259460 253972 259512 253978
rect 259460 253914 259512 253920
rect 258724 244384 258776 244390
rect 258724 244326 258776 244332
rect 258736 180266 258764 244326
rect 258724 180260 258776 180266
rect 258724 180202 258776 180208
rect 258724 171352 258776 171358
rect 258724 171294 258776 171300
rect 258080 137964 258132 137970
rect 258080 137906 258132 137912
rect 258736 132394 258764 171294
rect 259000 169516 259052 169522
rect 259000 169458 259052 169464
rect 259012 132462 259040 169458
rect 259472 150414 259500 253914
rect 260116 177313 260144 393314
rect 262864 389224 262916 389230
rect 262864 389166 262916 389172
rect 260840 291304 260892 291310
rect 260840 291246 260892 291252
rect 260196 220108 260248 220114
rect 260196 220050 260248 220056
rect 260102 177304 260158 177313
rect 260102 177239 260158 177248
rect 260208 176662 260236 220050
rect 260196 176656 260248 176662
rect 260196 176598 260248 176604
rect 260104 172712 260156 172718
rect 260104 172654 260156 172660
rect 259460 150408 259512 150414
rect 259460 150350 259512 150356
rect 259184 140956 259236 140962
rect 259184 140898 259236 140904
rect 259092 133204 259144 133210
rect 259092 133146 259144 133152
rect 259000 132456 259052 132462
rect 259000 132398 259052 132404
rect 258724 132388 258776 132394
rect 258724 132330 258776 132336
rect 258816 131300 258868 131306
rect 258816 131242 258868 131248
rect 258724 118788 258776 118794
rect 258724 118730 258776 118736
rect 257528 110424 257580 110430
rect 257528 110366 257580 110372
rect 257620 109200 257672 109206
rect 257620 109142 257672 109148
rect 257528 100836 257580 100842
rect 257528 100778 257580 100784
rect 257436 56024 257488 56030
rect 257436 55966 257488 55972
rect 257540 25566 257568 100778
rect 257632 35290 257660 109142
rect 257620 35284 257672 35290
rect 257620 35226 257672 35232
rect 257528 25560 257580 25566
rect 257528 25502 257580 25508
rect 257344 14544 257396 14550
rect 257344 14486 257396 14492
rect 256330 11792 256386 11801
rect 256330 11727 256386 11736
rect 255964 10328 256016 10334
rect 255964 10270 256016 10276
rect 253450 326 253888 354
rect 253450 -960 253562 326
rect 254646 -960 254758 480
rect 255842 354 255954 480
rect 256344 354 256372 11727
rect 258446 10976 258502 10985
rect 258446 10911 258448 10920
rect 258500 10911 258502 10920
rect 258448 10882 258500 10888
rect 256700 7744 256752 7750
rect 256700 7686 256752 7692
rect 256712 5506 256740 7686
rect 256700 5500 256752 5506
rect 256700 5442 256752 5448
rect 257068 5500 257120 5506
rect 257068 5442 257120 5448
rect 257080 480 257108 5442
rect 258736 4826 258764 118730
rect 258828 49026 258856 131242
rect 258908 131232 258960 131238
rect 258908 131174 258960 131180
rect 258920 55962 258948 131174
rect 259104 101998 259132 133146
rect 259196 119406 259224 140898
rect 260116 133890 260144 172654
rect 260196 162988 260248 162994
rect 260196 162930 260248 162936
rect 260104 133884 260156 133890
rect 260104 133826 260156 133832
rect 260208 124166 260236 162930
rect 260852 153202 260880 291246
rect 261576 157548 261628 157554
rect 261576 157490 261628 157496
rect 260840 153196 260892 153202
rect 260840 153138 260892 153144
rect 260378 146432 260434 146441
rect 260378 146367 260434 146376
rect 260196 124160 260248 124166
rect 260196 124102 260248 124108
rect 260104 122936 260156 122942
rect 260104 122878 260156 122884
rect 259184 119400 259236 119406
rect 259184 119342 259236 119348
rect 259092 101992 259144 101998
rect 259092 101934 259144 101940
rect 259000 100904 259052 100910
rect 259000 100846 259052 100852
rect 258908 55956 258960 55962
rect 258908 55898 258960 55904
rect 258816 49020 258868 49026
rect 258816 48962 258868 48968
rect 259012 26926 259040 100846
rect 259460 50380 259512 50386
rect 259460 50322 259512 50328
rect 259000 26920 259052 26926
rect 259000 26862 259052 26868
rect 259368 10940 259420 10946
rect 259368 10882 259420 10888
rect 259380 10334 259408 10882
rect 259368 10328 259420 10334
rect 259368 10270 259420 10276
rect 258724 4820 258776 4826
rect 258724 4762 258776 4768
rect 259380 3505 259408 10270
rect 258262 3496 258318 3505
rect 258262 3431 258318 3440
rect 259366 3496 259422 3505
rect 259366 3431 259422 3440
rect 258276 480 258304 3431
rect 259472 480 259500 50322
rect 259552 26920 259604 26926
rect 259552 26862 259604 26868
rect 259564 6914 259592 26862
rect 260116 13122 260144 122878
rect 260196 120284 260248 120290
rect 260196 120226 260248 120232
rect 260208 19990 260236 120226
rect 260288 110492 260340 110498
rect 260288 110434 260340 110440
rect 260300 53174 260328 110434
rect 260392 109002 260420 146367
rect 260930 136640 260986 136649
rect 260930 136575 260986 136584
rect 260944 135318 260972 136575
rect 261114 136232 261170 136241
rect 261114 136167 261170 136176
rect 261128 135386 261156 136167
rect 261116 135380 261168 135386
rect 261116 135322 261168 135328
rect 260932 135312 260984 135318
rect 260932 135254 260984 135260
rect 261484 123140 261536 123146
rect 261484 123082 261536 123088
rect 260380 108996 260432 109002
rect 260380 108938 260432 108944
rect 261390 97880 261446 97889
rect 261390 97815 261446 97824
rect 260380 96756 260432 96762
rect 260380 96698 260432 96704
rect 260392 75206 260420 96698
rect 261404 96694 261432 97815
rect 261392 96688 261444 96694
rect 261392 96630 261444 96636
rect 260380 75200 260432 75206
rect 260380 75142 260432 75148
rect 260288 53168 260340 53174
rect 260288 53110 260340 53116
rect 260196 19984 260248 19990
rect 260196 19926 260248 19932
rect 260104 13116 260156 13122
rect 260104 13058 260156 13064
rect 261496 9042 261524 123082
rect 261588 120086 261616 157490
rect 261850 146160 261906 146169
rect 261850 146095 261906 146104
rect 261668 135516 261720 135522
rect 261668 135458 261720 135464
rect 261576 120080 261628 120086
rect 261576 120022 261628 120028
rect 261576 107840 261628 107846
rect 261576 107782 261628 107788
rect 261588 21486 261616 107782
rect 261680 65550 261708 135458
rect 261864 106282 261892 146095
rect 262876 106282 262904 389166
rect 282184 363656 282236 363662
rect 282184 363598 282236 363604
rect 269764 336048 269816 336054
rect 269764 335990 269816 335996
rect 268384 325032 268436 325038
rect 268384 324974 268436 324980
rect 267004 320952 267056 320958
rect 267004 320894 267056 320900
rect 265624 318164 265676 318170
rect 265624 318106 265676 318112
rect 264244 311908 264296 311914
rect 264244 311850 264296 311856
rect 262956 308508 263008 308514
rect 262956 308450 263008 308456
rect 262968 182986 262996 308450
rect 264256 185774 264284 311850
rect 264336 250572 264388 250578
rect 264336 250514 264388 250520
rect 264244 185768 264296 185774
rect 264244 185710 264296 185716
rect 262956 182980 263008 182986
rect 262956 182922 263008 182928
rect 264348 181626 264376 250514
rect 265636 183054 265664 318106
rect 265624 183048 265676 183054
rect 265624 182990 265676 182996
rect 264336 181620 264388 181626
rect 264336 181562 264388 181568
rect 264426 175400 264482 175409
rect 264426 175335 264482 175344
rect 263140 165776 263192 165782
rect 263140 165718 263192 165724
rect 263046 164928 263102 164937
rect 263046 164863 263102 164872
rect 262954 137456 263010 137465
rect 262954 137391 263010 137400
rect 261852 106276 261904 106282
rect 261852 106218 261904 106224
rect 262864 106276 262916 106282
rect 262864 106218 262916 106224
rect 261760 105052 261812 105058
rect 261760 104994 261812 105000
rect 261668 65544 261720 65550
rect 261668 65486 261720 65492
rect 261772 60110 261800 104994
rect 262864 103760 262916 103766
rect 262864 103702 262916 103708
rect 261760 60104 261812 60110
rect 261760 60046 261812 60052
rect 262220 42152 262272 42158
rect 262220 42094 262272 42100
rect 261576 21480 261628 21486
rect 261576 21422 261628 21428
rect 262232 16574 262260 42094
rect 262876 42090 262904 103702
rect 262864 42084 262916 42090
rect 262864 42026 262916 42032
rect 262232 16546 262536 16574
rect 261760 13252 261812 13258
rect 261760 13194 261812 13200
rect 261484 9036 261536 9042
rect 261484 8978 261536 8984
rect 259564 6886 260696 6914
rect 260668 480 260696 6886
rect 261772 480 261800 13194
rect 255842 326 256372 354
rect 255842 -960 255954 326
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 262968 15978 262996 137391
rect 263060 125526 263088 164863
rect 263152 130422 263180 165718
rect 264242 165064 264298 165073
rect 264242 164999 264298 165008
rect 263140 130416 263192 130422
rect 263140 130358 263192 130364
rect 264256 125594 264284 164999
rect 264334 145344 264390 145353
rect 264334 145279 264390 145288
rect 264244 125588 264296 125594
rect 264244 125530 264296 125536
rect 263048 125520 263100 125526
rect 263048 125462 263100 125468
rect 263138 122632 263194 122641
rect 263138 122567 263194 122576
rect 263048 107704 263100 107710
rect 263048 107646 263100 107652
rect 263060 47666 263088 107646
rect 263152 69698 263180 122567
rect 264244 121644 264296 121650
rect 264244 121586 264296 121592
rect 264256 121281 264284 121586
rect 264242 121272 264298 121281
rect 264242 121207 264298 121216
rect 264348 112470 264376 145279
rect 264440 142866 264468 175335
rect 265898 174992 265954 175001
rect 265898 174927 265954 174936
rect 265346 174176 265402 174185
rect 265346 174111 265402 174120
rect 265360 174078 265388 174111
rect 265348 174072 265400 174078
rect 265348 174014 265400 174020
rect 265806 174040 265862 174049
rect 265912 174010 265940 174927
rect 265990 174584 266046 174593
rect 265990 174519 266046 174528
rect 265806 173975 265862 173984
rect 265900 174004 265952 174010
rect 265820 173942 265848 173975
rect 265900 173946 265952 173952
rect 265808 173936 265860 173942
rect 265808 173878 265860 173884
rect 265254 173224 265310 173233
rect 265254 173159 265310 173168
rect 265268 172582 265296 173159
rect 265346 172816 265402 172825
rect 265346 172751 265402 172760
rect 265360 172718 265388 172751
rect 265348 172712 265400 172718
rect 265348 172654 265400 172660
rect 265808 172644 265860 172650
rect 265808 172586 265860 172592
rect 265256 172576 265308 172582
rect 265820 172553 265848 172586
rect 265256 172518 265308 172524
rect 265806 172544 265862 172553
rect 265806 172479 265862 172488
rect 265070 172000 265126 172009
rect 265070 171935 265126 171944
rect 265084 171154 265112 171935
rect 266004 171834 266032 174519
rect 265992 171828 266044 171834
rect 265992 171770 266044 171776
rect 265162 171592 265218 171601
rect 265162 171527 265218 171536
rect 265176 171358 265204 171527
rect 265164 171352 265216 171358
rect 265164 171294 265216 171300
rect 265346 171184 265402 171193
rect 265072 171148 265124 171154
rect 265346 171119 265402 171128
rect 265072 171090 265124 171096
rect 265254 170232 265310 170241
rect 265254 170167 265310 170176
rect 265268 169930 265296 170167
rect 265256 169924 265308 169930
rect 265256 169866 265308 169872
rect 265360 169522 265388 171119
rect 265438 170640 265494 170649
rect 265438 170575 265494 170584
rect 265452 169862 265480 170575
rect 265440 169856 265492 169862
rect 265440 169798 265492 169804
rect 265622 169824 265678 169833
rect 265622 169759 265624 169768
rect 265676 169759 265678 169768
rect 265624 169730 265676 169736
rect 265348 169516 265400 169522
rect 265348 169458 265400 169464
rect 265898 169416 265954 169425
rect 265898 169351 265954 169360
rect 265438 169008 265494 169017
rect 265438 168943 265494 168952
rect 265346 168600 265402 168609
rect 265346 168535 265402 168544
rect 265360 168502 265388 168535
rect 265348 168496 265400 168502
rect 265348 168438 265400 168444
rect 265254 167648 265310 167657
rect 265254 167583 265310 167592
rect 265268 167210 265296 167583
rect 265256 167204 265308 167210
rect 265256 167146 265308 167152
rect 265162 167104 265218 167113
rect 265162 167039 265218 167048
rect 265176 163538 265204 167039
rect 265452 164898 265480 168943
rect 265806 168464 265862 168473
rect 265912 168434 265940 169351
rect 265806 168399 265862 168408
rect 265900 168428 265952 168434
rect 265820 167686 265848 168399
rect 265900 168370 265952 168376
rect 265808 167680 265860 167686
rect 265808 167622 265860 167628
rect 265530 167240 265586 167249
rect 265530 167175 265586 167184
rect 265544 167074 265572 167175
rect 265532 167068 265584 167074
rect 265532 167010 265584 167016
rect 265622 166424 265678 166433
rect 265622 166359 265678 166368
rect 265636 165714 265664 166359
rect 265898 166016 265954 166025
rect 265898 165951 265954 165960
rect 265808 165776 265860 165782
rect 265806 165744 265808 165753
rect 265860 165744 265862 165753
rect 265624 165708 265676 165714
rect 265806 165679 265862 165688
rect 265624 165650 265676 165656
rect 265912 165646 265940 165951
rect 265900 165640 265952 165646
rect 265900 165582 265952 165588
rect 265440 164892 265492 164898
rect 265440 164834 265492 164840
rect 265990 163840 266046 163849
rect 265990 163775 266046 163784
rect 265164 163532 265216 163538
rect 265164 163474 265216 163480
rect 265622 163432 265678 163441
rect 265622 163367 265678 163376
rect 265530 163024 265586 163033
rect 265636 162994 265664 163367
rect 265530 162959 265586 162968
rect 265624 162988 265676 162994
rect 265544 162926 265572 162959
rect 265624 162930 265676 162936
rect 265532 162920 265584 162926
rect 265438 162888 265494 162897
rect 265532 162862 265584 162868
rect 265438 162823 265494 162832
rect 264520 161628 264572 161634
rect 264520 161570 264572 161576
rect 264532 161265 264560 161570
rect 264518 161256 264574 161265
rect 264518 161191 264574 161200
rect 265346 160848 265402 160857
rect 265346 160783 265402 160792
rect 265360 160206 265388 160783
rect 265348 160200 265400 160206
rect 265348 160142 265400 160148
rect 265162 157448 265218 157457
rect 265162 157383 265218 157392
rect 265176 156670 265204 157383
rect 265452 157334 265480 162823
rect 265714 162072 265770 162081
rect 265714 162007 265770 162016
rect 265728 161566 265756 162007
rect 265806 161664 265862 161673
rect 265806 161599 265862 161608
rect 265716 161560 265768 161566
rect 265716 161502 265768 161508
rect 265820 161498 265848 161599
rect 265808 161492 265860 161498
rect 265808 161434 265860 161440
rect 265622 160440 265678 160449
rect 265622 160375 265678 160384
rect 265636 160274 265664 160375
rect 265624 160268 265676 160274
rect 265624 160210 265676 160216
rect 265806 160168 265862 160177
rect 265806 160103 265808 160112
rect 265860 160103 265862 160112
rect 265808 160074 265860 160080
rect 265898 159488 265954 159497
rect 265898 159423 265954 159432
rect 265806 159080 265862 159089
rect 265806 159015 265862 159024
rect 265820 158846 265848 159015
rect 265808 158840 265860 158846
rect 265714 158808 265770 158817
rect 265808 158782 265860 158788
rect 265714 158743 265716 158752
rect 265768 158743 265770 158752
rect 265716 158714 265768 158720
rect 265714 158264 265770 158273
rect 265714 158199 265770 158208
rect 265622 157856 265678 157865
rect 265622 157791 265678 157800
rect 265636 157418 265664 157791
rect 265728 157486 265756 158199
rect 265912 157554 265940 159423
rect 266004 159390 266032 163775
rect 265992 159384 266044 159390
rect 265992 159326 266044 159332
rect 265900 157548 265952 157554
rect 265900 157490 265952 157496
rect 265716 157480 265768 157486
rect 265716 157422 265768 157428
rect 265624 157412 265676 157418
rect 265624 157354 265676 157360
rect 265360 157306 265480 157334
rect 265164 156664 265216 156670
rect 265164 156606 265216 156612
rect 265360 155310 265388 157306
rect 265530 156904 265586 156913
rect 265530 156839 265586 156848
rect 265544 156058 265572 156839
rect 265898 156496 265954 156505
rect 265898 156431 265954 156440
rect 265532 156052 265584 156058
rect 265532 155994 265584 156000
rect 265912 155990 265940 156431
rect 265990 156088 266046 156097
rect 265990 156023 266046 156032
rect 265900 155984 265952 155990
rect 265900 155926 265952 155932
rect 265530 155680 265586 155689
rect 265530 155615 265586 155624
rect 265348 155304 265400 155310
rect 265348 155246 265400 155252
rect 265254 149696 265310 149705
rect 265254 149631 265310 149640
rect 265268 149190 265296 149631
rect 265256 149184 265308 149190
rect 265256 149126 265308 149132
rect 265438 148336 265494 148345
rect 265438 148271 265494 148280
rect 265070 147928 265126 147937
rect 265070 147863 265126 147872
rect 265084 146985 265112 147863
rect 265452 147694 265480 148271
rect 265440 147688 265492 147694
rect 265440 147630 265492 147636
rect 265070 146976 265126 146985
rect 265070 146911 265126 146920
rect 265438 146568 265494 146577
rect 265438 146503 265494 146512
rect 264520 143744 264572 143750
rect 264520 143686 264572 143692
rect 264428 142860 264480 142866
rect 264428 142802 264480 142808
rect 264426 141536 264482 141545
rect 264426 141471 264482 141480
rect 264440 140894 264468 141471
rect 264428 140888 264480 140894
rect 264428 140830 264480 140836
rect 264426 138272 264482 138281
rect 264426 138207 264482 138216
rect 264440 138174 264468 138207
rect 264428 138168 264480 138174
rect 264428 138110 264480 138116
rect 264426 137864 264482 137873
rect 264426 137799 264482 137808
rect 264440 136678 264468 137799
rect 264428 136672 264480 136678
rect 264428 136614 264480 136620
rect 264426 135960 264482 135969
rect 264426 135895 264482 135904
rect 264440 135454 264468 135895
rect 264428 135448 264480 135454
rect 264428 135390 264480 135396
rect 264428 128444 264480 128450
rect 264428 128386 264480 128392
rect 264440 128217 264468 128386
rect 264426 128208 264482 128217
rect 264426 128143 264482 128152
rect 264428 127016 264480 127022
rect 264428 126958 264480 126964
rect 264440 126857 264468 126958
rect 264426 126848 264482 126857
rect 264426 126783 264482 126792
rect 264426 124672 264482 124681
rect 264426 124607 264482 124616
rect 264336 112464 264388 112470
rect 264336 112406 264388 112412
rect 264242 112160 264298 112169
rect 264242 112095 264298 112104
rect 263140 69692 263192 69698
rect 263140 69634 263192 69640
rect 263048 47660 263100 47666
rect 263048 47602 263100 47608
rect 264256 31142 264284 112095
rect 264334 110936 264390 110945
rect 264334 110871 264390 110880
rect 264348 39438 264376 110871
rect 264440 58750 264468 124607
rect 264532 111790 264560 143686
rect 264612 140956 264664 140962
rect 264612 140898 264664 140904
rect 264624 140593 264652 140898
rect 264610 140584 264666 140593
rect 264610 140519 264666 140528
rect 265254 139768 265310 139777
rect 265254 139703 265310 139712
rect 265268 139534 265296 139703
rect 265256 139528 265308 139534
rect 265256 139470 265308 139476
rect 265452 138938 265480 146503
rect 265544 145586 265572 155615
rect 265806 155272 265862 155281
rect 266004 155242 266032 156023
rect 265806 155207 265862 155216
rect 265992 155236 266044 155242
rect 265820 154630 265848 155207
rect 265992 155178 266044 155184
rect 265990 154728 266046 154737
rect 265990 154663 266046 154672
rect 265808 154624 265860 154630
rect 265714 154592 265770 154601
rect 265808 154566 265860 154572
rect 265714 154527 265770 154536
rect 265728 152522 265756 154527
rect 265898 153912 265954 153921
rect 266004 153882 266032 154663
rect 265898 153847 265954 153856
rect 265992 153876 266044 153882
rect 265806 153504 265862 153513
rect 265806 153439 265862 153448
rect 265820 153338 265848 153439
rect 265808 153332 265860 153338
rect 265808 153274 265860 153280
rect 265912 153270 265940 153847
rect 265992 153818 266044 153824
rect 265900 153264 265952 153270
rect 265806 153232 265862 153241
rect 265900 153206 265952 153212
rect 265806 153167 265862 153176
rect 265716 152516 265768 152522
rect 265716 152458 265768 152464
rect 265820 152425 265848 153167
rect 266082 152688 266138 152697
rect 266082 152623 266138 152632
rect 265806 152416 265862 152425
rect 265806 152351 265862 152360
rect 265990 152144 266046 152153
rect 265990 152079 266046 152088
rect 265806 151872 265862 151881
rect 265806 151807 265808 151816
rect 265860 151807 265862 151816
rect 265808 151778 265860 151784
rect 265898 151328 265954 151337
rect 265898 151263 265954 151272
rect 265806 150920 265862 150929
rect 265806 150855 265862 150864
rect 265820 150550 265848 150855
rect 265808 150544 265860 150550
rect 265808 150486 265860 150492
rect 265912 150482 265940 151263
rect 265900 150476 265952 150482
rect 265900 150418 265952 150424
rect 265898 150104 265954 150113
rect 265898 150039 265954 150048
rect 265806 149152 265862 149161
rect 265912 149122 265940 150039
rect 266004 149734 266032 152079
rect 265992 149728 266044 149734
rect 265992 149670 266044 149676
rect 265806 149087 265862 149096
rect 265900 149116 265952 149122
rect 265714 148744 265770 148753
rect 265714 148679 265770 148688
rect 265728 147762 265756 148679
rect 265820 148374 265848 149087
rect 265900 149058 265952 149064
rect 265808 148368 265860 148374
rect 265808 148310 265860 148316
rect 265716 147756 265768 147762
rect 265716 147698 265768 147704
rect 265714 147112 265770 147121
rect 265714 147047 265770 147056
rect 265728 146334 265756 147047
rect 265716 146328 265768 146334
rect 265716 146270 265768 146276
rect 265898 145752 265954 145761
rect 265898 145687 265954 145696
rect 265532 145580 265584 145586
rect 265532 145522 265584 145528
rect 265808 145104 265860 145110
rect 265808 145046 265860 145052
rect 265820 144945 265848 145046
rect 265912 145042 265940 145687
rect 265900 145036 265952 145042
rect 265900 144978 265952 144984
rect 265806 144936 265862 144945
rect 265806 144871 265862 144880
rect 265530 144528 265586 144537
rect 265530 144463 265586 144472
rect 265544 143682 265572 144463
rect 265714 143984 265770 143993
rect 265714 143919 265770 143928
rect 265532 143676 265584 143682
rect 265532 143618 265584 143624
rect 265728 142934 265756 143919
rect 266096 143750 266124 152623
rect 266174 146704 266230 146713
rect 266174 146639 266230 146648
rect 266084 143744 266136 143750
rect 266084 143686 266136 143692
rect 265808 143608 265860 143614
rect 265806 143576 265808 143585
rect 265860 143576 265862 143585
rect 265806 143511 265862 143520
rect 266082 143168 266138 143177
rect 266082 143103 266138 143112
rect 265716 142928 265768 142934
rect 265716 142870 265768 142876
rect 265530 142760 265586 142769
rect 265530 142695 265586 142704
rect 265544 142254 265572 142695
rect 265622 142352 265678 142361
rect 265622 142287 265678 142296
rect 265532 142248 265584 142254
rect 265532 142190 265584 142196
rect 265636 142186 265664 142287
rect 265714 142216 265770 142225
rect 265624 142180 265676 142186
rect 265714 142151 265770 142160
rect 265624 142122 265676 142128
rect 265728 140078 265756 142151
rect 265806 140992 265862 141001
rect 265806 140927 265862 140936
rect 265820 140826 265848 140927
rect 265808 140820 265860 140826
rect 265808 140762 265860 140768
rect 265898 140176 265954 140185
rect 265898 140111 265954 140120
rect 265716 140072 265768 140078
rect 265716 140014 265768 140020
rect 265716 139936 265768 139942
rect 265716 139878 265768 139884
rect 265452 138910 265572 138938
rect 265438 138816 265494 138825
rect 265438 138751 265494 138760
rect 265162 138408 265218 138417
rect 265162 138343 265218 138352
rect 265176 138106 265204 138343
rect 265164 138100 265216 138106
rect 265164 138042 265216 138048
rect 265452 138038 265480 138751
rect 265440 138032 265492 138038
rect 265544 138014 265572 138910
rect 265544 137986 265664 138014
rect 265440 137974 265492 137980
rect 265532 134020 265584 134026
rect 265532 133962 265584 133968
rect 265544 133929 265572 133962
rect 265530 133920 265586 133929
rect 265530 133855 265586 133864
rect 265440 131232 265492 131238
rect 265438 131200 265440 131209
rect 265492 131200 265494 131209
rect 265438 131135 265494 131144
rect 265254 130248 265310 130257
rect 265254 130183 265310 130192
rect 265268 129810 265296 130183
rect 265256 129804 265308 129810
rect 265256 129746 265308 129752
rect 265636 124302 265664 137986
rect 265728 137290 265756 139878
rect 265912 139466 265940 140111
rect 265900 139460 265952 139466
rect 265900 139402 265952 139408
rect 266096 138014 266124 143103
rect 266188 139942 266216 146639
rect 266176 139936 266228 139942
rect 266176 139878 266228 139884
rect 266004 137986 266124 138014
rect 265716 137284 265768 137290
rect 265716 137226 265768 137232
rect 265808 135516 265860 135522
rect 265808 135458 265860 135464
rect 265820 135425 265848 135458
rect 265806 135416 265862 135425
rect 265806 135351 265862 135360
rect 265806 134600 265862 134609
rect 265806 134535 265862 134544
rect 265714 134192 265770 134201
rect 265714 134127 265770 134136
rect 265728 134094 265756 134127
rect 265716 134088 265768 134094
rect 265716 134030 265768 134036
rect 265820 133958 265848 134535
rect 265808 133952 265860 133958
rect 265808 133894 265860 133900
rect 265898 133240 265954 133249
rect 266004 133210 266032 137986
rect 266082 137048 266138 137057
rect 266082 136983 266138 136992
rect 265898 133175 265954 133184
rect 265992 133204 266044 133210
rect 265714 132832 265770 132841
rect 265714 132767 265770 132776
rect 265728 132530 265756 132767
rect 265912 132598 265940 133175
rect 265992 133146 266044 133152
rect 265900 132592 265952 132598
rect 265806 132560 265862 132569
rect 265716 132524 265768 132530
rect 265900 132534 265952 132540
rect 265806 132495 265862 132504
rect 265716 132466 265768 132472
rect 265714 131608 265770 131617
rect 265714 131543 265770 131552
rect 265728 131306 265756 131543
rect 265716 131300 265768 131306
rect 265716 131242 265768 131248
rect 265714 128616 265770 128625
rect 265714 128551 265770 128560
rect 265728 128382 265756 128551
rect 265716 128376 265768 128382
rect 265716 128318 265768 128324
rect 264612 124296 264664 124302
rect 264612 124238 264664 124244
rect 265624 124296 265676 124302
rect 265624 124238 265676 124244
rect 264520 111784 264572 111790
rect 264520 111726 264572 111732
rect 264624 104854 264652 124238
rect 265622 120864 265678 120873
rect 265622 120799 265678 120808
rect 265530 120456 265586 120465
rect 265530 120391 265586 120400
rect 265544 120290 265572 120391
rect 265532 120284 265584 120290
rect 265532 120226 265584 120232
rect 265636 120154 265664 120799
rect 265716 120216 265768 120222
rect 265714 120184 265716 120193
rect 265768 120184 265770 120193
rect 265624 120148 265676 120154
rect 265714 120119 265770 120128
rect 265624 120090 265676 120096
rect 265622 119504 265678 119513
rect 265622 119439 265678 119448
rect 265636 118726 265664 119439
rect 265714 118824 265770 118833
rect 265714 118759 265716 118768
rect 265768 118759 265770 118768
rect 265716 118730 265768 118736
rect 265624 118720 265676 118726
rect 265624 118662 265676 118668
rect 265346 117872 265402 117881
rect 265346 117807 265402 117816
rect 265360 117366 265388 117807
rect 265714 117464 265770 117473
rect 265714 117399 265716 117408
rect 265768 117399 265770 117408
rect 265716 117370 265768 117376
rect 265348 117360 265400 117366
rect 265348 117302 265400 117308
rect 265622 117328 265678 117337
rect 265622 117263 265678 117272
rect 265254 115288 265310 115297
rect 265254 115223 265310 115232
rect 265268 114578 265296 115223
rect 265256 114572 265308 114578
rect 265256 114514 265308 114520
rect 265254 113928 265310 113937
rect 265254 113863 265310 113872
rect 265268 113286 265296 113863
rect 265256 113280 265308 113286
rect 265256 113222 265308 113228
rect 265162 109712 265218 109721
rect 265162 109647 265218 109656
rect 265176 109138 265204 109647
rect 265530 109304 265586 109313
rect 265530 109239 265586 109248
rect 265164 109132 265216 109138
rect 265164 109074 265216 109080
rect 265544 109070 265572 109239
rect 265532 109064 265584 109070
rect 265532 109006 265584 109012
rect 265162 108760 265218 108769
rect 265162 108695 265218 108704
rect 265176 107710 265204 108695
rect 265164 107704 265216 107710
rect 265164 107646 265216 107652
rect 265530 106720 265586 106729
rect 265530 106655 265586 106664
rect 265544 106418 265572 106655
rect 265532 106412 265584 106418
rect 265532 106354 265584 106360
rect 265530 105768 265586 105777
rect 265530 105703 265586 105712
rect 265544 105058 265572 105703
rect 265532 105052 265584 105058
rect 265532 104994 265584 105000
rect 264612 104848 264664 104854
rect 264612 104790 264664 104796
rect 264518 104544 264574 104553
rect 264518 104479 264574 104488
rect 264532 62830 264560 104479
rect 265162 102776 265218 102785
rect 265162 102711 265218 102720
rect 264612 102400 264664 102406
rect 264612 102342 264664 102348
rect 264624 101969 264652 102342
rect 265176 102202 265204 102711
rect 265164 102196 265216 102202
rect 265164 102138 265216 102144
rect 264610 101960 264666 101969
rect 264610 101895 264666 101904
rect 265346 101416 265402 101425
rect 265346 101351 265402 101360
rect 265360 100842 265388 101351
rect 265530 100872 265586 100881
rect 265348 100836 265400 100842
rect 265530 100807 265586 100816
rect 265348 100778 265400 100784
rect 265544 100774 265572 100807
rect 265532 100768 265584 100774
rect 265532 100710 265584 100716
rect 265532 99544 265584 99550
rect 265530 99512 265532 99521
rect 265584 99512 265586 99521
rect 265530 99447 265586 99456
rect 265636 99374 265664 117263
rect 265714 116104 265770 116113
rect 265714 116039 265770 116048
rect 265728 116006 265756 116039
rect 265716 116000 265768 116006
rect 265716 115942 265768 115948
rect 265714 114744 265770 114753
rect 265714 114679 265770 114688
rect 265728 114646 265756 114679
rect 265716 114640 265768 114646
rect 265716 114582 265768 114588
rect 265714 113520 265770 113529
rect 265714 113455 265770 113464
rect 265728 113354 265756 113455
rect 265716 113348 265768 113354
rect 265716 113290 265768 113296
rect 265714 113248 265770 113257
rect 265714 113183 265716 113192
rect 265768 113183 265770 113192
rect 265716 113154 265768 113160
rect 265714 111888 265770 111897
rect 265714 111823 265716 111832
rect 265768 111823 265770 111832
rect 265716 111794 265768 111800
rect 265714 110528 265770 110537
rect 265714 110463 265716 110472
rect 265768 110463 265770 110472
rect 265716 110434 265768 110440
rect 265714 110120 265770 110129
rect 265714 110055 265770 110064
rect 265728 109206 265756 110055
rect 265716 109200 265768 109206
rect 265716 109142 265768 109148
rect 265714 107944 265770 107953
rect 265714 107879 265716 107888
rect 265768 107879 265770 107888
rect 265716 107850 265768 107856
rect 265716 107772 265768 107778
rect 265716 107714 265768 107720
rect 265728 107681 265756 107714
rect 265714 107672 265770 107681
rect 265714 107607 265770 107616
rect 265714 106584 265770 106593
rect 265714 106519 265770 106528
rect 265728 106350 265756 106519
rect 265716 106344 265768 106350
rect 265716 106286 265768 106292
rect 265714 105360 265770 105369
rect 265714 105295 265770 105304
rect 265728 104922 265756 105295
rect 265716 104916 265768 104922
rect 265716 104858 265768 104864
rect 265714 104000 265770 104009
rect 265714 103935 265770 103944
rect 265728 103698 265756 103935
rect 265716 103692 265768 103698
rect 265716 103634 265768 103640
rect 265714 102368 265770 102377
rect 265714 102303 265770 102312
rect 265728 102270 265756 102303
rect 265716 102264 265768 102270
rect 265716 102206 265768 102212
rect 265714 101008 265770 101017
rect 265714 100943 265770 100952
rect 265728 100910 265756 100943
rect 265716 100904 265768 100910
rect 265716 100846 265768 100852
rect 265714 100192 265770 100201
rect 265714 100127 265770 100136
rect 265728 99482 265756 100127
rect 265716 99476 265768 99482
rect 265716 99418 265768 99424
rect 265636 99346 265756 99374
rect 265622 98424 265678 98433
rect 265622 98359 265678 98368
rect 264610 98288 264666 98297
rect 264610 98223 264666 98232
rect 264624 98122 264652 98223
rect 264612 98116 264664 98122
rect 264612 98058 264664 98064
rect 265636 98054 265664 98359
rect 265624 98048 265676 98054
rect 265624 97990 265676 97996
rect 264610 97472 264666 97481
rect 264610 97407 264666 97416
rect 264624 96762 264652 97407
rect 265622 97064 265678 97073
rect 265622 96999 265678 97008
rect 264612 96756 264664 96762
rect 264612 96698 264664 96704
rect 265530 95704 265586 95713
rect 265530 95639 265586 95648
rect 265544 95266 265572 95639
rect 265532 95260 265584 95266
rect 265532 95202 265584 95208
rect 264520 62824 264572 62830
rect 264520 62766 264572 62772
rect 264428 58744 264480 58750
rect 264428 58686 264480 58692
rect 264428 55888 264480 55894
rect 264428 55830 264480 55836
rect 264336 39432 264388 39438
rect 264336 39374 264388 39380
rect 264244 31136 264296 31142
rect 264244 31078 264296 31084
rect 263600 24200 263652 24206
rect 263600 24142 263652 24148
rect 263612 19310 263640 24142
rect 263600 19304 263652 19310
rect 263600 19246 263652 19252
rect 263612 16574 263640 19246
rect 263612 16546 264192 16574
rect 262956 15972 263008 15978
rect 262956 15914 263008 15920
rect 264164 480 264192 16546
rect 264440 13258 264468 55830
rect 264428 13252 264480 13258
rect 264428 13194 264480 13200
rect 264980 8968 265032 8974
rect 264980 8910 265032 8916
rect 264992 3913 265020 8910
rect 265636 6186 265664 96999
rect 265728 40730 265756 99346
rect 265820 64258 265848 132495
rect 265898 132016 265954 132025
rect 265898 131951 265954 131960
rect 265912 131170 265940 131951
rect 265900 131164 265952 131170
rect 265900 131106 265952 131112
rect 265898 127256 265954 127265
rect 265898 127191 265954 127200
rect 265912 127090 265940 127191
rect 265900 127084 265952 127090
rect 265900 127026 265952 127032
rect 265898 126032 265954 126041
rect 265898 125967 265954 125976
rect 265912 125662 265940 125967
rect 265900 125656 265952 125662
rect 265900 125598 265952 125604
rect 265898 124264 265954 124273
rect 265898 124199 265900 124208
rect 265952 124199 265954 124208
rect 265900 124170 265952 124176
rect 265990 123856 266046 123865
rect 265990 123791 266046 123800
rect 265898 123448 265954 123457
rect 265898 123383 265954 123392
rect 265912 123146 265940 123383
rect 265900 123140 265952 123146
rect 265900 123082 265952 123088
rect 265898 123040 265954 123049
rect 265898 122975 265954 122984
rect 265912 122942 265940 122975
rect 265900 122936 265952 122942
rect 265900 122878 265952 122884
rect 266004 122874 266032 123791
rect 265992 122868 266044 122874
rect 265992 122810 266044 122816
rect 265990 122088 266046 122097
rect 265990 122023 266046 122032
rect 265898 121680 265954 121689
rect 265898 121615 265954 121624
rect 265912 121514 265940 121615
rect 266004 121582 266032 122023
rect 265992 121576 266044 121582
rect 265992 121518 266044 121524
rect 265900 121508 265952 121514
rect 265900 121450 265952 121456
rect 266096 118694 266124 136983
rect 265912 118666 266124 118694
rect 265912 89010 265940 118666
rect 265990 118280 266046 118289
rect 265990 118215 266046 118224
rect 266004 117502 266032 118215
rect 265992 117496 266044 117502
rect 265992 117438 266044 117444
rect 266082 116920 266138 116929
rect 266082 116855 266138 116864
rect 265990 116512 266046 116521
rect 265990 116447 266046 116456
rect 266004 116074 266032 116447
rect 266096 116142 266124 116855
rect 266084 116136 266136 116142
rect 266084 116078 266136 116084
rect 265992 116068 266044 116074
rect 265992 116010 266044 116016
rect 265990 114880 266046 114889
rect 265990 114815 266046 114824
rect 266004 114714 266032 114815
rect 265992 114708 266044 114714
rect 265992 114650 266044 114656
rect 265990 111344 266046 111353
rect 265990 111279 266046 111288
rect 266004 110634 266032 111279
rect 265992 110628 266044 110634
rect 265992 110570 266044 110576
rect 265990 108352 266046 108361
rect 265990 108287 266046 108296
rect 266004 107846 266032 108287
rect 265992 107840 266044 107846
rect 265992 107782 266044 107788
rect 265992 104984 266044 104990
rect 265990 104952 265992 104961
rect 266044 104952 266046 104961
rect 265990 104887 266046 104896
rect 265990 104136 266046 104145
rect 265990 104071 266046 104080
rect 266004 103766 266032 104071
rect 265992 103760 266044 103766
rect 265992 103702 266044 103708
rect 266082 103184 266138 103193
rect 266082 103119 266138 103128
rect 266096 102338 266124 103119
rect 266084 102332 266136 102338
rect 266084 102274 266136 102280
rect 265990 99784 266046 99793
rect 265990 99719 266046 99728
rect 266004 99414 266032 99719
rect 265992 99408 266044 99414
rect 265992 99350 266044 99356
rect 266082 98832 266138 98841
rect 266082 98767 266138 98776
rect 266096 98190 266124 98767
rect 266084 98184 266136 98190
rect 266084 98126 266136 98132
rect 265900 89004 265952 89010
rect 265900 88946 265952 88952
rect 265808 64252 265860 64258
rect 265808 64194 265860 64200
rect 265716 40724 265768 40730
rect 265716 40666 265768 40672
rect 266360 36576 266412 36582
rect 266360 36518 266412 36524
rect 266372 16574 266400 36518
rect 266372 16546 266584 16574
rect 265624 6180 265676 6186
rect 265624 6122 265676 6128
rect 264978 3904 265034 3913
rect 264978 3839 265034 3848
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 3839
rect 266556 480 266584 16546
rect 267016 3534 267044 320894
rect 267096 318096 267148 318102
rect 267096 318038 267148 318044
rect 267108 61402 267136 318038
rect 268396 177478 268424 324974
rect 269776 182918 269804 335990
rect 269856 327820 269908 327826
rect 269856 327762 269908 327768
rect 269764 182912 269816 182918
rect 269764 182854 269816 182860
rect 269868 181830 269896 327762
rect 271144 311160 271196 311166
rect 271144 311102 271196 311108
rect 269948 298240 270000 298246
rect 269948 298182 270000 298188
rect 269856 181824 269908 181830
rect 269856 181766 269908 181772
rect 269960 178673 269988 298182
rect 271156 184346 271184 311102
rect 276664 302252 276716 302258
rect 276664 302194 276716 302200
rect 273904 292664 273956 292670
rect 273904 292606 273956 292612
rect 272524 282940 272576 282946
rect 272524 282882 272576 282888
rect 271236 251932 271288 251938
rect 271236 251874 271288 251880
rect 271144 184340 271196 184346
rect 271144 184282 271196 184288
rect 271248 178770 271276 251874
rect 272536 180470 272564 282882
rect 272616 201000 272668 201006
rect 272616 200942 272668 200948
rect 272524 180464 272576 180470
rect 272524 180406 272576 180412
rect 272628 178974 272656 200942
rect 273916 180402 273944 292606
rect 273996 291440 274048 291446
rect 273996 291382 274048 291388
rect 273904 180396 273956 180402
rect 273904 180338 273956 180344
rect 274008 180334 274036 291382
rect 275284 217388 275336 217394
rect 275284 217330 275336 217336
rect 274088 187060 274140 187066
rect 274088 187002 274140 187008
rect 273996 180328 274048 180334
rect 273996 180270 274048 180276
rect 272616 178968 272668 178974
rect 272616 178910 272668 178916
rect 271236 178764 271288 178770
rect 271236 178706 271288 178712
rect 269946 178664 270002 178673
rect 269946 178599 270002 178608
rect 268384 177472 268436 177478
rect 268384 177414 268436 177420
rect 274100 176186 274128 187002
rect 275296 177614 275324 217330
rect 275284 177608 275336 177614
rect 275284 177550 275336 177556
rect 276676 177449 276704 302194
rect 279424 299600 279476 299606
rect 279424 299542 279476 299548
rect 278044 298172 278096 298178
rect 278044 298114 278096 298120
rect 276756 236768 276808 236774
rect 276756 236710 276808 236716
rect 276768 179042 276796 236710
rect 276848 229764 276900 229770
rect 276848 229706 276900 229712
rect 276756 179036 276808 179042
rect 276756 178978 276808 178984
rect 276662 177440 276718 177449
rect 276662 177375 276718 177384
rect 274088 176180 274140 176186
rect 274088 176122 274140 176128
rect 276860 175982 276888 229706
rect 278056 177682 278084 298114
rect 278136 277500 278188 277506
rect 278136 277442 278188 277448
rect 278148 188630 278176 277442
rect 278228 202156 278280 202162
rect 278228 202098 278280 202104
rect 278136 188624 278188 188630
rect 278136 188566 278188 188572
rect 278044 177676 278096 177682
rect 278044 177618 278096 177624
rect 278240 176118 278268 202098
rect 278320 193996 278372 194002
rect 278320 193938 278372 193944
rect 278228 176112 278280 176118
rect 278228 176054 278280 176060
rect 276848 175976 276900 175982
rect 276848 175918 276900 175924
rect 278332 175817 278360 193938
rect 279436 180794 279464 299542
rect 280896 277432 280948 277438
rect 280896 277374 280948 277380
rect 280804 258120 280856 258126
rect 280804 258062 280856 258068
rect 279516 243024 279568 243030
rect 279516 242966 279568 242972
rect 279528 188698 279556 242966
rect 279516 188692 279568 188698
rect 279516 188634 279568 188640
rect 280344 188556 280396 188562
rect 280344 188498 280396 188504
rect 280160 188420 280212 188426
rect 280160 188362 280212 188368
rect 279436 180766 279648 180794
rect 279424 177404 279476 177410
rect 279424 177346 279476 177352
rect 278318 175808 278374 175817
rect 278318 175743 278374 175752
rect 279330 175808 279386 175817
rect 279330 175743 279386 175752
rect 279344 174457 279372 175743
rect 279436 175273 279464 177346
rect 279516 176656 279568 176662
rect 279516 176598 279568 176604
rect 279528 175817 279556 176598
rect 279620 176050 279648 180766
rect 279608 176044 279660 176050
rect 279608 175986 279660 175992
rect 279514 175808 279570 175817
rect 279514 175743 279570 175752
rect 279422 175264 279478 175273
rect 279422 175199 279478 175208
rect 279330 174448 279386 174457
rect 279330 174383 279386 174392
rect 280172 136377 280200 188362
rect 280252 185836 280304 185842
rect 280252 185778 280304 185784
rect 280264 147801 280292 185778
rect 280356 156369 280384 188498
rect 280816 166326 280844 258062
rect 280908 198150 280936 277374
rect 282196 273970 282224 363598
rect 283012 301096 283064 301102
rect 283012 301038 283064 301044
rect 282918 298208 282974 298217
rect 282918 298143 282974 298152
rect 282276 287768 282328 287774
rect 282276 287710 282328 287716
rect 282184 273964 282236 273970
rect 282184 273906 282236 273912
rect 281724 232620 281776 232626
rect 281724 232562 281776 232568
rect 280896 198144 280948 198150
rect 280896 198086 280948 198092
rect 281630 196616 281686 196625
rect 281630 196551 281686 196560
rect 281540 176180 281592 176186
rect 281540 176122 281592 176128
rect 281552 172417 281580 176122
rect 281538 172408 281594 172417
rect 281538 172343 281594 172352
rect 281644 168609 281672 196551
rect 281630 168600 281686 168609
rect 281630 168535 281686 168544
rect 280804 166320 280856 166326
rect 280804 166262 280856 166268
rect 281632 166320 281684 166326
rect 281632 166262 281684 166268
rect 280342 156360 280398 156369
rect 280342 156295 280398 156304
rect 281540 155984 281592 155990
rect 281540 155926 281592 155932
rect 281552 152425 281580 155926
rect 281538 152416 281594 152425
rect 281538 152351 281594 152360
rect 280250 147792 280306 147801
rect 280250 147727 280306 147736
rect 280158 136368 280214 136377
rect 280158 136303 280214 136312
rect 281644 130937 281672 166262
rect 281630 130928 281686 130937
rect 281630 130863 281686 130872
rect 281630 130112 281686 130121
rect 281630 130047 281686 130056
rect 281644 129878 281672 130047
rect 281632 129872 281684 129878
rect 281632 129814 281684 129820
rect 281632 128308 281684 128314
rect 281632 128250 281684 128256
rect 281644 127809 281672 128250
rect 281630 127800 281686 127809
rect 281630 127735 281686 127744
rect 267278 125080 267334 125089
rect 267278 125015 267334 125024
rect 267188 106276 267240 106282
rect 267188 106218 267240 106224
rect 267096 61396 267148 61402
rect 267096 61338 267148 61344
rect 267200 58682 267228 106218
rect 267292 94518 267320 125015
rect 281632 121372 281684 121378
rect 281632 121314 281684 121320
rect 281644 120193 281672 121314
rect 281630 120184 281686 120193
rect 281630 120119 281686 120128
rect 281630 114064 281686 114073
rect 281630 113999 281686 114008
rect 280250 113248 280306 113257
rect 280250 113183 280306 113192
rect 280158 108624 280214 108633
rect 280158 108559 280214 108568
rect 279330 96656 279386 96665
rect 279330 96591 279386 96600
rect 267280 94512 267332 94518
rect 267280 94454 267332 94460
rect 270972 93838 271000 96016
rect 270960 93832 271012 93838
rect 270960 93774 271012 93780
rect 270972 93498 271000 93774
rect 276952 93702 276980 96016
rect 279344 95169 279372 96591
rect 279330 95160 279386 95169
rect 280172 95130 280200 108559
rect 279330 95095 279386 95104
rect 280160 95124 280212 95130
rect 280160 95066 280212 95072
rect 280264 95062 280292 113183
rect 281540 107908 281592 107914
rect 281540 107850 281592 107856
rect 281552 107817 281580 107850
rect 281538 107808 281594 107817
rect 281538 107743 281594 107752
rect 280342 104816 280398 104825
rect 280342 104751 280398 104760
rect 280252 95056 280304 95062
rect 280252 94998 280304 95004
rect 276940 93696 276992 93702
rect 276940 93638 276992 93644
rect 270960 93492 271012 93498
rect 270960 93434 271012 93440
rect 280356 92274 280384 104751
rect 281538 102504 281594 102513
rect 281538 102439 281594 102448
rect 280436 101448 280488 101454
rect 280436 101390 280488 101396
rect 280344 92268 280396 92274
rect 280344 92210 280396 92216
rect 276020 86284 276072 86290
rect 276020 86226 276072 86232
rect 273260 80708 273312 80714
rect 273260 80650 273312 80656
rect 269120 75200 269172 75206
rect 269120 75142 269172 75148
rect 267188 58676 267240 58682
rect 267188 58618 267240 58624
rect 268384 57248 268436 57254
rect 268384 57190 268436 57196
rect 268396 20670 268424 57190
rect 267740 20664 267792 20670
rect 267740 20606 267792 20612
rect 268384 20664 268436 20670
rect 268384 20606 268436 20612
rect 267752 16574 267780 20606
rect 269132 16574 269160 75142
rect 271880 58676 271932 58682
rect 271880 58618 271932 58624
rect 269764 44872 269816 44878
rect 269764 44814 269816 44820
rect 267752 16546 268424 16574
rect 269132 16546 269712 16574
rect 267004 3528 267056 3534
rect 267004 3470 267056 3476
rect 267740 3324 267792 3330
rect 267740 3266 267792 3272
rect 267752 480 267780 3266
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 269684 3482 269712 16546
rect 269776 4146 269804 44814
rect 270500 21412 270552 21418
rect 270500 21354 270552 21360
rect 270512 16574 270540 21354
rect 271892 16574 271920 58618
rect 270512 16546 270816 16574
rect 271892 16546 272472 16574
rect 269764 4140 269816 4146
rect 269764 4082 269816 4088
rect 269684 3454 270080 3482
rect 270052 480 270080 3454
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272444 480 272472 16546
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 80650
rect 273352 19984 273404 19990
rect 273352 19926 273404 19932
rect 273364 19242 273392 19926
rect 273352 19236 273404 19242
rect 273352 19178 273404 19184
rect 273364 3330 273392 19178
rect 276032 3602 276060 86226
rect 278044 77988 278096 77994
rect 278044 77930 278096 77936
rect 276664 60036 276716 60042
rect 276664 59978 276716 59984
rect 276676 28966 276704 59978
rect 276112 28960 276164 28966
rect 276112 28902 276164 28908
rect 276664 28960 276716 28966
rect 276664 28902 276716 28908
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 274824 3528 274876 3534
rect 276124 3482 276152 28902
rect 278056 9654 278084 77930
rect 280252 61396 280304 61402
rect 280252 61338 280304 61344
rect 278044 9648 278096 9654
rect 278044 9590 278096 9596
rect 278320 9648 278372 9654
rect 278320 9590 278372 9596
rect 276756 3596 276808 3602
rect 276756 3538 276808 3544
rect 274824 3470 274876 3476
rect 273352 3324 273404 3330
rect 273352 3266 273404 3272
rect 274836 480 274864 3470
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 3538
rect 278332 480 278360 9590
rect 280264 2990 280292 61338
rect 280448 16574 280476 101390
rect 281552 96422 281580 102439
rect 281540 96416 281592 96422
rect 281540 96358 281592 96364
rect 281644 92410 281672 113999
rect 281736 100881 281764 232562
rect 282288 221610 282316 287710
rect 282276 221604 282328 221610
rect 282276 221546 282328 221552
rect 282736 171080 282788 171086
rect 282736 171022 282788 171028
rect 282748 170105 282776 171022
rect 282828 171012 282880 171018
rect 282828 170954 282880 170960
rect 282840 170921 282868 170954
rect 282826 170912 282882 170921
rect 282826 170847 282882 170856
rect 282734 170096 282790 170105
rect 282734 170031 282790 170040
rect 281906 169416 281962 169425
rect 281906 169351 281962 169360
rect 281920 168910 281948 169351
rect 281908 168904 281960 168910
rect 281908 168846 281960 168852
rect 281908 168360 281960 168366
rect 281908 168302 281960 168308
rect 281920 167793 281948 168302
rect 282368 168292 282420 168298
rect 282368 168234 282420 168240
rect 281906 167784 281962 167793
rect 281906 167719 281962 167728
rect 282380 167113 282408 168234
rect 282366 167104 282422 167113
rect 282366 167039 282422 167048
rect 282092 167000 282144 167006
rect 282092 166942 282144 166948
rect 282104 166297 282132 166942
rect 282090 166288 282146 166297
rect 282090 166223 282146 166232
rect 282092 165572 282144 165578
rect 282092 165514 282144 165520
rect 282104 164801 282132 165514
rect 282366 165472 282422 165481
rect 282366 165407 282422 165416
rect 282090 164792 282146 164801
rect 282090 164727 282146 164736
rect 282380 164286 282408 165407
rect 282368 164280 282420 164286
rect 282368 164222 282420 164228
rect 282184 164212 282236 164218
rect 282184 164154 282236 164160
rect 282196 163169 282224 164154
rect 282828 164144 282880 164150
rect 282828 164086 282880 164092
rect 282840 163985 282868 164086
rect 282826 163976 282882 163985
rect 282826 163911 282882 163920
rect 282182 163160 282238 163169
rect 282182 163095 282238 163104
rect 282092 162852 282144 162858
rect 282092 162794 282144 162800
rect 282104 162489 282132 162794
rect 282828 162784 282880 162790
rect 282828 162726 282880 162732
rect 282090 162480 282146 162489
rect 282090 162415 282146 162424
rect 282840 161673 282868 162726
rect 282826 161664 282882 161673
rect 282826 161599 282882 161608
rect 282736 161424 282788 161430
rect 282736 161366 282788 161372
rect 282748 160177 282776 161366
rect 282826 160848 282882 160857
rect 282826 160783 282882 160792
rect 282840 160478 282868 160783
rect 282828 160472 282880 160478
rect 282828 160414 282880 160420
rect 282734 160168 282790 160177
rect 282734 160103 282790 160112
rect 282092 160064 282144 160070
rect 282092 160006 282144 160012
rect 282104 159361 282132 160006
rect 282090 159352 282146 159361
rect 282090 159287 282146 159296
rect 282736 158704 282788 158710
rect 282736 158646 282788 158652
rect 282748 157865 282776 158646
rect 282828 158636 282880 158642
rect 282828 158578 282880 158584
rect 282840 158545 282868 158578
rect 282826 158536 282882 158545
rect 282826 158471 282882 158480
rect 282734 157856 282790 157865
rect 282734 157791 282790 157800
rect 282092 157344 282144 157350
rect 282092 157286 282144 157292
rect 282104 157049 282132 157286
rect 282090 157040 282146 157049
rect 282090 156975 282146 156984
rect 282368 155916 282420 155922
rect 282368 155858 282420 155864
rect 282092 155848 282144 155854
rect 282092 155790 282144 155796
rect 282104 155553 282132 155790
rect 282090 155544 282146 155553
rect 282090 155479 282146 155488
rect 282380 154737 282408 155858
rect 282366 154728 282422 154737
rect 282366 154663 282422 154672
rect 282460 154556 282512 154562
rect 282460 154498 282512 154504
rect 281908 154216 281960 154222
rect 281908 154158 281960 154164
rect 281920 154057 281948 154158
rect 281906 154048 281962 154057
rect 281906 153983 281962 153992
rect 282472 153241 282500 154498
rect 282458 153232 282514 153241
rect 282458 153167 282514 153176
rect 281908 151768 281960 151774
rect 281906 151736 281908 151745
rect 281960 151736 281962 151745
rect 281906 151671 281962 151680
rect 282276 151156 282328 151162
rect 282276 151098 282328 151104
rect 282288 150929 282316 151098
rect 282274 150920 282330 150929
rect 282274 150855 282330 150864
rect 282736 150408 282788 150414
rect 282736 150350 282788 150356
rect 282748 149433 282776 150350
rect 282828 150340 282880 150346
rect 282828 150282 282880 150288
rect 282840 150113 282868 150282
rect 282826 150104 282882 150113
rect 282826 150039 282882 150048
rect 282734 149424 282790 149433
rect 282734 149359 282790 149368
rect 282828 149048 282880 149054
rect 282828 148990 282880 148996
rect 282840 148617 282868 148990
rect 282826 148608 282882 148617
rect 282826 148543 282882 148552
rect 282828 147620 282880 147626
rect 282828 147562 282880 147568
rect 282840 147121 282868 147562
rect 282826 147112 282882 147121
rect 282826 147047 282882 147056
rect 282826 146296 282882 146305
rect 282826 146231 282828 146240
rect 282880 146231 282882 146240
rect 282828 146202 282880 146208
rect 282736 146192 282788 146198
rect 282736 146134 282788 146140
rect 282748 145489 282776 146134
rect 282734 145480 282790 145489
rect 282734 145415 282790 145424
rect 282736 144900 282788 144906
rect 282736 144842 282788 144848
rect 282748 143993 282776 144842
rect 282828 144832 282880 144838
rect 282826 144800 282828 144809
rect 282880 144800 282882 144809
rect 282826 144735 282882 144744
rect 282734 143984 282790 143993
rect 282734 143919 282790 143928
rect 282092 143540 282144 143546
rect 282092 143482 282144 143488
rect 282104 143177 282132 143482
rect 282090 143168 282146 143177
rect 282090 143103 282146 143112
rect 282828 142520 282880 142526
rect 282826 142488 282828 142497
rect 282880 142488 282882 142497
rect 282826 142423 282882 142432
rect 282736 142112 282788 142118
rect 282736 142054 282788 142060
rect 282748 140865 282776 142054
rect 282826 141672 282882 141681
rect 282826 141607 282882 141616
rect 282840 141370 282868 141607
rect 282828 141364 282880 141370
rect 282828 141306 282880 141312
rect 282734 140856 282790 140865
rect 282734 140791 282790 140800
rect 282828 140752 282880 140758
rect 282828 140694 282880 140700
rect 282840 140185 282868 140694
rect 282826 140176 282882 140185
rect 282826 140111 282882 140120
rect 282736 139392 282788 139398
rect 282736 139334 282788 139340
rect 282826 139360 282882 139369
rect 282748 138553 282776 139334
rect 282826 139295 282828 139304
rect 282880 139295 282882 139304
rect 282828 139266 282880 139272
rect 282734 138544 282790 138553
rect 282734 138479 282790 138488
rect 282828 137964 282880 137970
rect 282828 137906 282880 137912
rect 282840 137873 282868 137906
rect 282826 137864 282882 137873
rect 282276 137828 282328 137834
rect 282826 137799 282882 137808
rect 282276 137770 282328 137776
rect 282288 137057 282316 137770
rect 282274 137048 282330 137057
rect 282274 136983 282330 136992
rect 282368 136604 282420 136610
rect 282368 136546 282420 136552
rect 282380 135561 282408 136546
rect 282366 135552 282422 135561
rect 282366 135487 282422 135496
rect 282736 135244 282788 135250
rect 282736 135186 282788 135192
rect 282748 134065 282776 135186
rect 282828 135176 282880 135182
rect 282828 135118 282880 135124
rect 282840 134745 282868 135118
rect 282826 134736 282882 134745
rect 282826 134671 282882 134680
rect 282734 134056 282790 134065
rect 282734 133991 282790 134000
rect 282000 133884 282052 133890
rect 282000 133826 282052 133832
rect 282012 133249 282040 133826
rect 282184 133476 282236 133482
rect 282184 133418 282236 133424
rect 281998 133240 282054 133249
rect 281998 133175 282054 133184
rect 282196 123185 282224 133418
rect 282828 132456 282880 132462
rect 282274 132424 282330 132433
rect 282828 132398 282880 132404
rect 282274 132359 282330 132368
rect 282288 131374 282316 132359
rect 282840 131753 282868 132398
rect 282826 131744 282882 131753
rect 282826 131679 282882 131688
rect 282276 131368 282328 131374
rect 282276 131310 282328 131316
rect 282828 129736 282880 129742
rect 282828 129678 282880 129684
rect 282840 128625 282868 129678
rect 282826 128616 282882 128625
rect 282826 128551 282882 128560
rect 282276 127492 282328 127498
rect 282276 127434 282328 127440
rect 282288 127129 282316 127434
rect 282274 127120 282330 127129
rect 282274 127055 282330 127064
rect 282828 126948 282880 126954
rect 282828 126890 282880 126896
rect 282840 126313 282868 126890
rect 282826 126304 282882 126313
rect 282826 126239 282882 126248
rect 282828 125588 282880 125594
rect 282828 125530 282880 125536
rect 282840 125497 282868 125530
rect 282826 125488 282882 125497
rect 282826 125423 282882 125432
rect 282182 123176 282238 123185
rect 282182 123111 282238 123120
rect 282828 122732 282880 122738
rect 282828 122674 282880 122680
rect 282840 121689 282868 122674
rect 282826 121680 282882 121689
rect 282826 121615 282882 121624
rect 281908 121440 281960 121446
rect 281908 121382 281960 121388
rect 281920 120873 281948 121382
rect 281906 120864 281962 120873
rect 281906 120799 281962 120808
rect 282092 120080 282144 120086
rect 282092 120022 282144 120028
rect 282104 119377 282132 120022
rect 282090 119368 282146 119377
rect 282090 119303 282146 119312
rect 282460 118652 282512 118658
rect 282460 118594 282512 118600
rect 282472 117881 282500 118594
rect 282826 118552 282882 118561
rect 282826 118487 282882 118496
rect 282840 118046 282868 118487
rect 282828 118040 282880 118046
rect 282828 117982 282880 117988
rect 282458 117872 282514 117881
rect 282458 117807 282514 117816
rect 282552 117292 282604 117298
rect 282552 117234 282604 117240
rect 282564 116385 282592 117234
rect 282550 116376 282606 116385
rect 282550 116311 282606 116320
rect 282552 115932 282604 115938
rect 282552 115874 282604 115880
rect 282564 114753 282592 115874
rect 282828 115864 282880 115870
rect 282828 115806 282880 115812
rect 282840 115569 282868 115806
rect 282826 115560 282882 115569
rect 282826 115495 282882 115504
rect 282550 114744 282606 114753
rect 282550 114679 282606 114688
rect 282092 113144 282144 113150
rect 282092 113086 282144 113092
rect 282104 112441 282132 113086
rect 282090 112432 282146 112441
rect 282090 112367 282146 112376
rect 282828 111784 282880 111790
rect 282828 111726 282880 111732
rect 282840 110945 282868 111726
rect 282826 110936 282882 110945
rect 282826 110871 282882 110880
rect 282276 110424 282328 110430
rect 282276 110366 282328 110372
rect 282288 109449 282316 110366
rect 282274 109440 282330 109449
rect 282274 109375 282330 109384
rect 282826 107128 282882 107137
rect 282932 107114 282960 298143
rect 283024 122505 283052 301038
rect 287336 286340 287388 286346
rect 287336 286282 287388 286288
rect 287152 264988 287204 264994
rect 287152 264930 287204 264936
rect 284300 262336 284352 262342
rect 284300 262278 284352 262284
rect 283104 252612 283156 252618
rect 283104 252554 283156 252560
rect 283116 155990 283144 252554
rect 283196 203720 283248 203726
rect 283196 203662 283248 203668
rect 283104 155984 283156 155990
rect 283104 155926 283156 155932
rect 283010 122496 283066 122505
rect 283010 122431 283066 122440
rect 283208 107914 283236 203662
rect 284312 133482 284340 262278
rect 284392 233912 284444 233918
rect 284392 233854 284444 233860
rect 284404 151774 284432 233854
rect 285680 206304 285732 206310
rect 285680 206246 285732 206252
rect 284484 184408 284536 184414
rect 284484 184350 284536 184356
rect 284392 151768 284444 151774
rect 284392 151710 284444 151716
rect 284300 133476 284352 133482
rect 284300 133418 284352 133424
rect 283196 107908 283248 107914
rect 283196 107850 283248 107856
rect 282882 107086 282960 107114
rect 282826 107063 282882 107072
rect 284496 104854 284524 184350
rect 285692 137834 285720 206246
rect 285956 191140 286008 191146
rect 285956 191082 286008 191088
rect 285864 189848 285916 189854
rect 285864 189790 285916 189796
rect 285772 184272 285824 184278
rect 285772 184214 285824 184220
rect 285680 137828 285732 137834
rect 285680 137770 285732 137776
rect 285784 127498 285812 184214
rect 285876 151162 285904 189790
rect 285968 154222 285996 191082
rect 287060 176112 287112 176118
rect 287060 176054 287112 176060
rect 287072 168910 287100 176054
rect 287060 168904 287112 168910
rect 287060 168846 287112 168852
rect 285956 154216 286008 154222
rect 285956 154158 286008 154164
rect 285864 151156 285916 151162
rect 285864 151098 285916 151104
rect 287164 141370 287192 264930
rect 287244 178968 287296 178974
rect 287244 178910 287296 178916
rect 287152 141364 287204 141370
rect 287152 141306 287204 141312
rect 287060 127628 287112 127634
rect 287060 127570 287112 127576
rect 285772 127492 285824 127498
rect 285772 127434 285824 127440
rect 282000 104848 282052 104854
rect 282000 104790 282052 104796
rect 284484 104848 284536 104854
rect 284484 104790 284536 104796
rect 282012 104009 282040 104790
rect 281998 104000 282054 104009
rect 281998 103935 282054 103944
rect 282828 102128 282880 102134
rect 282828 102070 282880 102076
rect 282840 101697 282868 102070
rect 282826 101688 282882 101697
rect 282826 101623 282882 101632
rect 281722 100872 281778 100881
rect 281722 100807 281778 100816
rect 281722 100192 281778 100201
rect 281722 100127 281778 100136
rect 281632 92404 281684 92410
rect 281632 92346 281684 92352
rect 281736 92342 281764 100127
rect 284300 100020 284352 100026
rect 284300 99962 284352 99968
rect 281906 97880 281962 97889
rect 281906 97815 281962 97824
rect 281920 93770 281948 97815
rect 281908 93764 281960 93770
rect 281908 93706 281960 93712
rect 281724 92336 281776 92342
rect 281724 92278 281776 92284
rect 283564 29844 283616 29850
rect 283564 29786 283616 29792
rect 280448 16546 280752 16574
rect 279516 2984 279568 2990
rect 279516 2926 279568 2932
rect 280252 2984 280304 2990
rect 280252 2926 280304 2932
rect 279528 480 279556 2926
rect 280724 480 280752 16546
rect 283576 12442 283604 29786
rect 283104 12436 283156 12442
rect 283104 12378 283156 12384
rect 283564 12436 283616 12442
rect 283564 12378 283616 12384
rect 281908 11756 281960 11762
rect 281908 11698 281960 11704
rect 281920 6866 281948 11698
rect 281908 6860 281960 6866
rect 281908 6802 281960 6808
rect 281920 480 281948 6802
rect 283116 480 283144 12378
rect 284312 480 284340 99962
rect 286324 62824 286376 62830
rect 286324 62766 286376 62772
rect 286336 16574 286364 62766
rect 287072 16574 287100 127570
rect 287256 118046 287284 178910
rect 287348 142526 287376 286282
rect 288532 238196 288584 238202
rect 288532 238138 288584 238144
rect 288440 205012 288492 205018
rect 288440 204954 288492 204960
rect 287336 142520 287388 142526
rect 287336 142462 287388 142468
rect 288452 129878 288480 204954
rect 288544 164286 288572 238138
rect 290096 235272 290148 235278
rect 290096 235214 290148 235220
rect 289912 185904 289964 185910
rect 289912 185846 289964 185852
rect 288624 180464 288676 180470
rect 288624 180406 288676 180412
rect 288532 164280 288584 164286
rect 288532 164222 288584 164228
rect 288636 131374 288664 180406
rect 288716 177676 288768 177682
rect 288716 177618 288768 177624
rect 288728 160478 288756 177618
rect 289820 176044 289872 176050
rect 289820 175986 289872 175992
rect 289832 171018 289860 175986
rect 289820 171012 289872 171018
rect 289820 170954 289872 170960
rect 288716 160472 288768 160478
rect 288716 160414 288768 160420
rect 289924 147626 289952 185846
rect 290004 179036 290056 179042
rect 290004 178978 290056 178984
rect 290016 168298 290044 178978
rect 290004 168292 290056 168298
rect 290004 168234 290056 168240
rect 289912 147620 289964 147626
rect 289912 147562 289964 147568
rect 288624 131368 288676 131374
rect 288624 131310 288676 131316
rect 288440 129872 288492 129878
rect 288440 129814 288492 129820
rect 287244 118040 287296 118046
rect 287244 117982 287296 117988
rect 290108 102134 290136 235214
rect 291292 186992 291344 186998
rect 291292 186934 291344 186940
rect 291200 184204 291252 184210
rect 291200 184146 291252 184152
rect 291212 146198 291240 184146
rect 291304 171086 291332 186934
rect 291384 175976 291436 175982
rect 291384 175918 291436 175924
rect 291292 171080 291344 171086
rect 291292 171022 291344 171028
rect 291396 164150 291424 175918
rect 291384 164144 291436 164150
rect 291384 164086 291436 164092
rect 291200 146192 291252 146198
rect 291200 146134 291252 146140
rect 290096 102128 290148 102134
rect 290096 102070 290148 102076
rect 291856 89078 291884 397462
rect 298744 392012 298796 392018
rect 298744 391954 298796 391960
rect 297364 354000 297416 354006
rect 297364 353942 297416 353948
rect 295984 329112 296036 329118
rect 295984 329054 296036 329060
rect 293222 307048 293278 307057
rect 293222 306983 293278 306992
rect 292672 191344 292724 191350
rect 292672 191286 292724 191292
rect 292580 177540 292632 177546
rect 292580 177482 292632 177488
rect 292592 125594 292620 177482
rect 292684 165578 292712 191286
rect 292764 188692 292816 188698
rect 292764 188634 292816 188640
rect 292672 165572 292724 165578
rect 292672 165514 292724 165520
rect 292776 162790 292804 188634
rect 292764 162784 292816 162790
rect 292764 162726 292816 162732
rect 292580 125588 292632 125594
rect 292580 125530 292632 125536
rect 291844 89072 291896 89078
rect 291844 89014 291896 89020
rect 291200 83564 291252 83570
rect 291200 83506 291252 83512
rect 288440 29640 288492 29646
rect 288440 29582 288492 29588
rect 287704 28280 287756 28286
rect 287704 28222 287756 28228
rect 286336 16546 286640 16574
rect 287072 16546 287376 16574
rect 286612 4049 286640 16546
rect 286598 4040 286654 4049
rect 286598 3975 286654 3984
rect 285404 3460 285456 3466
rect 285404 3402 285456 3408
rect 285416 480 285444 3402
rect 286612 480 286640 3975
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 287716 3466 287744 28222
rect 288452 16574 288480 29582
rect 289084 25560 289136 25566
rect 289084 25502 289136 25508
rect 288452 16546 289032 16574
rect 287704 3460 287756 3466
rect 287704 3402 287756 3408
rect 289004 480 289032 16546
rect 289096 3534 289124 25502
rect 291212 16574 291240 83506
rect 291212 16546 291424 16574
rect 289084 3528 289136 3534
rect 289084 3470 289136 3476
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 290200 480 290228 3470
rect 291396 480 291424 16546
rect 293236 13802 293264 306983
rect 293960 284436 294012 284442
rect 293960 284378 294012 284384
rect 293972 161430 294000 284378
rect 295432 196716 295484 196722
rect 295432 196658 295484 196664
rect 294052 195492 294104 195498
rect 294052 195434 294104 195440
rect 293960 161424 294012 161430
rect 293960 161366 294012 161372
rect 294064 110430 294092 195434
rect 294144 180260 294196 180266
rect 294144 180202 294196 180208
rect 294156 120086 294184 180202
rect 295340 178900 295392 178906
rect 295340 178842 295392 178848
rect 294236 177608 294288 177614
rect 294236 177550 294288 177556
rect 294248 150346 294276 177550
rect 294236 150340 294288 150346
rect 294236 150282 294288 150288
rect 294144 120080 294196 120086
rect 294144 120022 294196 120028
rect 295352 113150 295380 178842
rect 295444 168366 295472 196658
rect 295524 185632 295576 185638
rect 295524 185574 295576 185580
rect 295432 168360 295484 168366
rect 295432 168302 295484 168308
rect 295536 167006 295564 185574
rect 295524 167000 295576 167006
rect 295524 166942 295576 166948
rect 295996 135930 296024 329054
rect 296720 202292 296772 202298
rect 296720 202234 296772 202240
rect 295984 135924 296036 135930
rect 295984 135866 296036 135872
rect 295340 113144 295392 113150
rect 295340 113086 295392 113092
rect 296732 111790 296760 202234
rect 296904 183116 296956 183122
rect 296904 183058 296956 183064
rect 296812 181756 296864 181762
rect 296812 181698 296864 181704
rect 296824 142118 296852 181698
rect 296916 149054 296944 183058
rect 296904 149048 296956 149054
rect 296904 148990 296956 148996
rect 296812 142112 296864 142118
rect 296812 142054 296864 142060
rect 296720 111784 296772 111790
rect 296720 111726 296772 111732
rect 294052 110424 294104 110430
rect 294052 110366 294104 110372
rect 293960 102808 294012 102814
rect 293960 102750 294012 102756
rect 293224 13796 293276 13802
rect 293224 13738 293276 13744
rect 292580 3596 292632 3602
rect 292580 3538 292632 3544
rect 292592 480 292620 3538
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 13738
rect 293972 3482 294000 102750
rect 297376 66230 297404 353942
rect 298100 301028 298152 301034
rect 298100 300970 298152 300976
rect 298112 162858 298140 300970
rect 298192 201136 298244 201142
rect 298192 201078 298244 201084
rect 298100 162852 298152 162858
rect 298100 162794 298152 162800
rect 298204 135182 298232 201078
rect 298284 181484 298336 181490
rect 298284 181426 298336 181432
rect 298296 144838 298324 181426
rect 298284 144832 298336 144838
rect 298284 144774 298336 144780
rect 298192 135176 298244 135182
rect 298192 135118 298244 135124
rect 298756 92342 298784 391954
rect 300124 324964 300176 324970
rect 300124 324906 300176 324912
rect 299480 221604 299532 221610
rect 299480 221546 299532 221552
rect 299492 139330 299520 221546
rect 299572 203652 299624 203658
rect 299572 203594 299624 203600
rect 299584 164218 299612 203594
rect 299572 164212 299624 164218
rect 299572 164154 299624 164160
rect 300136 141438 300164 324906
rect 302884 322312 302936 322318
rect 302884 322254 302936 322260
rect 300952 296744 301004 296750
rect 300952 296686 301004 296692
rect 300860 266416 300912 266422
rect 300860 266358 300912 266364
rect 300216 181688 300268 181694
rect 300216 181630 300268 181636
rect 300124 141432 300176 141438
rect 300124 141374 300176 141380
rect 299480 139324 299532 139330
rect 299480 139266 299532 139272
rect 298744 92336 298796 92342
rect 298744 92278 298796 92284
rect 298100 90364 298152 90370
rect 298100 90306 298152 90312
rect 298112 87009 298140 90306
rect 300228 89010 300256 181630
rect 300872 158642 300900 266358
rect 300860 158636 300912 158642
rect 300860 158578 300912 158584
rect 300860 144220 300912 144226
rect 300860 144162 300912 144168
rect 300216 89004 300268 89010
rect 300216 88946 300268 88952
rect 298098 87000 298154 87009
rect 298098 86935 298154 86944
rect 299664 66904 299716 66910
rect 299662 66872 299664 66881
rect 299716 66872 299718 66881
rect 299662 66807 299718 66816
rect 296720 66224 296772 66230
rect 296720 66166 296772 66172
rect 297364 66224 297416 66230
rect 297364 66166 297416 66172
rect 295340 64320 295392 64326
rect 295340 64262 295392 64268
rect 294142 31104 294198 31113
rect 294142 31039 294144 31048
rect 294196 31039 294198 31048
rect 294144 31010 294196 31016
rect 294156 26234 294184 31010
rect 294064 26206 294184 26234
rect 294064 3602 294092 26206
rect 294052 3596 294104 3602
rect 294052 3538 294104 3544
rect 295352 3534 295380 64262
rect 296732 16574 296760 66166
rect 298100 40724 298152 40730
rect 298100 40666 298152 40672
rect 296732 16546 297312 16574
rect 295340 3528 295392 3534
rect 293972 3454 294920 3482
rect 295340 3470 295392 3476
rect 296074 3496 296130 3505
rect 294892 480 294920 3454
rect 296074 3431 296130 3440
rect 296088 480 296116 3431
rect 297284 480 297312 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 40666
rect 300872 16574 300900 144162
rect 300964 135250 300992 296686
rect 301504 221536 301556 221542
rect 301504 221478 301556 221484
rect 301044 198144 301096 198150
rect 301044 198086 301096 198092
rect 300952 135244 301004 135250
rect 300952 135186 301004 135192
rect 301056 126954 301084 198086
rect 301044 126948 301096 126954
rect 301044 126890 301096 126896
rect 301516 109002 301544 221478
rect 302240 209160 302292 209166
rect 302240 209102 302292 209108
rect 302252 117298 302280 209102
rect 302332 198008 302384 198014
rect 302332 197950 302384 197956
rect 302240 117292 302292 117298
rect 302240 117234 302292 117240
rect 302344 115870 302372 197950
rect 302424 180396 302476 180402
rect 302424 180338 302476 180344
rect 302436 158710 302464 180338
rect 302424 158704 302476 158710
rect 302424 158646 302476 158652
rect 302332 115864 302384 115870
rect 302332 115806 302384 115812
rect 301504 108996 301556 109002
rect 301504 108938 301556 108944
rect 302240 87644 302292 87650
rect 302240 87586 302292 87592
rect 300872 16546 301544 16574
rect 300766 3496 300822 3505
rect 300766 3431 300822 3440
rect 299664 3188 299716 3194
rect 299664 3130 299716 3136
rect 299676 480 299704 3130
rect 300780 480 300808 3431
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 302252 3194 302280 87586
rect 302896 47598 302924 322254
rect 303620 299532 303672 299538
rect 303620 299474 303672 299480
rect 303632 121378 303660 299474
rect 303712 225616 303764 225622
rect 303712 225558 303764 225564
rect 303724 122738 303752 225558
rect 303804 180328 303856 180334
rect 303804 180270 303856 180276
rect 303816 157350 303844 180270
rect 303804 157344 303856 157350
rect 303804 157286 303856 157292
rect 303712 122732 303764 122738
rect 303712 122674 303764 122680
rect 303620 121372 303672 121378
rect 303620 121314 303672 121320
rect 304276 85542 304304 401610
rect 322940 395344 322992 395350
rect 322940 395286 322992 395292
rect 313924 388476 313976 388482
rect 313924 388418 313976 388424
rect 309784 333260 309836 333266
rect 309784 333202 309836 333208
rect 306380 300960 306432 300966
rect 306380 300902 306432 300908
rect 305644 284980 305696 284986
rect 305644 284922 305696 284928
rect 305000 260908 305052 260914
rect 305000 260850 305052 260856
rect 305012 137970 305040 260850
rect 305092 198076 305144 198082
rect 305092 198018 305144 198024
rect 305000 137964 305052 137970
rect 305000 137906 305052 137912
rect 305104 118658 305132 198018
rect 305184 188352 305236 188358
rect 305184 188294 305236 188300
rect 305196 139398 305224 188294
rect 305184 139392 305236 139398
rect 305184 139334 305236 139340
rect 305656 126274 305684 284922
rect 306392 136610 306420 300902
rect 308404 273964 308456 273970
rect 308404 273906 308456 273912
rect 307760 210452 307812 210458
rect 307760 210394 307812 210400
rect 306472 195356 306524 195362
rect 306472 195298 306524 195304
rect 306380 136604 306432 136610
rect 306380 136546 306432 136552
rect 305644 126268 305696 126274
rect 305644 126210 305696 126216
rect 305092 118652 305144 118658
rect 305092 118594 305144 118600
rect 306484 115938 306512 195298
rect 306564 188624 306616 188630
rect 306564 188566 306616 188572
rect 306576 155854 306604 188566
rect 307024 168428 307076 168434
rect 307024 168370 307076 168376
rect 306564 155848 306616 155854
rect 306564 155790 306616 155796
rect 306472 115932 306524 115938
rect 306472 115874 306524 115880
rect 304264 85536 304316 85542
rect 304264 85478 304316 85484
rect 305000 85536 305052 85542
rect 305000 85478 305052 85484
rect 305012 84862 305040 85478
rect 305000 84856 305052 84862
rect 305000 84798 305052 84804
rect 302884 47592 302936 47598
rect 302884 47534 302936 47540
rect 302896 16574 302924 47534
rect 302896 16546 303200 16574
rect 302240 3188 302292 3194
rect 302240 3130 302292 3136
rect 303172 480 303200 16546
rect 305012 3534 305040 84798
rect 306746 8256 306802 8265
rect 306746 8191 306802 8200
rect 306760 7614 306788 8191
rect 307036 7682 307064 168370
rect 307772 143546 307800 210394
rect 307944 200864 307996 200870
rect 307944 200806 307996 200812
rect 307852 182844 307904 182850
rect 307852 182786 307904 182792
rect 307760 143540 307812 143546
rect 307760 143482 307812 143488
rect 307864 128314 307892 182786
rect 307956 155922 307984 200806
rect 307944 155916 307996 155922
rect 307944 155858 307996 155864
rect 307852 128308 307904 128314
rect 307852 128250 307904 128256
rect 307024 7676 307076 7682
rect 307024 7618 307076 7624
rect 306748 7608 306800 7614
rect 306748 7550 306800 7556
rect 304356 3528 304408 3534
rect 304356 3470 304408 3476
rect 305000 3528 305052 3534
rect 305000 3470 305052 3476
rect 305550 3496 305606 3505
rect 304368 480 304396 3470
rect 305550 3431 305606 3440
rect 305564 480 305592 3431
rect 306760 480 306788 7550
rect 308416 4146 308444 273906
rect 309140 220176 309192 220182
rect 309140 220118 309192 220124
rect 309152 140758 309180 220118
rect 309232 194064 309284 194070
rect 309232 194006 309284 194012
rect 309140 140752 309192 140758
rect 309140 140694 309192 140700
rect 309244 121446 309272 194006
rect 309324 188488 309376 188494
rect 309324 188430 309376 188436
rect 309336 129742 309364 188430
rect 309796 153882 309824 333202
rect 311900 295384 311952 295390
rect 311900 295326 311952 295332
rect 310520 251252 310572 251258
rect 310520 251194 310572 251200
rect 309784 153876 309836 153882
rect 309784 153818 309836 153824
rect 310532 150414 310560 251194
rect 311164 243568 311216 243574
rect 311164 243510 311216 243516
rect 310612 205148 310664 205154
rect 310612 205090 310664 205096
rect 310520 150408 310572 150414
rect 310520 150350 310572 150356
rect 310624 133890 310652 205090
rect 310704 185700 310756 185706
rect 310704 185642 310756 185648
rect 310716 154562 310744 185642
rect 310704 154556 310756 154562
rect 310704 154498 310756 154504
rect 310612 133884 310664 133890
rect 310612 133826 310664 133832
rect 309784 133204 309836 133210
rect 309784 133146 309836 133152
rect 309324 129736 309376 129742
rect 309324 129678 309376 129684
rect 309232 121440 309284 121446
rect 309232 121382 309284 121388
rect 309232 49088 309284 49094
rect 309230 49056 309232 49065
rect 309284 49056 309286 49065
rect 309230 48991 309286 49000
rect 308404 4140 308456 4146
rect 308404 4082 308456 4088
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 354 308026 480
rect 308416 354 308444 4082
rect 309796 3534 309824 133146
rect 311176 104854 311204 243510
rect 311912 146266 311940 295326
rect 311992 276140 312044 276146
rect 311992 276082 312044 276088
rect 311900 146260 311952 146266
rect 311900 146202 311952 146208
rect 312004 144906 312032 276082
rect 313280 238128 313332 238134
rect 313280 238070 313332 238076
rect 312544 178832 312596 178838
rect 312544 178774 312596 178780
rect 311992 144900 312044 144906
rect 311992 144842 312044 144848
rect 312556 128314 312584 178774
rect 313292 160070 313320 238070
rect 313280 160064 313332 160070
rect 313280 160006 313332 160012
rect 313936 145586 313964 388418
rect 318064 351212 318116 351218
rect 318064 351154 318116 351160
rect 316774 338736 316830 338745
rect 316774 338671 316830 338680
rect 314660 294024 314712 294030
rect 314660 293966 314712 293972
rect 314108 181824 314160 181830
rect 314108 181766 314160 181772
rect 314016 166320 314068 166326
rect 314016 166262 314068 166268
rect 313924 145580 313976 145586
rect 313924 145522 313976 145528
rect 312544 128308 312596 128314
rect 312544 128250 312596 128256
rect 311900 124908 311952 124914
rect 311900 124850 311952 124856
rect 311164 104848 311216 104854
rect 311164 104790 311216 104796
rect 311808 72480 311860 72486
rect 311808 72422 311860 72428
rect 311820 69698 311848 72422
rect 311164 69692 311216 69698
rect 311164 69634 311216 69640
rect 311808 69692 311860 69698
rect 311808 69634 311860 69640
rect 311176 16574 311204 69634
rect 311912 16574 311940 124850
rect 313280 50448 313332 50454
rect 313280 50390 313332 50396
rect 313292 16574 313320 50390
rect 314028 50386 314056 166262
rect 314120 76566 314148 181766
rect 314672 132462 314700 293966
rect 316684 279472 316736 279478
rect 316684 279414 316736 279420
rect 315304 256012 315356 256018
rect 315304 255954 315356 255960
rect 314660 132456 314712 132462
rect 314660 132398 314712 132404
rect 315316 120086 315344 255954
rect 315304 120080 315356 120086
rect 315304 120022 315356 120028
rect 316040 111104 316092 111110
rect 316040 111046 316092 111052
rect 314108 76560 314160 76566
rect 314108 76502 314160 76508
rect 314660 73840 314712 73846
rect 314660 73782 314712 73788
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 311176 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 310242 11792 310298 11801
rect 310242 11727 310298 11736
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309784 3528 309836 3534
rect 309784 3470 309836 3476
rect 309060 480 309088 3470
rect 310256 480 310284 11727
rect 311452 480 311480 16546
rect 307914 326 308444 354
rect 307914 -960 308026 326
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 73782
rect 316052 3482 316080 111046
rect 316696 97986 316724 279414
rect 316788 159390 316816 338671
rect 316868 183048 316920 183054
rect 316868 182990 316920 182996
rect 316776 159384 316828 159390
rect 316776 159326 316828 159332
rect 316684 97980 316736 97986
rect 316684 97922 316736 97928
rect 316880 91050 316908 182990
rect 318076 95266 318104 351154
rect 320824 348424 320876 348430
rect 320824 348366 320876 348372
rect 319444 182980 319496 182986
rect 319444 182922 319496 182928
rect 318156 160744 318208 160750
rect 318156 160686 318208 160692
rect 318064 95260 318116 95266
rect 318064 95202 318116 95208
rect 316868 91044 316920 91050
rect 316868 90986 316920 90992
rect 317420 75880 317472 75886
rect 317420 75822 317472 75828
rect 316132 32496 316184 32502
rect 316132 32438 316184 32444
rect 316144 3602 316172 32438
rect 317432 16574 317460 75822
rect 318168 75206 318196 160686
rect 318800 117972 318852 117978
rect 318800 117914 318852 117920
rect 318156 75200 318208 75206
rect 318156 75142 318208 75148
rect 318812 16574 318840 117914
rect 319456 100706 319484 182922
rect 320836 131782 320864 348366
rect 322204 337408 322256 337414
rect 322204 337350 322256 337356
rect 320916 172576 320968 172582
rect 320916 172518 320968 172524
rect 320824 131776 320876 131782
rect 320824 131718 320876 131724
rect 319444 100700 319496 100706
rect 319444 100642 319496 100648
rect 320180 35284 320232 35290
rect 320180 35226 320232 35232
rect 320192 16574 320220 35226
rect 320928 32434 320956 172518
rect 322216 142866 322244 337350
rect 322296 173936 322348 173942
rect 322296 173878 322348 173884
rect 322204 142860 322256 142866
rect 322204 142802 322256 142808
rect 322204 68332 322256 68338
rect 322204 68274 322256 68280
rect 320916 32428 320968 32434
rect 320916 32370 320968 32376
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 316132 3596 316184 3602
rect 316132 3538 316184 3544
rect 317328 3596 317380 3602
rect 317328 3538 317380 3544
rect 316052 3454 316264 3482
rect 316236 480 316264 3454
rect 317340 480 317368 3538
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322216 4146 322244 68274
rect 322308 35222 322336 173878
rect 322952 75886 322980 395286
rect 334716 389836 334768 389842
rect 334716 389778 334768 389784
rect 327724 386436 327776 386442
rect 327724 386378 327776 386384
rect 324964 385076 325016 385082
rect 324964 385018 325016 385024
rect 323584 295996 323636 296002
rect 323584 295938 323636 295944
rect 323596 149734 323624 295938
rect 323676 181620 323728 181626
rect 323676 181562 323728 181568
rect 323584 149728 323636 149734
rect 323584 149670 323636 149676
rect 323688 126954 323716 181562
rect 324976 158030 325004 385018
rect 326344 303748 326396 303754
rect 326344 303690 326396 303696
rect 325148 177472 325200 177478
rect 325148 177414 325200 177420
rect 325056 171148 325108 171154
rect 325056 171090 325108 171096
rect 324964 158024 325016 158030
rect 324964 157966 325016 157972
rect 323676 126948 323728 126954
rect 323676 126890 323728 126896
rect 323032 116612 323084 116618
rect 323032 116554 323084 116560
rect 322940 75880 322992 75886
rect 322940 75822 322992 75828
rect 322296 35216 322348 35222
rect 322296 35158 322348 35164
rect 322204 4140 322256 4146
rect 322204 4082 322256 4088
rect 322112 3596 322164 3602
rect 322112 3538 322164 3544
rect 322124 480 322152 3538
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323044 354 323072 116554
rect 324320 82136 324372 82142
rect 324320 82078 324372 82084
rect 324332 3534 324360 82078
rect 324412 38004 324464 38010
rect 324412 37946 324464 37952
rect 324320 3528 324372 3534
rect 324320 3470 324372 3476
rect 324424 480 324452 37946
rect 325068 37942 325096 171090
rect 325160 83502 325188 177414
rect 325700 123480 325752 123486
rect 325700 123422 325752 123428
rect 325148 83496 325200 83502
rect 325148 83438 325200 83444
rect 325056 37936 325108 37942
rect 325056 37878 325108 37884
rect 325712 16574 325740 123422
rect 326356 95130 326384 303690
rect 327736 164898 327764 386378
rect 331864 372632 331916 372638
rect 331864 372574 331916 372580
rect 330484 254584 330536 254590
rect 330484 254526 330536 254532
rect 329104 193928 329156 193934
rect 329104 193870 329156 193876
rect 327816 167068 327868 167074
rect 327816 167010 327868 167016
rect 327724 164892 327776 164898
rect 327724 164834 327776 164840
rect 327724 138712 327776 138718
rect 327724 138654 327776 138660
rect 327736 111110 327764 138654
rect 327724 111104 327776 111110
rect 327724 111046 327776 111052
rect 326344 95124 326396 95130
rect 326344 95066 326396 95072
rect 327080 89072 327132 89078
rect 327080 89014 327132 89020
rect 327092 16574 327120 89014
rect 327828 39370 327856 167010
rect 329116 96558 329144 193870
rect 330496 115938 330524 254526
rect 331876 136610 331904 372574
rect 334624 307148 334676 307154
rect 334624 307090 334676 307096
rect 331956 302932 332008 302938
rect 331956 302874 332008 302880
rect 331864 136604 331916 136610
rect 331864 136546 331916 136552
rect 330484 115932 330536 115938
rect 330484 115874 330536 115880
rect 329840 111104 329892 111110
rect 329840 111046 329892 111052
rect 329104 96552 329156 96558
rect 329104 96494 329156 96500
rect 328460 76560 328512 76566
rect 328460 76502 328512 76508
rect 327816 39364 327868 39370
rect 327816 39306 327868 39312
rect 328472 16574 328500 76502
rect 329852 16574 329880 111046
rect 331968 93809 331996 302874
rect 333336 178764 333388 178770
rect 333336 178706 333388 178712
rect 333244 175296 333296 175302
rect 333244 175238 333296 175244
rect 332048 151088 332100 151094
rect 332048 151030 332100 151036
rect 331954 93800 332010 93809
rect 331954 93735 332010 93744
rect 332060 83570 332088 151030
rect 332048 83564 332100 83570
rect 332048 83506 332100 83512
rect 331220 83496 331272 83502
rect 331220 83438 331272 83444
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325620 480 325648 3470
rect 323278 354 323390 480
rect 323044 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330404 480 330432 16546
rect 331232 3602 331260 83438
rect 333256 68921 333284 175238
rect 333348 107642 333376 178706
rect 333336 107636 333388 107642
rect 333336 107578 333388 107584
rect 332598 68912 332654 68921
rect 332598 68847 332654 68856
rect 333242 68912 333298 68921
rect 333242 68847 333298 68856
rect 331220 3596 331272 3602
rect 331220 3538 331272 3544
rect 332612 3534 332640 68847
rect 334636 40050 334664 307090
rect 334728 137290 334756 389778
rect 336016 147014 336044 405719
rect 341524 403028 341576 403034
rect 341524 402970 341576 402976
rect 338118 401704 338174 401713
rect 338118 401639 338174 401648
rect 336096 320884 336148 320890
rect 336096 320826 336148 320832
rect 336108 156126 336136 320826
rect 336278 202192 336334 202201
rect 336278 202127 336334 202136
rect 336188 163532 336240 163538
rect 336188 163474 336240 163480
rect 336096 156120 336148 156126
rect 336096 156062 336148 156068
rect 336004 147008 336056 147014
rect 336004 146950 336056 146956
rect 334716 137284 334768 137290
rect 334716 137226 334768 137232
rect 335360 79620 335412 79626
rect 335360 79562 335412 79568
rect 333980 40044 334032 40050
rect 333980 39986 334032 39992
rect 334624 40044 334676 40050
rect 334624 39986 334676 39992
rect 333992 16574 334020 39986
rect 335372 16574 335400 79562
rect 336200 36582 336228 163474
rect 336292 102134 336320 202127
rect 337476 191412 337528 191418
rect 337476 191354 337528 191360
rect 337384 136604 337436 136610
rect 337384 136546 337436 136552
rect 336280 102128 336332 102134
rect 336280 102070 336332 102076
rect 337396 37262 337424 136546
rect 337488 92410 337516 191354
rect 337476 92404 337528 92410
rect 337476 92346 337528 92352
rect 338132 80034 338160 401639
rect 340144 356720 340196 356726
rect 340144 356662 340196 356668
rect 338764 340196 338816 340202
rect 338764 340138 338816 340144
rect 338212 147008 338264 147014
rect 338212 146950 338264 146956
rect 338120 80028 338172 80034
rect 338120 79970 338172 79976
rect 338132 79626 338160 79970
rect 338120 79620 338172 79626
rect 338120 79562 338172 79568
rect 338120 42220 338172 42226
rect 338120 42162 338172 42168
rect 337384 37256 337436 37262
rect 337384 37198 337436 37204
rect 337396 36922 337424 37198
rect 336740 36916 336792 36922
rect 336740 36858 336792 36864
rect 337384 36916 337436 36922
rect 337384 36858 337436 36864
rect 336188 36576 336240 36582
rect 336188 36518 336240 36524
rect 336752 16574 336780 36858
rect 338132 16574 338160 42162
rect 338224 40730 338252 146950
rect 338302 134464 338358 134473
rect 338302 134399 338358 134408
rect 338316 134065 338344 134399
rect 338302 134056 338358 134065
rect 338302 133991 338358 134000
rect 338316 123486 338344 133991
rect 338776 124166 338804 340138
rect 339500 164892 339552 164898
rect 339500 164834 339552 164840
rect 339512 164286 339540 164834
rect 339500 164280 339552 164286
rect 339500 164222 339552 164228
rect 338764 124160 338816 124166
rect 338764 124102 338816 124108
rect 338304 123480 338356 123486
rect 338304 123422 338356 123428
rect 339512 42158 339540 164222
rect 340156 94994 340184 356662
rect 340880 159384 340932 159390
rect 340880 159326 340932 159332
rect 340144 94988 340196 94994
rect 340144 94930 340196 94936
rect 340892 80714 340920 159326
rect 340972 135924 341024 135930
rect 340972 135866 341024 135872
rect 340984 135318 341012 135866
rect 340972 135312 341024 135318
rect 340972 135254 341024 135260
rect 340984 116618 341012 135254
rect 340972 116612 341024 116618
rect 340972 116554 341024 116560
rect 340880 80708 340932 80714
rect 340880 80650 340932 80656
rect 340144 49020 340196 49026
rect 340144 48962 340196 48968
rect 339500 42152 339552 42158
rect 339500 42094 339552 42100
rect 338212 40724 338264 40730
rect 338212 40666 338264 40672
rect 333992 16546 334664 16574
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 332600 3528 332652 3534
rect 332600 3470 332652 3476
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 332692 3460 332744 3466
rect 332692 3402 332744 3408
rect 331588 3392 331640 3398
rect 331588 3334 331640 3340
rect 331600 480 331628 3334
rect 332704 480 332732 3402
rect 333900 480 333928 3470
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336292 480 336320 16546
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 339500 14544 339552 14550
rect 339500 14486 339552 14492
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 14486
rect 340156 3534 340184 48962
rect 341536 41410 341564 402970
rect 349802 381848 349858 381857
rect 349802 381783 349858 381792
rect 342904 379568 342956 379574
rect 342904 379510 342956 379516
rect 341616 305652 341668 305658
rect 341616 305594 341668 305600
rect 341628 151910 341656 305594
rect 342260 300144 342312 300150
rect 342260 300086 342312 300092
rect 341616 151904 341668 151910
rect 341616 151846 341668 151852
rect 342272 151774 342300 300086
rect 342352 158024 342404 158030
rect 342352 157966 342404 157972
rect 342364 157486 342392 157966
rect 342352 157480 342404 157486
rect 342352 157422 342404 157428
rect 342260 151768 342312 151774
rect 342260 151710 342312 151716
rect 342272 151094 342300 151710
rect 342260 151088 342312 151094
rect 342260 151030 342312 151036
rect 342260 149728 342312 149734
rect 342260 149670 342312 149676
rect 342272 149190 342300 149670
rect 342260 149184 342312 149190
rect 342260 149126 342312 149132
rect 342272 102814 342300 149126
rect 342260 102808 342312 102814
rect 342260 102750 342312 102756
rect 342364 86290 342392 157422
rect 342916 95062 342944 379510
rect 346400 378820 346452 378826
rect 346400 378762 346452 378768
rect 343640 319456 343692 319462
rect 343640 319398 343692 319404
rect 343652 161430 343680 319398
rect 345020 316736 345072 316742
rect 345020 316678 345072 316684
rect 344282 188320 344338 188329
rect 344282 188255 344338 188264
rect 343640 161424 343692 161430
rect 343640 161366 343692 161372
rect 343652 160750 343680 161366
rect 343640 160744 343692 160750
rect 343640 160686 343692 160692
rect 343640 156120 343692 156126
rect 343640 156062 343692 156068
rect 343652 101454 343680 156062
rect 343824 141432 343876 141438
rect 343824 141374 343876 141380
rect 343732 137284 343784 137290
rect 343732 137226 343784 137232
rect 343744 136746 343772 137226
rect 343732 136740 343784 136746
rect 343732 136682 343784 136688
rect 343744 117978 343772 136682
rect 343836 124914 343864 141374
rect 343824 124908 343876 124914
rect 343824 124850 343876 124856
rect 343732 117972 343784 117978
rect 343732 117914 343784 117920
rect 344296 110430 344324 188255
rect 345032 163538 345060 316678
rect 345664 308440 345716 308446
rect 345664 308382 345716 308388
rect 345020 163532 345072 163538
rect 345020 163474 345072 163480
rect 345020 153876 345072 153882
rect 345020 153818 345072 153824
rect 344928 143608 344980 143614
rect 344928 143550 344980 143556
rect 344940 140049 344968 143550
rect 344926 140040 344982 140049
rect 344926 139975 344982 139984
rect 344284 110424 344336 110430
rect 344284 110366 344336 110372
rect 343640 101448 343692 101454
rect 343640 101390 343692 101396
rect 345032 100026 345060 153818
rect 345112 152108 345164 152114
rect 345112 152050 345164 152056
rect 345124 151910 345152 152050
rect 345112 151904 345164 151910
rect 345112 151846 345164 151852
rect 345124 127634 345152 151846
rect 345204 131776 345256 131782
rect 345204 131718 345256 131724
rect 345112 127628 345164 127634
rect 345112 127570 345164 127576
rect 345216 111110 345244 131718
rect 345204 111104 345256 111110
rect 345204 111046 345256 111052
rect 345020 100020 345072 100026
rect 345020 99962 345072 99968
rect 342904 95056 342956 95062
rect 342904 94998 342956 95004
rect 345676 93702 345704 308382
rect 346306 145888 346362 145897
rect 346306 145823 346362 145832
rect 346320 144226 346348 145823
rect 346308 144220 346360 144226
rect 346308 144162 346360 144168
rect 346412 142154 346440 378762
rect 346582 352608 346638 352617
rect 346582 352543 346638 352552
rect 346492 349852 346544 349858
rect 346492 349794 346544 349800
rect 346504 145897 346532 349794
rect 346596 190454 346624 352543
rect 348424 341556 348476 341562
rect 348424 341498 348476 341504
rect 346596 190426 346716 190454
rect 346688 166326 346716 190426
rect 347320 180192 347372 180198
rect 347320 180134 347372 180140
rect 347042 169688 347098 169697
rect 347042 169623 347098 169632
rect 347056 168434 347084 169623
rect 347044 168428 347096 168434
rect 347044 168370 347096 168376
rect 346676 166320 346728 166326
rect 346860 166320 346912 166326
rect 346676 166262 346728 166268
rect 346858 166288 346860 166297
rect 346912 166288 346914 166297
rect 346858 166223 346914 166232
rect 346676 163532 346728 163538
rect 346676 163474 346728 163480
rect 346688 162897 346716 163474
rect 346674 162888 346730 162897
rect 346674 162823 346730 162832
rect 347044 156120 347096 156126
rect 347042 156088 347044 156097
rect 347096 156088 347098 156097
rect 347042 156023 347098 156032
rect 346674 154456 346730 154465
rect 346674 154391 346730 154400
rect 346688 153882 346716 154391
rect 346676 153876 346728 153882
rect 346676 153818 346728 153824
rect 346582 152688 346638 152697
rect 346582 152623 346638 152632
rect 346596 152114 346624 152623
rect 346584 152108 346636 152114
rect 346584 152050 346636 152056
rect 346676 151768 346728 151774
rect 346676 151710 346728 151716
rect 346688 151065 346716 151710
rect 346674 151056 346730 151065
rect 346674 150991 346730 151000
rect 346674 147656 346730 147665
rect 346674 147591 346730 147600
rect 346688 146946 346716 147591
rect 346676 146940 346728 146946
rect 346676 146882 346728 146888
rect 346490 145888 346546 145897
rect 346490 145823 346546 145832
rect 346676 145580 346728 145586
rect 346676 145522 346728 145528
rect 346688 144265 346716 145522
rect 346674 144256 346730 144265
rect 346674 144191 346730 144200
rect 346688 143614 346716 144191
rect 346676 143608 346728 143614
rect 346676 143550 346728 143556
rect 346584 142860 346636 142866
rect 346584 142802 346636 142808
rect 346596 142633 346624 142802
rect 346582 142624 346638 142633
rect 346582 142559 346638 142568
rect 346412 142126 346532 142154
rect 346504 141522 346532 142126
rect 346412 141494 346532 141522
rect 346412 138718 346440 141494
rect 346492 141432 346544 141438
rect 346492 141374 346544 141380
rect 346504 140865 346532 141374
rect 346490 140856 346546 140865
rect 346490 140791 346546 140800
rect 346400 138712 346452 138718
rect 346400 138654 346452 138660
rect 346596 133210 346624 142559
rect 347134 139224 347190 139233
rect 347134 139159 347190 139168
rect 347148 138718 347176 139159
rect 347136 138712 347188 138718
rect 347136 138654 347188 138660
rect 346674 137456 346730 137465
rect 346674 137391 346730 137400
rect 346688 136746 346716 137391
rect 346676 136740 346728 136746
rect 346676 136682 346728 136688
rect 346584 133204 346636 133210
rect 346584 133146 346636 133152
rect 347044 120080 347096 120086
rect 347044 120022 347096 120028
rect 347056 118833 347084 120022
rect 347042 118824 347098 118833
rect 347042 118759 347098 118768
rect 347332 117201 347360 180134
rect 347502 174720 347558 174729
rect 347502 174655 347558 174664
rect 347516 173942 347544 174655
rect 347504 173936 347556 173942
rect 347504 173878 347556 173884
rect 347502 173088 347558 173097
rect 347502 173023 347558 173032
rect 347516 172582 347544 173023
rect 347504 172576 347556 172582
rect 347504 172518 347556 172524
rect 347502 171320 347558 171329
rect 347502 171255 347558 171264
rect 347516 171154 347544 171255
rect 347504 171148 347556 171154
rect 347504 171090 347556 171096
rect 347502 167920 347558 167929
rect 347502 167855 347558 167864
rect 347516 167074 347544 167855
rect 347504 167068 347556 167074
rect 347504 167010 347556 167016
rect 347502 164520 347558 164529
rect 347502 164455 347558 164464
rect 347516 164286 347544 164455
rect 347504 164280 347556 164286
rect 347504 164222 347556 164228
rect 347504 161424 347556 161430
rect 347504 161366 347556 161372
rect 347516 161129 347544 161366
rect 347502 161120 347558 161129
rect 347502 161055 347558 161064
rect 347502 159488 347558 159497
rect 347502 159423 347558 159432
rect 347516 159390 347544 159423
rect 347504 159384 347556 159390
rect 347504 159326 347556 159332
rect 347502 157856 347558 157865
rect 347502 157791 347558 157800
rect 347516 157486 347544 157791
rect 347504 157480 347556 157486
rect 347504 157422 347556 157428
rect 347502 149288 347558 149297
rect 347502 149223 347558 149232
rect 347516 149190 347544 149223
rect 347504 149184 347556 149190
rect 347504 149126 347556 149132
rect 347502 135824 347558 135833
rect 347502 135759 347558 135768
rect 347516 135318 347544 135759
rect 347504 135312 347556 135318
rect 347504 135254 347556 135260
rect 347410 132424 347466 132433
rect 347410 132359 347466 132368
rect 347424 131782 347452 132359
rect 347412 131776 347464 131782
rect 347412 131718 347464 131724
rect 347686 128480 347742 128489
rect 347686 128415 347742 128424
rect 347700 126954 347728 128415
rect 347964 128308 348016 128314
rect 347964 128250 348016 128256
rect 347976 127401 348004 128250
rect 347962 127392 348018 127401
rect 347962 127327 348018 127336
rect 347688 126948 347740 126954
rect 347688 126890 347740 126896
rect 347688 126268 347740 126274
rect 347688 126210 347740 126216
rect 347700 125633 347728 126210
rect 347686 125624 347742 125633
rect 347686 125559 347742 125568
rect 347318 117192 347374 117201
rect 347318 117127 347374 117136
rect 347504 115932 347556 115938
rect 347504 115874 347556 115880
rect 347516 115433 347544 115874
rect 347502 115424 347558 115433
rect 347502 115359 347558 115368
rect 347044 110424 347096 110430
rect 347042 110392 347044 110401
rect 347096 110392 347098 110401
rect 347042 110327 347098 110336
rect 347504 108996 347556 109002
rect 347504 108938 347556 108944
rect 347516 108769 347544 108938
rect 347502 108760 347558 108769
rect 347502 108695 347558 108704
rect 347504 107636 347556 107642
rect 347504 107578 347556 107584
rect 347516 107001 347544 107578
rect 347502 106992 347558 107001
rect 347502 106927 347558 106936
rect 347044 104848 347096 104854
rect 347044 104790 347096 104796
rect 347056 103601 347084 104790
rect 347042 103592 347098 103601
rect 347042 103527 347098 103536
rect 347228 102128 347280 102134
rect 347228 102070 347280 102076
rect 347240 101969 347268 102070
rect 347226 101960 347282 101969
rect 347226 101895 347282 101904
rect 347504 100700 347556 100706
rect 347504 100642 347556 100648
rect 347516 100201 347544 100642
rect 347502 100192 347558 100201
rect 347502 100127 347558 100136
rect 347504 97980 347556 97986
rect 347504 97922 347556 97928
rect 347516 96937 347544 97922
rect 347502 96928 347558 96937
rect 347502 96863 347558 96872
rect 347700 93838 347728 125559
rect 347688 93832 347740 93838
rect 347688 93774 347740 93780
rect 345664 93696 345716 93702
rect 345664 93638 345716 93644
rect 348436 92750 348464 341498
rect 349068 231872 349120 231878
rect 349068 231814 349120 231820
rect 348976 186992 349028 186998
rect 348976 186934 349028 186940
rect 348882 127392 348938 127401
rect 348882 127327 348938 127336
rect 348896 96626 348924 127327
rect 348988 124166 349016 186934
rect 348976 124160 349028 124166
rect 348976 124102 349028 124108
rect 348988 124001 349016 124102
rect 348974 123992 349030 124001
rect 348974 123927 349030 123936
rect 349080 122777 349108 231814
rect 349158 131064 349214 131073
rect 349158 130999 349214 131008
rect 349172 130665 349200 130999
rect 349158 130656 349214 130665
rect 349158 130591 349214 130600
rect 349066 122768 349122 122777
rect 349066 122703 349122 122712
rect 348884 96620 348936 96626
rect 348884 96562 348936 96568
rect 348424 92744 348476 92750
rect 348424 92686 348476 92692
rect 342352 86284 342404 86290
rect 342352 86226 342404 86232
rect 345020 86284 345072 86290
rect 345020 86226 345072 86232
rect 342260 80708 342312 80714
rect 342260 80650 342312 80656
rect 340880 41404 340932 41410
rect 340880 41346 340932 41352
rect 341524 41404 341576 41410
rect 341524 41346 341576 41352
rect 340892 3534 340920 41346
rect 340972 35216 341024 35222
rect 340972 35158 341024 35164
rect 340144 3528 340196 3534
rect 340144 3470 340196 3476
rect 340880 3528 340932 3534
rect 340880 3470 340932 3476
rect 340984 480 341012 35158
rect 342272 16574 342300 80650
rect 343638 47560 343694 47569
rect 343638 47495 343694 47504
rect 343652 16574 343680 47495
rect 345032 16574 345060 86226
rect 347780 50380 347832 50386
rect 347780 50322 347832 50328
rect 347792 16574 347820 50322
rect 349172 33114 349200 130591
rect 349816 93770 349844 381783
rect 372620 376780 372672 376786
rect 372620 376722 372672 376728
rect 349896 344344 349948 344350
rect 349896 344286 349948 344292
rect 349804 93764 349856 93770
rect 349804 93706 349856 93712
rect 349908 93634 349936 344286
rect 358084 327752 358136 327758
rect 358084 327694 358136 327700
rect 353944 303000 353996 303006
rect 353944 302942 353996 302948
rect 352564 292596 352616 292602
rect 352564 292538 352616 292544
rect 350816 185632 350868 185638
rect 350816 185574 350868 185580
rect 350828 175522 350856 185574
rect 352576 177478 352604 292538
rect 352564 177472 352616 177478
rect 352564 177414 352616 177420
rect 353300 177336 353352 177342
rect 353300 177278 353352 177284
rect 353312 175522 353340 177278
rect 353956 175982 353984 302942
rect 356060 253224 356112 253230
rect 356060 253166 356112 253172
rect 353944 175976 353996 175982
rect 353944 175918 353996 175924
rect 356072 175522 356100 253166
rect 358096 190454 358124 327694
rect 360844 287700 360896 287706
rect 360844 287642 360896 287648
rect 359462 226944 359518 226953
rect 359462 226879 359518 226888
rect 358096 190426 358216 190454
rect 358084 184204 358136 184210
rect 358084 184146 358136 184152
rect 358096 175522 358124 184146
rect 358188 178770 358216 190426
rect 359476 180198 359504 226879
rect 360856 182850 360884 287642
rect 365720 283620 365772 283626
rect 365720 283562 365772 283568
rect 363604 218748 363656 218754
rect 363604 218690 363656 218696
rect 360844 182844 360896 182850
rect 360844 182786 360896 182792
rect 361304 181484 361356 181490
rect 361304 181426 361356 181432
rect 359464 180192 359516 180198
rect 359464 180134 359516 180140
rect 358176 178764 358228 178770
rect 358176 178706 358228 178712
rect 361316 175522 361344 181426
rect 363616 177410 363644 218690
rect 363788 180260 363840 180266
rect 363788 180202 363840 180208
rect 363604 177404 363656 177410
rect 363604 177346 363656 177352
rect 363800 175522 363828 180202
rect 350828 175494 351256 175522
rect 353312 175494 353648 175522
rect 356072 175494 356132 175522
rect 358096 175494 358524 175522
rect 361008 175494 361344 175522
rect 363492 175494 363828 175522
rect 365732 175522 365760 283562
rect 371884 261520 371936 261526
rect 371884 261462 371936 261468
rect 370504 259480 370556 259486
rect 370504 259422 370556 259428
rect 367100 247784 367152 247790
rect 367100 247726 367152 247732
rect 367112 190454 367140 247726
rect 369860 196648 369912 196654
rect 369860 196590 369912 196596
rect 369872 190454 369900 196590
rect 367112 190426 367968 190454
rect 369872 190426 370452 190454
rect 367940 175522 367968 190426
rect 370424 175522 370452 190426
rect 370516 177342 370544 259422
rect 370504 177336 370556 177342
rect 370504 177278 370556 177284
rect 371896 176050 371924 261462
rect 372632 190454 372660 376722
rect 372632 190426 372844 190454
rect 371884 176044 371936 176050
rect 371884 175986 371936 175992
rect 372816 175522 372844 190426
rect 374656 184210 374684 563654
rect 377404 456816 377456 456822
rect 377404 456758 377456 456764
rect 375380 247716 375432 247722
rect 375380 247658 375432 247664
rect 374644 184204 374696 184210
rect 374644 184146 374696 184152
rect 375392 175522 375420 247658
rect 377416 234569 377444 456758
rect 379520 264240 379572 264246
rect 379520 264182 379572 264188
rect 376758 234560 376814 234569
rect 376758 234495 376814 234504
rect 377402 234560 377458 234569
rect 377402 234495 377458 234504
rect 376772 180266 376800 234495
rect 378140 228472 378192 228478
rect 378140 228414 378192 228420
rect 376760 180260 376812 180266
rect 376760 180202 376812 180208
rect 378152 175522 378180 228414
rect 379532 190454 379560 264182
rect 379532 190426 380204 190454
rect 380176 175522 380204 190426
rect 381556 185638 381584 702782
rect 386432 700330 386460 702782
rect 397472 702545 397500 703520
rect 413664 702982 413692 703520
rect 413652 702976 413704 702982
rect 413652 702918 413704 702924
rect 429856 702846 429884 703520
rect 462332 702914 462360 703520
rect 462320 702908 462372 702914
rect 462320 702850 462372 702856
rect 424968 702840 425020 702846
rect 424968 702782 425020 702788
rect 429844 702840 429896 702846
rect 429844 702782 429896 702788
rect 397458 702536 397514 702545
rect 397458 702471 397514 702480
rect 424980 700330 425008 702782
rect 478524 702778 478552 703520
rect 478512 702772 478564 702778
rect 478512 702714 478564 702720
rect 494808 702710 494836 703520
rect 494796 702704 494848 702710
rect 494796 702646 494848 702652
rect 527192 702642 527220 703520
rect 527180 702636 527232 702642
rect 527180 702578 527232 702584
rect 465724 702568 465776 702574
rect 465724 702510 465776 702516
rect 465736 700330 465764 702510
rect 543476 702506 543504 703520
rect 559668 702574 559696 703520
rect 550548 702568 550600 702574
rect 550548 702510 550600 702516
rect 559656 702568 559708 702574
rect 559656 702510 559708 702516
rect 543464 702500 543516 702506
rect 543464 702442 543516 702448
rect 550560 700330 550588 702510
rect 386420 700324 386472 700330
rect 386420 700266 386472 700272
rect 424968 700324 425020 700330
rect 424968 700266 425020 700272
rect 465724 700324 465776 700330
rect 465724 700266 465776 700272
rect 550548 700324 550600 700330
rect 550548 700266 550600 700272
rect 457444 643748 457496 643754
rect 457444 643690 457496 643696
rect 429844 575544 429896 575550
rect 429844 575486 429896 575492
rect 429856 563718 429884 575486
rect 429844 563712 429896 563718
rect 429844 563654 429896 563660
rect 405740 511284 405792 511290
rect 405740 511226 405792 511232
rect 405752 510678 405780 511226
rect 405740 510672 405792 510678
rect 405740 510614 405792 510620
rect 395344 323604 395396 323610
rect 395344 323546 395396 323552
rect 385040 236700 385092 236706
rect 385040 236642 385092 236648
rect 382280 229832 382332 229838
rect 382280 229774 382332 229780
rect 382292 190454 382320 229774
rect 385052 190454 385080 236642
rect 391940 213240 391992 213246
rect 391940 213182 391992 213188
rect 389180 209840 389232 209846
rect 389180 209782 389232 209788
rect 387800 207664 387852 207670
rect 387800 207606 387852 207612
rect 382292 190426 382688 190454
rect 385052 190426 385172 190454
rect 381544 185632 381596 185638
rect 381544 185574 381596 185580
rect 382660 175522 382688 190426
rect 385144 175522 385172 190426
rect 387812 175522 387840 207606
rect 389192 190454 389220 209782
rect 391952 190454 391980 213182
rect 394698 191040 394754 191049
rect 394698 190975 394754 190984
rect 394712 190454 394740 190975
rect 389192 190426 390048 190454
rect 391952 190426 392532 190454
rect 394712 190426 394924 190454
rect 390020 175522 390048 190426
rect 392504 175522 392532 190426
rect 394896 175522 394924 190426
rect 395356 185638 395384 323546
rect 399484 322244 399536 322250
rect 399484 322186 399536 322192
rect 395344 185632 395396 185638
rect 395344 185574 395396 185580
rect 399496 178838 399524 322186
rect 403624 307080 403676 307086
rect 403624 307022 403676 307028
rect 400864 249076 400916 249082
rect 400864 249018 400916 249024
rect 400220 217320 400272 217326
rect 400220 217262 400272 217268
rect 399484 178832 399536 178838
rect 399484 178774 399536 178780
rect 397460 177472 397512 177478
rect 397460 177414 397512 177420
rect 397472 175522 397500 177414
rect 400232 175522 400260 217262
rect 400876 182986 400904 249018
rect 401600 211812 401652 211818
rect 401600 211754 401652 211760
rect 401612 190454 401640 211754
rect 401612 190426 402284 190454
rect 400864 182980 400916 182986
rect 400864 182922 400916 182928
rect 402256 175522 402284 190426
rect 403636 176730 403664 307022
rect 405752 181490 405780 510614
rect 421564 371272 421616 371278
rect 421564 371214 421616 371220
rect 409880 331900 409932 331906
rect 409880 331842 409932 331848
rect 407764 251864 407816 251870
rect 407764 251806 407816 251812
rect 407120 214600 407172 214606
rect 407120 214542 407172 214548
rect 407132 190454 407160 214542
rect 407132 190426 407252 190454
rect 405740 181484 405792 181490
rect 405740 181426 405792 181432
rect 403624 176724 403676 176730
rect 403624 176666 403676 176672
rect 404820 176724 404872 176730
rect 404820 176666 404872 176672
rect 404832 175522 404860 176666
rect 407224 175522 407252 190426
rect 407776 180266 407804 251806
rect 407764 180260 407816 180266
rect 407764 180202 407816 180208
rect 409892 175522 409920 331842
rect 416780 303680 416832 303686
rect 416780 303622 416832 303628
rect 414664 284368 414716 284374
rect 414664 284310 414716 284316
rect 413284 242956 413336 242962
rect 413284 242898 413336 242904
rect 411260 239420 411312 239426
rect 411260 239362 411312 239368
rect 411272 180794 411300 239362
rect 411904 232552 411956 232558
rect 411904 232494 411956 232500
rect 411916 183054 411944 232494
rect 411904 183048 411956 183054
rect 411904 182990 411956 182996
rect 411272 180766 412128 180794
rect 412100 175522 412128 180766
rect 413296 177546 413324 242898
rect 414020 215960 414072 215966
rect 414020 215902 414072 215908
rect 414032 190454 414060 215902
rect 414032 190426 414612 190454
rect 413284 177540 413336 177546
rect 413284 177482 413336 177488
rect 414584 175522 414612 190426
rect 414676 180334 414704 284310
rect 416792 190454 416820 303622
rect 418804 276072 418856 276078
rect 418804 276014 418856 276020
rect 417424 222896 417476 222902
rect 417424 222838 417476 222844
rect 416792 190426 417004 190454
rect 414664 180328 414716 180334
rect 414664 180270 414716 180276
rect 416976 175522 417004 190426
rect 417436 177614 417464 222838
rect 418816 178906 418844 276014
rect 419540 275324 419592 275330
rect 419540 275266 419592 275272
rect 418896 228404 418948 228410
rect 418896 228346 418948 228352
rect 418804 178900 418856 178906
rect 418804 178842 418856 178848
rect 417424 177608 417476 177614
rect 417424 177550 417476 177556
rect 418908 177478 418936 228346
rect 418896 177472 418948 177478
rect 418896 177414 418948 177420
rect 419552 175522 419580 275266
rect 421576 176118 421604 371214
rect 425704 330540 425756 330546
rect 425704 330482 425756 330488
rect 424416 181552 424468 181558
rect 424416 181494 424468 181500
rect 422300 177404 422352 177410
rect 422300 177346 422352 177352
rect 421564 176112 421616 176118
rect 421564 176054 421616 176060
rect 422312 175522 422340 177346
rect 424428 175522 424456 181494
rect 425716 176089 425744 330482
rect 453304 311908 453356 311914
rect 453304 311850 453356 311856
rect 445760 309868 445812 309874
rect 445760 309810 445812 309816
rect 433340 309800 433392 309806
rect 433340 309742 433392 309748
rect 428464 294636 428516 294642
rect 428464 294578 428516 294584
rect 428096 199504 428148 199510
rect 428096 199446 428148 199452
rect 425796 185632 425848 185638
rect 425796 185574 425848 185580
rect 425702 176080 425758 176089
rect 425702 176015 425758 176024
rect 425808 175914 425836 185574
rect 426900 177608 426952 177614
rect 426900 177550 426952 177556
rect 425796 175908 425848 175914
rect 425796 175850 425848 175856
rect 426912 175522 426940 177550
rect 365732 175494 365884 175522
rect 367940 175494 368368 175522
rect 370424 175494 370852 175522
rect 372816 175494 373244 175522
rect 375392 175494 375728 175522
rect 378152 175494 378212 175522
rect 380176 175494 380604 175522
rect 382660 175494 383088 175522
rect 385144 175494 385572 175522
rect 387812 175494 387964 175522
rect 390020 175494 390448 175522
rect 392504 175494 392932 175522
rect 394896 175494 395324 175522
rect 397472 175494 397808 175522
rect 400232 175494 400292 175522
rect 402256 175494 402684 175522
rect 404832 175494 405168 175522
rect 407224 175494 407652 175522
rect 409892 175494 410044 175522
rect 412100 175494 412528 175522
rect 414584 175494 415012 175522
rect 416976 175494 417404 175522
rect 419552 175494 419888 175522
rect 422312 175494 422372 175522
rect 424428 175494 424764 175522
rect 426912 175494 427248 175522
rect 427818 175264 427874 175273
rect 427818 175199 427820 175208
rect 427872 175199 427874 175208
rect 427820 175170 427872 175176
rect 427910 166968 427966 166977
rect 427910 166903 427966 166912
rect 349986 128480 350042 128489
rect 349986 128415 350042 128424
rect 349896 93628 349948 93634
rect 349896 93570 349948 93576
rect 350000 73166 350028 128415
rect 350552 96070 350612 96098
rect 351472 96070 351808 96098
rect 352760 96070 353096 96098
rect 354048 96070 354384 96098
rect 355336 96070 355672 96098
rect 356532 96070 356868 96098
rect 357820 96070 358156 96098
rect 359108 96070 359444 96098
rect 360304 96070 360732 96098
rect 361592 96070 361928 96098
rect 362972 96070 363216 96098
rect 364352 96070 364504 96098
rect 365732 96070 365792 96098
rect 366652 96070 366988 96098
rect 367112 96070 368276 96098
rect 368492 96070 369564 96098
rect 369872 96070 370852 96098
rect 371252 96070 372048 96098
rect 372632 96070 373336 96098
rect 374012 96070 374624 96098
rect 375392 96070 375912 96098
rect 376772 96070 377108 96098
rect 378152 96070 378396 96098
rect 379532 96070 379684 96098
rect 380912 96070 380972 96098
rect 381372 96070 382168 96098
rect 382292 96070 383456 96098
rect 383672 96070 384744 96098
rect 385052 96070 386032 96098
rect 386432 96070 387228 96098
rect 388180 96070 388516 96098
rect 389468 96070 389804 96098
rect 390664 96070 391092 96098
rect 391952 96070 392380 96098
rect 393332 96070 393576 96098
rect 394712 96070 394864 96098
rect 396092 96070 396152 96098
rect 397104 96070 397440 96098
rect 397564 96070 398636 96098
rect 399588 96070 399924 96098
rect 400876 96070 401212 96098
rect 401612 96070 402500 96098
rect 402992 96070 403696 96098
rect 404372 96070 404984 96098
rect 406028 96070 406272 96098
rect 407132 96070 407560 96098
rect 408512 96070 408756 96098
rect 409892 96070 410044 96098
rect 411272 96070 411332 96098
rect 412284 96070 412620 96098
rect 413020 96070 413816 96098
rect 414032 96070 415104 96098
rect 415412 96070 416392 96098
rect 416792 96070 417680 96098
rect 418172 96070 418876 96098
rect 419552 96070 420164 96098
rect 420932 96070 421452 96098
rect 422312 96070 422740 96098
rect 423692 96070 423936 96098
rect 425072 96070 425224 96098
rect 426452 96070 426512 96098
rect 427464 96070 427800 96098
rect 350552 93854 350580 96070
rect 350552 93826 350672 93854
rect 349988 73160 350040 73166
rect 349988 73102 350040 73108
rect 349252 42084 349304 42090
rect 349252 42026 349304 42032
rect 349160 33108 349212 33114
rect 349160 33050 349212 33056
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 347792 16546 348096 16574
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 342180 480 342208 3470
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346952 3596 347004 3602
rect 346952 3538 347004 3544
rect 346964 480 346992 3538
rect 348068 480 348096 16546
rect 349160 4276 349212 4282
rect 349160 4218 349212 4224
rect 349172 3466 349200 4218
rect 349160 3460 349212 3466
rect 349160 3402 349212 3408
rect 349264 480 349292 42026
rect 350644 14482 350672 93826
rect 351472 93498 351500 96070
rect 351460 93492 351512 93498
rect 351460 93434 351512 93440
rect 352012 92336 352064 92342
rect 352012 92278 352064 92284
rect 352024 91798 352052 92278
rect 352760 91798 352788 96070
rect 354048 92750 354076 96070
rect 353300 92744 353352 92750
rect 353300 92686 353352 92692
rect 354036 92744 354088 92750
rect 354036 92686 354088 92692
rect 352012 91792 352064 91798
rect 352012 91734 352064 91740
rect 352748 91792 352800 91798
rect 352748 91734 352800 91740
rect 351920 89004 351972 89010
rect 351920 88946 351972 88952
rect 350632 14476 350684 14482
rect 350632 14418 350684 14424
rect 351932 3534 351960 88946
rect 352024 42226 352052 91734
rect 352012 42220 352064 42226
rect 352012 42162 352064 42168
rect 353312 4282 353340 92686
rect 355336 89078 355364 96070
rect 356532 93702 356560 96070
rect 357820 93854 357848 96070
rect 359108 93854 359136 96070
rect 360304 93854 360332 96070
rect 357452 93826 357848 93854
rect 358832 93826 359136 93854
rect 360212 93826 360332 93854
rect 356520 93696 356572 93702
rect 356520 93638 356572 93644
rect 356532 92546 356560 93638
rect 356060 92540 356112 92546
rect 356060 92482 356112 92488
rect 356520 92540 356572 92546
rect 356520 92482 356572 92488
rect 355324 89072 355376 89078
rect 355324 89014 355376 89020
rect 356072 38010 356100 92482
rect 357452 92478 357480 93826
rect 358832 93634 358860 93826
rect 360212 93770 360240 93826
rect 360200 93764 360252 93770
rect 360200 93706 360252 93712
rect 358820 93628 358872 93634
rect 358820 93570 358872 93576
rect 357440 92472 357492 92478
rect 357440 92414 357492 92420
rect 356060 38004 356112 38010
rect 356060 37946 356112 37952
rect 356704 37936 356756 37942
rect 356704 37878 356756 37884
rect 353300 4276 353352 4282
rect 353300 4218 353352 4224
rect 356716 3602 356744 37878
rect 357452 35290 357480 92414
rect 357440 35284 357492 35290
rect 357440 35226 357492 35232
rect 358832 32502 358860 93570
rect 360212 50454 360240 93706
rect 360200 50448 360252 50454
rect 360200 50390 360252 50396
rect 361592 49094 361620 96070
rect 361580 49088 361632 49094
rect 361580 49030 361632 49036
rect 358820 32496 358872 32502
rect 358820 32438 358872 32444
rect 362972 7614 363000 96070
rect 364352 47598 364380 96070
rect 365732 87650 365760 96070
rect 366652 90370 366680 96070
rect 366640 90364 366692 90370
rect 366640 90306 366692 90312
rect 365720 87644 365772 87650
rect 365720 87586 365772 87592
rect 364340 47592 364392 47598
rect 364340 47534 364392 47540
rect 367112 31074 367140 96070
rect 367100 31068 367152 31074
rect 367100 31010 367152 31016
rect 368492 29646 368520 96070
rect 368480 29640 368532 29646
rect 368480 29582 368532 29588
rect 369872 28286 369900 96070
rect 369860 28280 369912 28286
rect 369860 28222 369912 28228
rect 362960 7608 363012 7614
rect 362960 7550 363012 7556
rect 371252 6866 371280 96070
rect 372632 77994 372660 96070
rect 372620 77988 372672 77994
rect 372620 77930 372672 77936
rect 374012 25566 374040 96070
rect 374000 25560 374052 25566
rect 374000 25502 374052 25508
rect 375392 21418 375420 96070
rect 375380 21412 375432 21418
rect 375380 21354 375432 21360
rect 376772 19990 376800 96070
rect 376760 19984 376812 19990
rect 376760 19926 376812 19932
rect 378152 19310 378180 96070
rect 379532 26926 379560 96070
rect 379520 26920 379572 26926
rect 379520 26862 379572 26868
rect 378140 19304 378192 19310
rect 378140 19246 378192 19252
rect 371240 6860 371292 6866
rect 371240 6802 371292 6808
rect 380912 5506 380940 96070
rect 381372 84194 381400 96070
rect 381004 84166 381400 84194
rect 381004 24274 381032 84166
rect 380992 24268 381044 24274
rect 380992 24210 381044 24216
rect 382292 17270 382320 96070
rect 383672 22778 383700 96070
rect 383660 22772 383712 22778
rect 383660 22714 383712 22720
rect 382280 17264 382332 17270
rect 382280 17206 382332 17212
rect 385052 15910 385080 96070
rect 386432 44878 386460 96070
rect 388180 89010 388208 96070
rect 389468 95266 389496 96070
rect 389456 95260 389508 95266
rect 389456 95202 389508 95208
rect 388442 90400 388498 90409
rect 388442 90335 388498 90344
rect 388168 89004 388220 89010
rect 388168 88946 388220 88952
rect 386420 44872 386472 44878
rect 386420 44814 386472 44820
rect 385040 15904 385092 15910
rect 385040 15846 385092 15852
rect 380900 5500 380952 5506
rect 380900 5442 380952 5448
rect 356704 3596 356756 3602
rect 356704 3538 356756 3544
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 351920 3528 351972 3534
rect 351920 3470 351972 3476
rect 350460 480 350488 3470
rect 388456 3466 388484 90335
rect 389468 84194 389496 95202
rect 390664 93809 390692 96070
rect 390650 93800 390706 93809
rect 390650 93735 390706 93744
rect 390664 84194 390692 93735
rect 391952 91050 391980 96070
rect 391940 91044 391992 91050
rect 391940 90986 391992 90992
rect 389192 84166 389496 84194
rect 390572 84166 390692 84194
rect 389192 37942 389220 84166
rect 390572 80714 390600 84166
rect 390560 80708 390612 80714
rect 390560 80650 390612 80656
rect 389180 37936 389232 37942
rect 389180 37878 389232 37884
rect 391952 14550 391980 90986
rect 393332 80034 393360 96070
rect 394712 92410 394740 96070
rect 396092 92546 396120 96070
rect 397104 94994 397132 96070
rect 396172 94988 396224 94994
rect 396172 94930 396224 94936
rect 397092 94988 397144 94994
rect 397092 94930 397144 94936
rect 395344 92540 395396 92546
rect 395344 92482 395396 92488
rect 396080 92540 396132 92546
rect 396080 92482 396132 92488
rect 394700 92404 394752 92410
rect 394700 92346 394752 92352
rect 393320 80028 393372 80034
rect 393320 79970 393372 79976
rect 394712 49026 394740 92346
rect 395356 76566 395384 92482
rect 396184 84194 396212 94930
rect 396724 92540 396776 92546
rect 396724 92482 396776 92488
rect 396092 84166 396212 84194
rect 396092 82142 396120 84166
rect 396080 82136 396132 82142
rect 396080 82078 396132 82084
rect 395344 76560 395396 76566
rect 395344 76502 395396 76508
rect 396736 75886 396764 92482
rect 397564 84194 397592 96070
rect 399484 93152 399536 93158
rect 399484 93094 399536 93100
rect 397472 84166 397592 84194
rect 397472 83502 397500 84166
rect 397460 83496 397512 83502
rect 397460 83438 397512 83444
rect 396724 75880 396776 75886
rect 396724 75822 396776 75828
rect 399496 66910 399524 93094
rect 399588 92546 399616 96070
rect 400876 95062 400904 96070
rect 400220 95056 400272 95062
rect 400220 94998 400272 95004
rect 400864 95056 400916 95062
rect 400864 94998 400916 95004
rect 399576 92540 399628 92546
rect 399576 92482 399628 92488
rect 400232 73846 400260 94998
rect 400220 73840 400272 73846
rect 400220 73782 400272 73788
rect 401612 69698 401640 96070
rect 401600 69692 401652 69698
rect 401600 69634 401652 69640
rect 402992 68338 403020 96070
rect 404372 84862 404400 96070
rect 406028 93158 406056 96070
rect 406016 93152 406068 93158
rect 406016 93094 406068 93100
rect 406384 92540 406436 92546
rect 406384 92482 406436 92488
rect 404360 84856 404412 84862
rect 404360 84798 404412 84804
rect 402980 68332 403032 68338
rect 402980 68274 403032 68280
rect 399484 66904 399536 66910
rect 399484 66846 399536 66852
rect 394700 49020 394752 49026
rect 394700 48962 394752 48968
rect 391940 14544 391992 14550
rect 391940 14486 391992 14492
rect 406396 13802 406424 92482
rect 407132 66230 407160 96070
rect 408512 92546 408540 96070
rect 408500 92540 408552 92546
rect 408500 92482 408552 92488
rect 407120 66224 407172 66230
rect 407120 66166 407172 66172
rect 409892 64190 409920 96070
rect 411272 93854 411300 96070
rect 411272 93826 411392 93854
rect 410524 93152 410576 93158
rect 410524 93094 410576 93100
rect 409880 64184 409932 64190
rect 409880 64126 409932 64132
rect 410536 43586 410564 93094
rect 411260 89004 411312 89010
rect 411260 88946 411312 88952
rect 410524 43580 410576 43586
rect 410524 43522 410576 43528
rect 406384 13796 406436 13802
rect 406384 13738 406436 13744
rect 411272 12442 411300 88946
rect 411364 62830 411392 93826
rect 412284 89010 412312 96070
rect 412272 89004 412324 89010
rect 412272 88946 412324 88952
rect 413020 84194 413048 96070
rect 412652 84166 413048 84194
rect 411352 62824 411404 62830
rect 411352 62766 411404 62772
rect 412652 61402 412680 84166
rect 412640 61396 412692 61402
rect 412640 61338 412692 61344
rect 414032 60042 414060 96070
rect 414020 60036 414072 60042
rect 414020 59978 414072 59984
rect 415412 58682 415440 96070
rect 415400 58676 415452 58682
rect 415400 58618 415452 58624
rect 416792 57254 416820 96070
rect 416780 57248 416832 57254
rect 416780 57190 416832 57196
rect 411260 12436 411312 12442
rect 411260 12378 411312 12384
rect 418172 8974 418200 96070
rect 419552 55894 419580 96070
rect 419540 55888 419592 55894
rect 419540 55830 419592 55836
rect 420932 10334 420960 96070
rect 422312 54534 422340 96070
rect 422300 54528 422352 54534
rect 422300 54470 422352 54476
rect 423692 53106 423720 96070
rect 423680 53100 423732 53106
rect 423680 53042 423732 53048
rect 425072 51814 425100 96070
rect 426452 93854 426480 96070
rect 426452 93826 426572 93854
rect 425060 51808 425112 51814
rect 425060 51750 425112 51756
rect 426544 46306 426572 93826
rect 427464 93158 427492 96070
rect 427634 95976 427690 95985
rect 427634 95911 427690 95920
rect 427648 95198 427676 95911
rect 427636 95192 427688 95198
rect 427636 95134 427688 95140
rect 427452 93152 427504 93158
rect 427452 93094 427504 93100
rect 426532 46300 426584 46306
rect 426532 46242 426584 46248
rect 427924 41410 427952 166903
rect 428002 165744 428058 165753
rect 428002 165679 428058 165688
rect 428016 86290 428044 165679
rect 428108 126313 428136 199446
rect 428476 133793 428504 294578
rect 430948 271176 431000 271182
rect 430948 271118 431000 271124
rect 430762 231160 430818 231169
rect 430762 231095 430818 231104
rect 429476 204944 429528 204950
rect 429476 204886 429528 204892
rect 429384 178832 429436 178838
rect 429384 178774 429436 178780
rect 429292 175908 429344 175914
rect 429292 175850 429344 175856
rect 429198 173360 429254 173369
rect 429198 173295 429254 173304
rect 429108 166864 429160 166870
rect 429108 166806 429160 166812
rect 429120 166161 429148 166806
rect 429106 166152 429162 166161
rect 429106 166087 429162 166096
rect 428462 133784 428518 133793
rect 428462 133719 428518 133728
rect 428094 126304 428150 126313
rect 428094 126239 428150 126248
rect 428094 99376 428150 99385
rect 428094 99311 428150 99320
rect 428108 96558 428136 99311
rect 428186 98288 428242 98297
rect 428186 98223 428242 98232
rect 428096 96552 428148 96558
rect 428096 96494 428148 96500
rect 428200 95130 428228 98223
rect 428188 95124 428240 95130
rect 428188 95066 428240 95072
rect 428004 86284 428056 86290
rect 428004 86226 428056 86232
rect 427912 41404 427964 41410
rect 427912 41346 427964 41352
rect 429212 37262 429240 173295
rect 429304 168881 429332 175850
rect 429396 172281 429424 178774
rect 429382 172272 429438 172281
rect 429382 172207 429438 172216
rect 429396 171193 429424 172207
rect 429382 171184 429438 171193
rect 429382 171119 429438 171128
rect 429290 168872 429346 168881
rect 429290 168807 429346 168816
rect 429290 167784 429346 167793
rect 429290 167719 429346 167728
rect 429304 40050 429332 167719
rect 429382 140856 429438 140865
rect 429382 140791 429438 140800
rect 429292 40044 429344 40050
rect 429292 39986 429344 39992
rect 429200 37256 429252 37262
rect 429200 37198 429252 37204
rect 429396 34474 429424 140791
rect 429488 138961 429516 204886
rect 430580 178696 430632 178702
rect 430580 178638 430632 178644
rect 430592 173233 430620 178638
rect 430672 176112 430724 176118
rect 430672 176054 430724 176060
rect 430578 173224 430634 173233
rect 430578 173159 430634 173168
rect 430592 172582 430620 173159
rect 430580 172576 430632 172582
rect 430580 172518 430632 172524
rect 430684 169969 430712 176054
rect 430670 169960 430726 169969
rect 430670 169895 430726 169904
rect 430670 165064 430726 165073
rect 430670 164999 430726 165008
rect 430580 164212 430632 164218
rect 430580 164154 430632 164160
rect 430592 163985 430620 164154
rect 430578 163976 430634 163985
rect 430578 163911 430634 163920
rect 430580 162852 430632 162858
rect 430580 162794 430632 162800
rect 430592 162489 430620 162794
rect 430578 162480 430634 162489
rect 430578 162415 430634 162424
rect 430580 162240 430632 162246
rect 430580 162182 430632 162188
rect 430592 161945 430620 162182
rect 430578 161936 430634 161945
rect 430578 161871 430634 161880
rect 430580 161424 430632 161430
rect 430580 161366 430632 161372
rect 430592 160993 430620 161366
rect 430578 160984 430634 160993
rect 430578 160919 430634 160928
rect 430580 160064 430632 160070
rect 430580 160006 430632 160012
rect 430592 159769 430620 160006
rect 430578 159760 430634 159769
rect 430578 159695 430634 159704
rect 430580 158704 430632 158710
rect 430580 158646 430632 158652
rect 430592 158545 430620 158646
rect 430578 158536 430634 158545
rect 430578 158471 430634 158480
rect 430580 157344 430632 157350
rect 430580 157286 430632 157292
rect 430592 157185 430620 157286
rect 430578 157176 430634 157185
rect 430578 157111 430634 157120
rect 430580 155848 430632 155854
rect 430580 155790 430632 155796
rect 430592 155689 430620 155790
rect 430578 155680 430634 155689
rect 430578 155615 430634 155624
rect 430580 154556 430632 154562
rect 430580 154498 430632 154504
rect 430592 154193 430620 154498
rect 430578 154184 430634 154193
rect 430578 154119 430634 154128
rect 430580 153196 430632 153202
rect 430580 153138 430632 153144
rect 430592 152833 430620 153138
rect 430578 152824 430634 152833
rect 430578 152759 430634 152768
rect 430580 151768 430632 151774
rect 430580 151710 430632 151716
rect 430592 151609 430620 151710
rect 430578 151600 430634 151609
rect 430578 151535 430634 151544
rect 430580 150408 430632 150414
rect 430580 150350 430632 150356
rect 430592 150113 430620 150350
rect 430578 150104 430634 150113
rect 430578 150039 430634 150048
rect 430580 149048 430632 149054
rect 430580 148990 430632 148996
rect 430592 148617 430620 148990
rect 430578 148608 430634 148617
rect 430578 148543 430634 148552
rect 430580 146260 430632 146266
rect 430580 146202 430632 146208
rect 430592 146033 430620 146202
rect 430578 146024 430634 146033
rect 430578 145959 430634 145968
rect 430580 144900 430632 144906
rect 430580 144842 430632 144848
rect 430592 144537 430620 144842
rect 430578 144528 430634 144537
rect 430578 144463 430634 144472
rect 430578 142216 430634 142225
rect 430578 142151 430580 142160
rect 430632 142151 430634 142160
rect 430580 142122 430632 142128
rect 430580 140752 430632 140758
rect 430580 140694 430632 140700
rect 430592 140593 430620 140694
rect 430578 140584 430634 140593
rect 430578 140519 430634 140528
rect 429474 138952 429530 138961
rect 429474 138887 429530 138896
rect 429750 138952 429806 138961
rect 429750 138887 429806 138896
rect 429764 138038 429792 138887
rect 429752 138032 429804 138038
rect 429752 137974 429804 137980
rect 430578 137728 430634 137737
rect 430578 137663 430634 137672
rect 430592 137290 430620 137663
rect 430580 137284 430632 137290
rect 430580 137226 430632 137232
rect 430580 136604 430632 136610
rect 430580 136546 430632 136552
rect 430592 136377 430620 136546
rect 430578 136368 430634 136377
rect 430578 136303 430634 136312
rect 430580 135244 430632 135250
rect 430580 135186 430632 135192
rect 430592 135017 430620 135186
rect 430578 135008 430634 135017
rect 430578 134943 430634 134952
rect 430580 133884 430632 133890
rect 430580 133826 430632 133832
rect 430592 133793 430620 133826
rect 430578 133784 430634 133793
rect 430578 133719 430634 133728
rect 430580 132456 430632 132462
rect 430580 132398 430632 132404
rect 430592 132161 430620 132398
rect 430578 132152 430634 132161
rect 430578 132087 430634 132096
rect 430580 129736 430632 129742
rect 430580 129678 430632 129684
rect 430592 129441 430620 129678
rect 430578 129432 430634 129441
rect 430578 129367 430634 129376
rect 430580 125588 430632 125594
rect 430580 125530 430632 125536
rect 430592 125089 430620 125530
rect 430578 125080 430634 125089
rect 430578 125015 430634 125024
rect 430580 124160 430632 124166
rect 430580 124102 430632 124108
rect 430592 123865 430620 124102
rect 430578 123856 430634 123865
rect 430578 123791 430634 123800
rect 430580 122800 430632 122806
rect 430580 122742 430632 122748
rect 430592 122641 430620 122742
rect 430578 122632 430634 122641
rect 430578 122567 430634 122576
rect 430580 121440 430632 121446
rect 430578 121408 430580 121417
rect 430632 121408 430634 121417
rect 430578 121343 430634 121352
rect 430580 120896 430632 120902
rect 430580 120838 430632 120844
rect 430592 120601 430620 120838
rect 430578 120592 430634 120601
rect 430578 120527 430634 120536
rect 430580 119944 430632 119950
rect 430580 119886 430632 119892
rect 430592 119513 430620 119886
rect 430578 119504 430634 119513
rect 430578 119439 430634 119448
rect 430580 118448 430632 118454
rect 430580 118390 430632 118396
rect 430592 118153 430620 118390
rect 430578 118144 430634 118153
rect 430578 118079 430634 118088
rect 430580 117292 430632 117298
rect 430580 117234 430632 117240
rect 430592 117065 430620 117234
rect 430578 117056 430634 117065
rect 430578 116991 430634 117000
rect 430580 115932 430632 115938
rect 430580 115874 430632 115880
rect 430592 115841 430620 115874
rect 430578 115832 430634 115841
rect 430578 115767 430634 115776
rect 430580 114436 430632 114442
rect 430580 114378 430632 114384
rect 430592 114209 430620 114378
rect 430578 114200 430634 114209
rect 430578 114135 430634 114144
rect 430580 111784 430632 111790
rect 430580 111726 430632 111732
rect 430592 111489 430620 111726
rect 430578 111480 430634 111489
rect 430578 111415 430634 111424
rect 430578 109032 430634 109041
rect 430578 108967 430580 108976
rect 430632 108967 430634 108976
rect 430580 108938 430632 108944
rect 430580 107636 430632 107642
rect 430580 107578 430632 107584
rect 430592 107137 430620 107578
rect 430578 107128 430634 107137
rect 430578 107063 430634 107072
rect 430580 106276 430632 106282
rect 430580 106218 430632 106224
rect 430592 105913 430620 106218
rect 430578 105904 430634 105913
rect 430578 105839 430634 105848
rect 430580 104848 430632 104854
rect 430580 104790 430632 104796
rect 430592 104689 430620 104790
rect 430578 104680 430634 104689
rect 430578 104615 430634 104624
rect 430580 103488 430632 103494
rect 430578 103456 430580 103465
rect 430632 103456 430634 103465
rect 430578 103391 430634 103400
rect 430580 102128 430632 102134
rect 430580 102070 430632 102076
rect 430592 101561 430620 102070
rect 430578 101552 430634 101561
rect 430578 101487 430634 101496
rect 430580 97980 430632 97986
rect 430580 97922 430632 97928
rect 430592 97889 430620 97922
rect 430578 97880 430634 97889
rect 430578 97815 430634 97824
rect 430684 42090 430712 164999
rect 430776 112713 430804 231095
rect 430856 155916 430908 155922
rect 430856 155858 430908 155864
rect 430868 155417 430896 155858
rect 430854 155408 430910 155417
rect 430854 155343 430910 155352
rect 430960 151814 430988 271118
rect 432144 260160 432196 260166
rect 432144 260102 432196 260108
rect 431960 246356 432012 246362
rect 431960 246298 432012 246304
rect 430960 151786 431172 151814
rect 430856 150340 430908 150346
rect 430856 150282 430908 150288
rect 430868 149841 430896 150282
rect 430854 149832 430910 149841
rect 430854 149767 430910 149776
rect 430856 144832 430908 144838
rect 430856 144774 430908 144780
rect 430868 144129 430896 144774
rect 430854 144120 430910 144129
rect 430854 144055 430910 144064
rect 430856 137964 430908 137970
rect 430856 137906 430908 137912
rect 430868 137465 430896 137906
rect 430854 137456 430910 137465
rect 430854 137391 430910 137400
rect 431144 136610 431172 151786
rect 431132 136604 431184 136610
rect 431132 136546 431184 136552
rect 430856 132388 430908 132394
rect 430856 132330 430908 132336
rect 430868 131889 430896 132330
rect 430854 131880 430910 131889
rect 430854 131815 430910 131824
rect 430856 114504 430908 114510
rect 430856 114446 430908 114452
rect 430868 113937 430896 114446
rect 430854 113928 430910 113937
rect 430854 113863 430910 113872
rect 430762 112704 430818 112713
rect 430762 112639 430818 112648
rect 431866 110392 431922 110401
rect 431972 110378 432000 246298
rect 432050 169960 432106 169969
rect 432050 169895 432106 169904
rect 431922 110350 432000 110378
rect 431866 110327 431922 110336
rect 430764 103420 430816 103426
rect 430764 103362 430816 103368
rect 430776 102785 430804 103362
rect 430762 102776 430818 102785
rect 430762 102711 430818 102720
rect 432064 50386 432092 169895
rect 432156 147529 432184 260102
rect 432236 199436 432288 199442
rect 432236 199378 432288 199384
rect 432142 147520 432198 147529
rect 432142 147455 432198 147464
rect 432248 118454 432276 199378
rect 433352 120902 433380 309742
rect 439504 298172 439556 298178
rect 439504 298114 439556 298120
rect 433524 242208 433576 242214
rect 433524 242150 433576 242156
rect 433432 178764 433484 178770
rect 433432 178706 433484 178712
rect 433444 166870 433472 178706
rect 433432 166864 433484 166870
rect 433432 166806 433484 166812
rect 433340 120896 433392 120902
rect 433340 120838 433392 120844
rect 433536 119950 433564 242150
rect 434720 238060 434772 238066
rect 434720 238002 434772 238008
rect 433616 172576 433668 172582
rect 433616 172518 433668 172524
rect 433524 119944 433576 119950
rect 433524 119886 433576 119892
rect 432236 118448 432288 118454
rect 432236 118390 432288 118396
rect 432052 50380 432104 50386
rect 432052 50322 432104 50328
rect 430672 42084 430724 42090
rect 430672 42026 430724 42032
rect 433628 35222 433656 172518
rect 434732 109002 434760 238002
rect 438952 224936 439004 224942
rect 438952 224878 439004 224884
rect 438964 224534 438992 224878
rect 439516 224534 439544 298114
rect 443000 231124 443052 231130
rect 443000 231066 443052 231072
rect 438952 224528 439004 224534
rect 438952 224470 439004 224476
rect 439504 224528 439556 224534
rect 439504 224470 439556 224476
rect 437572 195424 437624 195430
rect 437572 195366 437624 195372
rect 436100 195288 436152 195294
rect 436100 195230 436152 195236
rect 434812 192568 434864 192574
rect 434812 192510 434864 192516
rect 434824 115938 434852 192510
rect 434904 182912 434956 182918
rect 434904 182854 434956 182860
rect 434916 149054 434944 182854
rect 434996 177540 435048 177546
rect 434996 177482 435048 177488
rect 435008 162858 435036 177482
rect 434996 162852 435048 162858
rect 434996 162794 435048 162800
rect 436008 162852 436060 162858
rect 436008 162794 436060 162800
rect 436020 162178 436048 162794
rect 436008 162172 436060 162178
rect 436008 162114 436060 162120
rect 436112 150346 436140 195230
rect 436376 189780 436428 189786
rect 436376 189722 436428 189728
rect 436192 178900 436244 178906
rect 436192 178842 436244 178848
rect 436100 150340 436152 150346
rect 436100 150282 436152 150288
rect 434904 149048 434956 149054
rect 434904 148990 434956 148996
rect 436100 142180 436152 142186
rect 436100 142122 436152 142128
rect 434812 115932 434864 115938
rect 434812 115874 434864 115880
rect 434720 108996 434772 109002
rect 434720 108938 434772 108944
rect 436112 71738 436140 142122
rect 436204 137222 436232 178842
rect 436284 175976 436336 175982
rect 436284 175918 436336 175924
rect 436296 146266 436324 175918
rect 436388 164218 436416 189722
rect 437480 180192 437532 180198
rect 437480 180134 437532 180140
rect 436376 164212 436428 164218
rect 436376 164154 436428 164160
rect 436652 164212 436704 164218
rect 436652 164154 436704 164160
rect 436664 163538 436692 164154
rect 436652 163532 436704 163538
rect 436652 163474 436704 163480
rect 436284 146260 436336 146266
rect 436284 146202 436336 146208
rect 436744 138712 436796 138718
rect 436744 138654 436796 138660
rect 436652 138032 436704 138038
rect 436652 137974 436704 137980
rect 436664 137290 436692 137974
rect 436756 137970 436784 138654
rect 436744 137964 436796 137970
rect 436744 137906 436796 137912
rect 436652 137284 436704 137290
rect 436652 137226 436704 137232
rect 436192 137216 436244 137222
rect 436192 137158 436244 137164
rect 436744 137216 436796 137222
rect 436744 137158 436796 137164
rect 436756 100706 436784 137158
rect 437492 103426 437520 180134
rect 437584 121446 437612 195366
rect 438860 180124 438912 180130
rect 438860 180066 438912 180072
rect 437664 177336 437716 177342
rect 437664 177278 437716 177284
rect 437676 150414 437704 177278
rect 437664 150408 437716 150414
rect 437664 150350 437716 150356
rect 437572 121440 437624 121446
rect 437572 121382 437624 121388
rect 438872 106282 438900 180066
rect 438964 155854 438992 224470
rect 440240 221468 440292 221474
rect 440240 221410 440292 221416
rect 439136 203584 439188 203590
rect 439136 203526 439188 203532
rect 439044 180260 439096 180266
rect 439044 180202 439096 180208
rect 438952 155848 439004 155854
rect 438952 155790 439004 155796
rect 439056 125594 439084 180202
rect 439148 162246 439176 203526
rect 439136 162240 439188 162246
rect 439136 162182 439188 162188
rect 439148 161474 439176 162182
rect 439148 161446 439544 161474
rect 439044 125588 439096 125594
rect 439044 125530 439096 125536
rect 438860 106276 438912 106282
rect 438860 106218 438912 106224
rect 437480 103420 437532 103426
rect 437480 103362 437532 103368
rect 436744 100700 436796 100706
rect 436744 100642 436796 100648
rect 439516 86970 439544 161446
rect 440252 132394 440280 221410
rect 441712 189100 441764 189106
rect 441712 189042 441764 189048
rect 441620 177472 441672 177478
rect 441620 177414 441672 177420
rect 440332 176044 440384 176050
rect 440332 175986 440384 175992
rect 440240 132388 440292 132394
rect 440240 132330 440292 132336
rect 440344 103494 440372 175986
rect 440422 175944 440478 175953
rect 440422 175879 440478 175888
rect 440436 144838 440464 175879
rect 440424 144832 440476 144838
rect 440424 144774 440476 144780
rect 441632 104854 441660 177414
rect 441724 144906 441752 189042
rect 441712 144900 441764 144906
rect 441712 144842 441764 144848
rect 443012 107642 443040 231066
rect 443092 200796 443144 200802
rect 443092 200738 443144 200744
rect 443000 107636 443052 107642
rect 443000 107578 443052 107584
rect 441620 104848 441672 104854
rect 441620 104790 441672 104796
rect 440332 103488 440384 103494
rect 440332 103430 440384 103436
rect 443104 97986 443132 200738
rect 443184 183048 443236 183054
rect 443184 182990 443236 182996
rect 443196 124166 443224 182990
rect 444472 182844 444524 182850
rect 444472 182786 444524 182792
rect 444380 180328 444432 180334
rect 444380 180270 444432 180276
rect 444392 129742 444420 180270
rect 444484 161430 444512 182786
rect 444472 161424 444524 161430
rect 444472 161366 444524 161372
rect 444484 160138 444512 161366
rect 444472 160132 444524 160138
rect 444472 160074 444524 160080
rect 445772 140758 445800 309810
rect 450544 300892 450596 300898
rect 450544 300834 450596 300840
rect 448520 272536 448572 272542
rect 448520 272478 448572 272484
rect 446404 235340 446456 235346
rect 446404 235282 446456 235288
rect 446416 218754 446444 235282
rect 446404 218748 446456 218754
rect 446404 218690 446456 218696
rect 445852 184340 445904 184346
rect 445852 184282 445904 184288
rect 445760 140752 445812 140758
rect 445760 140694 445812 140700
rect 445772 140078 445800 140694
rect 445760 140072 445812 140078
rect 445760 140014 445812 140020
rect 444380 129736 444432 129742
rect 444380 129678 444432 129684
rect 443184 124160 443236 124166
rect 443184 124102 443236 124108
rect 445864 114442 445892 184282
rect 446416 135250 446444 218690
rect 447140 193860 447192 193866
rect 447140 193802 447192 193808
rect 446404 135244 446456 135250
rect 446404 135186 446456 135192
rect 447152 114510 447180 193802
rect 447784 160132 447836 160138
rect 447784 160074 447836 160080
rect 447796 126954 447824 160074
rect 447784 126948 447836 126954
rect 447784 126890 447836 126896
rect 447140 114504 447192 114510
rect 447140 114446 447192 114452
rect 445852 114436 445904 114442
rect 445852 114378 445904 114384
rect 448532 102134 448560 272478
rect 450556 206310 450584 300834
rect 453316 289134 453344 311850
rect 452660 289128 452712 289134
rect 452660 289070 452712 289076
rect 453304 289128 453356 289134
rect 453304 289070 453356 289076
rect 450544 206304 450596 206310
rect 450544 206246 450596 206252
rect 448612 185768 448664 185774
rect 448612 185710 448664 185716
rect 448624 117298 448652 185710
rect 449900 182980 449952 182986
rect 449900 182922 449952 182928
rect 449912 122806 449940 182922
rect 450556 158710 450584 206246
rect 451280 192500 451332 192506
rect 451280 192442 451332 192448
rect 450544 158704 450596 158710
rect 450544 158646 450596 158652
rect 449900 122800 449952 122806
rect 449900 122742 449952 122748
rect 448612 117292 448664 117298
rect 448612 117234 448664 117240
rect 451292 111790 451320 192442
rect 452672 132462 452700 289070
rect 454040 262268 454092 262274
rect 454040 262210 454092 262216
rect 454052 160070 454080 262210
rect 454040 160064 454092 160070
rect 454040 160006 454092 160012
rect 457456 153202 457484 643690
rect 460940 257372 460992 257378
rect 460940 257314 460992 257320
rect 457444 153196 457496 153202
rect 457444 153138 457496 153144
rect 460952 138718 460980 257314
rect 464344 162172 464396 162178
rect 464344 162114 464396 162120
rect 461676 139392 461728 139398
rect 461676 139334 461728 139340
rect 461688 138718 461716 139334
rect 460940 138712 460992 138718
rect 460940 138654 460992 138660
rect 461676 138712 461728 138718
rect 461676 138654 461728 138660
rect 452660 132456 452712 132462
rect 452660 132398 452712 132404
rect 451280 111784 451332 111790
rect 451280 111726 451332 111732
rect 448520 102128 448572 102134
rect 448520 102070 448572 102076
rect 443092 97980 443144 97986
rect 443092 97922 443144 97928
rect 439504 86964 439556 86970
rect 439504 86906 439556 86912
rect 436100 71732 436152 71738
rect 436100 71674 436152 71680
rect 464356 46918 464384 162114
rect 465736 151774 465764 700266
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 579618 683904 579674 683913
rect 579618 683839 579674 683848
rect 579632 683194 579660 683839
rect 579620 683188 579672 683194
rect 579620 683130 579672 683136
rect 579620 670744 579672 670750
rect 579988 670744 580040 670750
rect 579620 670686 579672 670692
rect 579986 670712 579988 670721
rect 580040 670712 580042 670721
rect 579632 643754 579660 670686
rect 579986 670647 580042 670656
rect 579620 643748 579672 643754
rect 579620 643690 579672 643696
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580276 594114 580304 697167
rect 580354 644056 580410 644065
rect 580354 643991 580410 644000
rect 580368 620265 580396 643991
rect 580354 620256 580410 620265
rect 580354 620191 580410 620200
rect 580354 617536 580410 617545
rect 580354 617471 580410 617480
rect 580264 594108 580316 594114
rect 580264 594050 580316 594056
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 556804 590708 556856 590714
rect 556804 590650 556856 590656
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 556816 554062 556844 590650
rect 580172 582412 580224 582418
rect 580172 582354 580224 582360
rect 580184 577697 580212 582354
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563718 580212 564295
rect 580172 563712 580224 563718
rect 580172 563654 580224 563660
rect 556804 554056 556856 554062
rect 556804 553998 556856 554004
rect 580368 538898 580396 617471
rect 580356 538892 580408 538898
rect 580356 538834 580408 538840
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 579804 525768 579856 525774
rect 579804 525710 579856 525716
rect 579816 524521 579844 525710
rect 579802 524512 579858 524521
rect 579802 524447 579858 524456
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580906 491328 580962 491337
rect 580906 491263 580962 491272
rect 580920 484673 580948 491263
rect 580906 484664 580962 484673
rect 580906 484599 580962 484608
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580908 431996 580960 432002
rect 580908 431938 580960 431944
rect 580920 431633 580948 431938
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580262 428496 580318 428505
rect 580262 428431 580318 428440
rect 580276 418305 580304 428431
rect 580262 418296 580318 418305
rect 580262 418231 580318 418240
rect 579618 404968 579674 404977
rect 579618 404903 579674 404912
rect 579632 404394 579660 404903
rect 579620 404388 579672 404394
rect 579620 404330 579672 404336
rect 579632 367810 579660 404330
rect 580262 378448 580318 378457
rect 580262 378383 580318 378392
rect 479524 367804 479576 367810
rect 479524 367746 479576 367752
rect 579620 367804 579672 367810
rect 579620 367746 579672 367752
rect 475384 192500 475436 192506
rect 475384 192442 475436 192448
rect 468484 178084 468536 178090
rect 468484 178026 468536 178032
rect 467104 164892 467156 164898
rect 467104 164834 467156 164840
rect 467116 160070 467144 164834
rect 467104 160064 467156 160070
rect 467104 160006 467156 160012
rect 465724 151768 465776 151774
rect 465724 151710 465776 151716
rect 468496 136610 468524 178026
rect 471244 163532 471296 163538
rect 471244 163474 471296 163480
rect 468484 136604 468536 136610
rect 468484 136546 468536 136552
rect 464344 46912 464396 46918
rect 464344 46854 464396 46860
rect 433616 35216 433668 35222
rect 433616 35158 433668 35164
rect 429384 34468 429436 34474
rect 429384 34410 429436 34416
rect 420920 10328 420972 10334
rect 420920 10270 420972 10276
rect 418160 8968 418212 8974
rect 418160 8910 418212 8916
rect 471256 6866 471284 163474
rect 475396 157350 475424 192442
rect 475384 157344 475436 157350
rect 475384 157286 475436 157292
rect 479536 154562 479564 367746
rect 579620 366376 579672 366382
rect 579620 366318 579672 366324
rect 579632 352578 579660 366318
rect 579802 365120 579858 365129
rect 579802 365055 579858 365064
rect 579816 364410 579844 365055
rect 579804 364404 579856 364410
rect 579804 364346 579856 364352
rect 580276 355366 580304 378383
rect 580264 355360 580316 355366
rect 580264 355302 580316 355308
rect 482284 352572 482336 352578
rect 482284 352514 482336 352520
rect 579620 352572 579672 352578
rect 579620 352514 579672 352520
rect 482296 155922 482324 352514
rect 579632 351937 579660 352514
rect 579618 351928 579674 351937
rect 579618 351863 579674 351872
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580276 306338 580304 325207
rect 580264 306332 580316 306338
rect 580264 306274 580316 306280
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580262 272232 580318 272241
rect 580262 272167 580318 272176
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 485044 258120 485096 258126
rect 485044 258062 485096 258068
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 482284 155916 482336 155922
rect 482284 155858 482336 155864
rect 479524 154556 479576 154562
rect 479524 154498 479576 154504
rect 485056 133890 485084 258062
rect 579986 245576 580042 245585
rect 579986 245511 580042 245520
rect 580000 244322 580028 245511
rect 579620 244316 579672 244322
rect 579620 244258 579672 244264
rect 579988 244316 580040 244322
rect 579988 244258 580040 244264
rect 579632 192506 579660 244258
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580184 231878 580212 232319
rect 580172 231872 580224 231878
rect 580172 231814 580224 231820
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218754 580212 218991
rect 580172 218748 580224 218754
rect 580172 218690 580224 218696
rect 580172 206304 580224 206310
rect 580172 206246 580224 206252
rect 580184 205737 580212 206246
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 579620 192500 579672 192506
rect 579620 192442 579672 192448
rect 580276 188329 580304 272167
rect 580906 192536 580962 192545
rect 580906 192471 580962 192480
rect 580262 188320 580318 188329
rect 580262 188255 580318 188264
rect 580920 186998 580948 192471
rect 580908 186992 580960 186998
rect 580908 186934 580960 186940
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 164898 580212 165815
rect 580172 164892 580224 164898
rect 580172 164834 580224 164840
rect 582378 152688 582434 152697
rect 582378 152623 582434 152632
rect 493324 140072 493376 140078
rect 493324 140014 493376 140020
rect 485044 133884 485096 133890
rect 485044 133826 485096 133832
rect 493336 20670 493364 140014
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580264 137284 580316 137290
rect 580264 137226 580316 137232
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580276 59673 580304 137226
rect 580354 112840 580410 112849
rect 580354 112775 580410 112784
rect 580368 96626 580396 112775
rect 580356 96620 580408 96626
rect 580356 96562 580408 96568
rect 582392 93838 582420 152623
rect 582380 93832 582432 93838
rect 582380 93774 582432 93780
rect 580262 59664 580318 59673
rect 580262 59599 580318 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 493324 20664 493376 20670
rect 493324 20606 493376 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 471244 6860 471296 6866
rect 471244 6802 471296 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 351644 3460 351696 3466
rect 351644 3402 351696 3408
rect 388444 3460 388496 3466
rect 388444 3402 388496 3408
rect 351656 480 351684 3402
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3514 671200 3570 671256
rect 3514 658144 3570 658200
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3330 579944 3386 580000
rect 3238 566888 3294 566944
rect 3422 553832 3478 553888
rect 3146 527856 3202 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3422 501744 3478 501800
rect 3422 475632 3478 475688
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 3422 449520 3478 449576
rect 32954 458768 33010 458824
rect 3514 423544 3570 423600
rect 3422 410488 3478 410544
rect 3422 397432 3478 397488
rect 3238 371320 3294 371376
rect 3330 358400 3386 358456
rect 2778 345344 2834 345400
rect 3238 319232 3294 319288
rect 3422 306212 3424 306232
rect 3424 306212 3476 306232
rect 3476 306212 3478 306232
rect 3422 306176 3478 306212
rect 29642 298288 29698 298344
rect 2778 293156 2780 293176
rect 2780 293156 2832 293176
rect 2832 293156 2834 293176
rect 2778 293120 2834 293156
rect 3422 267144 3478 267200
rect 3146 254088 3202 254144
rect 3146 241032 3202 241088
rect 3330 214920 3386 214976
rect 3330 201864 3386 201920
rect 3422 188808 3478 188864
rect 3422 162832 3478 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 2778 97552 2834 97608
rect 3146 84632 3202 84688
rect 9678 73752 9734 73808
rect 3422 71576 3478 71632
rect 18 69536 74 69592
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3238 32408 3294 32464
rect 3422 19352 3478 19408
rect 2870 17176 2926 17232
rect 8298 36488 8354 36544
rect 3422 6432 3478 6488
rect 23478 42064 23534 42120
rect 35714 451152 35770 451208
rect 39854 273400 39910 273456
rect 41326 392536 41382 392592
rect 41234 333920 41290 333976
rect 42706 454688 42762 454744
rect 43902 383152 43958 383208
rect 46754 537376 46810 537432
rect 45282 339632 45338 339688
rect 50894 583888 50950 583944
rect 48134 446392 48190 446448
rect 49422 449928 49478 449984
rect 41326 181328 41382 181384
rect 51906 387096 51962 387152
rect 50710 246880 50766 246936
rect 49698 72392 49754 72448
rect 38658 32408 38714 32464
rect 42798 26832 42854 26888
rect 52366 387096 52422 387152
rect 53746 482840 53802 482896
rect 53102 338000 53158 338056
rect 54942 386552 54998 386608
rect 57702 583752 57758 583808
rect 53470 190984 53526 191040
rect 57702 493348 57704 493368
rect 57704 493348 57756 493368
rect 57756 493348 57758 493368
rect 57702 493312 57758 493348
rect 56598 387776 56654 387832
rect 57702 453872 57758 453928
rect 58622 492632 58678 492688
rect 57886 438096 57942 438152
rect 56322 300056 56378 300112
rect 59266 480800 59322 480856
rect 58990 406952 59046 407008
rect 58990 405728 59046 405784
rect 58530 388320 58586 388376
rect 60462 469104 60518 469160
rect 60462 467880 60518 467936
rect 60186 365880 60242 365936
rect 56506 195200 56562 195256
rect 61750 445748 61752 445768
rect 61752 445748 61804 445768
rect 61804 445748 61806 445768
rect 61750 445712 61806 445748
rect 60646 334056 60702 334112
rect 63222 447344 63278 447400
rect 63498 491292 63554 491328
rect 63498 491272 63500 491292
rect 63500 491272 63552 491292
rect 63552 491272 63554 491292
rect 64418 437552 64474 437608
rect 64418 431976 64474 432032
rect 64510 431840 64566 431896
rect 64510 422320 64566 422376
rect 64510 412528 64566 412584
rect 64510 403008 64566 403064
rect 64510 400288 64566 400344
rect 61474 301416 61530 301472
rect 62026 265668 62082 265704
rect 62026 265648 62028 265668
rect 62028 265648 62080 265668
rect 62080 265648 62082 265668
rect 63314 179968 63370 180024
rect 64694 460808 64750 460864
rect 64694 451424 64750 451480
rect 64786 451152 64842 451208
rect 64786 447072 64842 447128
rect 67638 581304 67694 581360
rect 67822 580624 67878 580680
rect 67362 579128 67418 579184
rect 65614 466112 65670 466168
rect 65154 379480 65210 379536
rect 67270 564440 67326 564496
rect 66902 477400 66958 477456
rect 66902 476448 66958 476504
rect 66258 442992 66314 443048
rect 66902 382064 66958 382120
rect 67638 578448 67694 578504
rect 68190 577768 68246 577824
rect 67546 577088 67602 577144
rect 67638 575728 67694 575784
rect 67638 574368 67694 574424
rect 67730 573416 67786 573472
rect 67638 573008 67694 573064
rect 67914 571784 67970 571840
rect 68558 580624 68614 580680
rect 68742 576408 68798 576464
rect 68650 571784 68706 571840
rect 67822 571648 67878 571704
rect 68466 571648 68522 571704
rect 67638 570016 67694 570072
rect 67638 568928 67694 568984
rect 67730 568676 67786 568712
rect 67730 568656 67732 568676
rect 67732 568656 67784 568676
rect 67784 568656 67786 568676
rect 67730 567568 67786 567624
rect 67638 567160 67694 567216
rect 67638 565836 67640 565856
rect 67640 565836 67692 565856
rect 67692 565836 67694 565856
rect 67638 565800 67694 565836
rect 67638 564848 67694 564904
rect 67730 563488 67786 563544
rect 67638 563116 67640 563136
rect 67640 563116 67692 563136
rect 67692 563116 67694 563136
rect 67638 563080 67694 563116
rect 67638 562300 67640 562320
rect 67640 562300 67692 562320
rect 67692 562300 67694 562320
rect 67638 562264 67694 562300
rect 67638 562128 67694 562184
rect 67730 560768 67786 560824
rect 67638 560360 67694 560416
rect 67638 559408 67694 559464
rect 68282 557368 68338 557424
rect 67730 556688 67786 556744
rect 67638 556144 67694 556200
rect 67730 555328 67786 555384
rect 67638 554820 67640 554840
rect 67640 554820 67692 554840
rect 67692 554820 67694 554840
rect 67638 554784 67694 554820
rect 67638 553444 67694 553480
rect 67638 553424 67640 553444
rect 67640 553424 67692 553444
rect 67692 553424 67694 553444
rect 67638 552084 67694 552120
rect 67638 552064 67640 552084
rect 67640 552064 67692 552084
rect 67692 552064 67694 552084
rect 67638 551248 67694 551304
rect 67730 549888 67786 549944
rect 67638 549364 67694 549400
rect 67638 549344 67640 549364
rect 67640 549344 67692 549364
rect 67692 549344 67694 549364
rect 67638 547984 67694 548040
rect 67638 546508 67694 546544
rect 67638 546488 67640 546508
rect 67640 546488 67692 546508
rect 67692 546488 67694 546508
rect 67730 543904 67786 543960
rect 68282 543904 68338 543960
rect 68006 543224 68062 543280
rect 67638 542544 67694 542600
rect 67730 541728 67786 541784
rect 67638 541184 67694 541240
rect 67638 540096 67694 540152
rect 67638 487872 67694 487928
rect 67638 487212 67694 487248
rect 67638 487192 67640 487212
rect 67640 487192 67692 487212
rect 67692 487192 67694 487212
rect 67638 486512 67694 486568
rect 68098 485968 68154 486024
rect 67362 480528 67418 480584
rect 67638 485152 67694 485208
rect 67638 482568 67694 482624
rect 67638 481072 67694 481128
rect 67546 479848 67602 479904
rect 67454 478488 67510 478544
rect 67638 476992 67694 477048
rect 67638 475632 67694 475688
rect 67730 475088 67786 475144
rect 67638 474272 67694 474328
rect 67638 473592 67694 473648
rect 67638 472504 67694 472560
rect 67638 471008 67694 471064
rect 67546 470192 67602 470248
rect 67638 469648 67694 469704
rect 67638 468152 67694 468208
rect 67638 466792 67694 466848
rect 67270 466384 67326 466440
rect 67454 466384 67510 466440
rect 67454 465568 67510 465624
rect 67638 466112 67694 466168
rect 67638 464752 67694 464808
rect 67730 464208 67786 464264
rect 67638 462848 67694 462904
rect 67638 462712 67694 462768
rect 67638 461352 67694 461408
rect 67638 460672 67694 460728
rect 67730 460164 67732 460184
rect 67732 460164 67784 460184
rect 67784 460164 67786 460184
rect 67730 460128 67786 460164
rect 67638 459312 67694 459368
rect 67454 371728 67510 371784
rect 67086 345888 67142 345944
rect 67730 457272 67786 457328
rect 67638 456884 67694 456920
rect 67638 456864 67640 456884
rect 67640 456864 67692 456884
rect 67692 456864 67694 456884
rect 67638 455912 67694 455968
rect 67638 454708 67694 454744
rect 67638 454688 67640 454708
rect 67640 454688 67692 454708
rect 67692 454688 67694 454708
rect 67638 453364 67640 453384
rect 67640 453364 67692 453384
rect 67692 453364 67694 453384
rect 67638 453328 67694 453364
rect 67730 453192 67786 453248
rect 67638 449948 67694 449984
rect 67638 449928 67640 449948
rect 67640 449928 67692 449948
rect 67692 449928 67694 449948
rect 67638 449112 67694 449168
rect 67638 447752 67694 447808
rect 67638 446528 67694 446584
rect 67638 445052 67694 445088
rect 67638 445032 67640 445052
rect 67640 445032 67692 445052
rect 67692 445032 67694 445052
rect 68834 558864 68890 558920
rect 68926 550704 68982 550760
rect 68834 544448 68890 544504
rect 68374 484608 68430 484664
rect 68374 479732 68430 479768
rect 68374 479712 68376 479732
rect 68376 479712 68428 479732
rect 68428 479712 68430 479732
rect 68650 477128 68706 477184
rect 67638 443808 67694 443864
rect 68282 443808 68338 443864
rect 67730 442756 67732 442776
rect 67732 442756 67784 442776
rect 67784 442756 67786 442776
rect 67730 442720 67786 442756
rect 67638 441768 67694 441824
rect 67638 441124 67640 441144
rect 67640 441124 67692 441144
rect 67692 441124 67694 441144
rect 67638 441088 67694 441124
rect 67638 440988 67640 441008
rect 67640 440988 67692 441008
rect 67692 440988 67694 441008
rect 67638 440952 67694 440988
rect 69018 543224 69074 543280
rect 75090 583888 75146 583944
rect 81438 583752 81494 583808
rect 81806 583752 81862 583808
rect 88246 584024 88302 584080
rect 88982 583888 89038 583944
rect 91374 583752 91430 583808
rect 101862 582392 101918 582448
rect 100574 581712 100630 581768
rect 106186 572736 106242 572792
rect 69202 545128 69258 545184
rect 69202 485968 69258 486024
rect 69110 482840 69166 482896
rect 68926 451832 68982 451888
rect 68742 445032 68798 445088
rect 68834 401648 68890 401704
rect 68742 386144 68798 386200
rect 68834 384784 68890 384840
rect 68742 383424 68798 383480
rect 67638 382472 67694 382528
rect 67638 380704 67694 380760
rect 67638 379752 67694 379808
rect 68006 379616 68062 379672
rect 67638 378664 67694 378720
rect 67638 377032 67694 377088
rect 67638 375944 67694 376000
rect 67638 374620 67640 374640
rect 67640 374620 67692 374640
rect 67692 374620 67694 374640
rect 67638 374584 67694 374620
rect 67638 373224 67694 373280
rect 67638 372408 67694 372464
rect 67730 370232 67786 370288
rect 67638 369688 67694 369744
rect 67638 369008 67694 369064
rect 67914 367376 67970 367432
rect 68742 367376 68798 367432
rect 67638 366424 67694 366480
rect 68466 365744 68522 365800
rect 67638 363704 67694 363760
rect 67730 363568 67786 363624
rect 67362 353368 67418 353424
rect 67638 362344 67694 362400
rect 67638 361256 67694 361312
rect 67638 360576 67694 360632
rect 67638 359508 67694 359544
rect 68558 364656 68614 364712
rect 67638 359488 67640 359508
rect 67640 359488 67692 359508
rect 67692 359488 67694 359508
rect 67638 358128 67694 358184
rect 67638 357468 67694 357504
rect 67638 357448 67640 357468
rect 67640 357448 67692 357468
rect 67692 357448 67694 357468
rect 67638 356904 67694 356960
rect 67638 355816 67694 355872
rect 67638 354748 67694 354784
rect 67638 354728 67640 354748
rect 67640 354728 67692 354748
rect 67692 354728 67694 354748
rect 68558 352688 68614 352744
rect 67638 352588 67640 352608
rect 67640 352588 67692 352608
rect 67692 352588 67694 352608
rect 67638 352552 67694 352588
rect 68006 351212 68062 351248
rect 68006 351192 68008 351212
rect 68008 351192 68060 351212
rect 68060 351192 68062 351212
rect 67638 349852 67694 349888
rect 67638 349832 67640 349852
rect 67640 349832 67692 349852
rect 67692 349832 67694 349852
rect 67638 349172 67694 349208
rect 67638 349152 67640 349172
rect 67640 349152 67692 349172
rect 67692 349152 67694 349172
rect 67638 348492 67694 348528
rect 67638 348472 67640 348492
rect 67640 348472 67692 348492
rect 67692 348472 67694 348492
rect 67638 347248 67694 347304
rect 67638 345616 67694 345672
rect 67638 344392 67694 344448
rect 68006 344256 68062 344312
rect 67638 342896 67694 342952
rect 67638 341672 67694 341728
rect 68650 341572 68652 341592
rect 68652 341572 68704 341592
rect 68704 341572 68706 341592
rect 68650 341536 68706 341572
rect 68650 340584 68706 340640
rect 105726 543768 105782 543824
rect 69754 489912 69810 489968
rect 80334 538056 80390 538112
rect 80334 537376 80390 537432
rect 86130 498752 86186 498808
rect 92570 531936 92626 531992
rect 90362 497392 90418 497448
rect 86774 496168 86830 496224
rect 89626 496032 89682 496088
rect 87694 490592 87750 490648
rect 97078 536832 97134 536888
rect 95790 493312 95846 493368
rect 95054 490592 95110 490648
rect 97078 490456 97134 490512
rect 69846 489096 69902 489152
rect 99378 443672 99434 443728
rect 69110 436464 69166 436520
rect 70398 436056 70454 436112
rect 71042 438912 71098 438968
rect 69110 374176 69166 374232
rect 67546 323584 67602 323640
rect 67270 312568 67326 312624
rect 65982 295976 66038 296032
rect 67454 291080 67510 291136
rect 66902 289176 66958 289232
rect 68926 351192 68982 351248
rect 75182 438096 75238 438152
rect 77298 434560 77354 434616
rect 74630 387912 74686 387968
rect 78034 387776 78090 387832
rect 84198 438640 84254 438696
rect 84842 438640 84898 438696
rect 84198 437416 84254 437472
rect 85026 437452 85028 437472
rect 85028 437452 85080 437472
rect 85080 437452 85082 437472
rect 85026 437416 85082 437452
rect 83002 392536 83058 392592
rect 86222 386416 86278 386472
rect 94502 400968 94558 401024
rect 97078 437824 97134 437880
rect 99930 442448 99986 442504
rect 99654 438912 99710 438968
rect 96158 389816 96214 389872
rect 100942 537920 100998 537976
rect 101034 446528 101090 446584
rect 100758 441088 100814 441144
rect 100850 440136 100906 440192
rect 101954 480120 102010 480176
rect 101954 451188 101956 451208
rect 101956 451188 102008 451208
rect 102008 451188 102010 451208
rect 101954 451152 102010 451188
rect 103426 488688 103482 488744
rect 102874 488552 102930 488608
rect 103334 488008 103390 488064
rect 103610 487192 103666 487248
rect 103334 486512 103390 486568
rect 103426 486004 103428 486024
rect 103428 486004 103480 486024
rect 103480 486004 103482 486024
rect 103426 485968 103482 486004
rect 102230 485288 102286 485344
rect 102230 484608 102286 484664
rect 102230 483792 102286 483848
rect 102322 482568 102378 482624
rect 102230 482432 102286 482488
rect 102230 481480 102286 481536
rect 102322 481208 102378 481264
rect 102230 479848 102286 479904
rect 102874 477672 102930 477728
rect 102230 476992 102286 477048
rect 102414 477128 102470 477184
rect 102322 476448 102378 476504
rect 102230 475632 102286 475688
rect 102322 475088 102378 475144
rect 102230 474272 102286 474328
rect 102230 472912 102286 472968
rect 102322 472368 102378 472424
rect 102230 471552 102286 471608
rect 103426 474000 103482 474056
rect 102782 470192 102838 470248
rect 102230 469512 102286 469568
rect 102230 466792 102286 466848
rect 102230 466112 102286 466168
rect 102322 465432 102378 465488
rect 102230 462848 102286 462904
rect 102230 462032 102286 462088
rect 102322 461488 102378 461544
rect 102138 460672 102194 460728
rect 102138 459312 102194 459368
rect 102138 458632 102194 458688
rect 102138 456592 102194 456648
rect 102138 454708 102194 454744
rect 102138 454688 102140 454708
rect 102140 454688 102192 454708
rect 102192 454688 102194 454708
rect 102138 453872 102194 453928
rect 102138 451988 102194 452024
rect 102138 451968 102140 451988
rect 102140 451968 102192 451988
rect 102192 451968 102194 451988
rect 102138 449812 102194 449848
rect 102138 449792 102140 449812
rect 102140 449792 102192 449812
rect 102192 449792 102194 449812
rect 102138 447752 102194 447808
rect 102138 445168 102194 445224
rect 102138 443672 102194 443728
rect 102138 442312 102194 442368
rect 102322 460128 102378 460184
rect 102322 457952 102378 458008
rect 102874 454552 102930 454608
rect 103334 454552 103390 454608
rect 102322 453328 102378 453384
rect 102506 450608 102562 450664
rect 102322 449248 102378 449304
rect 102322 447888 102378 447944
rect 102322 445712 102378 445768
rect 102322 443808 102378 443864
rect 103334 391176 103390 391232
rect 103518 468968 103574 469024
rect 103518 464888 103574 464944
rect 103518 456048 103574 456104
rect 104714 464108 104716 464128
rect 104716 464108 104768 464128
rect 104768 464108 104770 464128
rect 104714 464072 104770 464108
rect 103426 389952 103482 390008
rect 101402 388864 101458 388920
rect 104898 481480 104954 481536
rect 104898 480256 104954 480312
rect 105358 450472 105414 450528
rect 105818 540368 105874 540424
rect 106922 584024 106978 584080
rect 106370 574640 106426 574696
rect 106278 560360 106334 560416
rect 108394 579400 108450 579456
rect 109130 581712 109186 581768
rect 108946 580760 109002 580816
rect 108854 580080 108910 580136
rect 108946 578720 109002 578776
rect 108946 578040 109002 578096
rect 108854 577516 108910 577552
rect 108854 577496 108856 577516
rect 108856 577496 108908 577516
rect 108908 577496 108910 577516
rect 108486 576680 108542 576736
rect 108946 576156 109002 576192
rect 108946 576136 108948 576156
rect 108948 576136 109000 576156
rect 109000 576136 109002 576156
rect 108946 573960 109002 574016
rect 107658 573280 107714 573336
rect 108946 571920 109002 571976
rect 107842 571376 107898 571432
rect 107750 557640 107806 557696
rect 107658 556280 107714 556336
rect 107014 551520 107070 551576
rect 106922 542000 106978 542056
rect 106646 462168 106702 462224
rect 106646 460944 106702 461000
rect 105726 447208 105782 447264
rect 108854 570560 108910 570616
rect 108946 570016 109002 570072
rect 108946 569200 109002 569256
rect 108946 567840 109002 567896
rect 108946 567196 108948 567216
rect 108948 567196 109000 567216
rect 109000 567196 109002 567216
rect 108946 567160 109002 567196
rect 108394 566480 108450 566536
rect 108946 565836 108948 565856
rect 108948 565836 109000 565856
rect 109000 565836 109002 565856
rect 108946 565800 109002 565836
rect 108946 565120 109002 565176
rect 108394 563896 108450 563952
rect 108946 562400 109002 562456
rect 108946 561040 109002 561096
rect 108210 560380 108266 560416
rect 108210 560360 108212 560380
rect 108212 560360 108264 560380
rect 108264 560360 108266 560380
rect 108854 559680 108910 559736
rect 108946 559020 109002 559056
rect 108946 559000 108948 559020
rect 108948 559000 109000 559020
rect 109000 559000 109002 559020
rect 108946 558320 109002 558376
rect 108946 556960 109002 557016
rect 108854 555736 108910 555792
rect 108946 554240 109002 554296
rect 108118 552880 108174 552936
rect 107842 552608 107898 552664
rect 107934 546760 107990 546816
rect 107842 540640 107898 540696
rect 108946 550840 109002 550896
rect 108854 550160 108910 550216
rect 108946 549480 109002 549536
rect 108946 548800 109002 548856
rect 108946 547440 109002 547496
rect 108946 546080 109002 546136
rect 108946 545400 109002 545456
rect 108946 543360 109002 543416
rect 108946 539960 109002 540016
rect 108302 471824 108358 471880
rect 108302 471008 108358 471064
rect 106922 395256 106978 395312
rect 106186 388456 106242 388512
rect 108486 465704 108542 465760
rect 108762 388320 108818 388376
rect 111798 583888 111854 583944
rect 111706 544448 111762 544504
rect 111798 494672 111854 494728
rect 113086 479440 113142 479496
rect 113178 442448 113234 442504
rect 112810 387912 112866 387968
rect 74814 385328 74870 385384
rect 114374 487192 114430 487248
rect 114282 389292 114338 389328
rect 114282 389272 114284 389292
rect 114284 389272 114336 389292
rect 114336 389272 114338 389292
rect 115294 385872 115350 385928
rect 115386 378528 115442 378584
rect 115294 377848 115350 377904
rect 69202 352688 69258 352744
rect 115938 451988 115994 452024
rect 115938 451968 115940 451988
rect 115940 451968 115992 451988
rect 115992 451968 115994 451988
rect 116030 383968 116086 384024
rect 115938 370232 115994 370288
rect 115294 344528 115350 344584
rect 71686 339904 71742 339960
rect 71318 338000 71374 338056
rect 71318 337320 71374 337376
rect 70398 333920 70454 333976
rect 70398 333240 70454 333296
rect 69110 311072 69166 311128
rect 68926 298152 68982 298208
rect 67638 291080 67694 291136
rect 67638 288768 67694 288824
rect 67730 288380 67786 288416
rect 67730 288360 67732 288380
rect 67732 288360 67784 288380
rect 67784 288360 67786 288380
rect 68190 288088 68246 288144
rect 69110 287000 69166 287056
rect 68926 286048 68982 286104
rect 67546 285368 67602 285424
rect 67638 284416 67694 284472
rect 68834 283736 68890 283792
rect 67730 283328 67786 283384
rect 67730 280472 67786 280528
rect 67638 280336 67694 280392
rect 67638 279112 67694 279168
rect 67638 277752 67694 277808
rect 68282 277616 68338 277672
rect 67730 276392 67786 276448
rect 67638 276256 67694 276312
rect 67730 275032 67786 275088
rect 67638 274896 67694 274952
rect 67638 273284 67694 273320
rect 67638 273264 67640 273284
rect 67640 273264 67692 273284
rect 67692 273264 67694 273284
rect 67638 272312 67694 272368
rect 68098 272176 68154 272232
rect 67730 271496 67786 271552
rect 67638 271124 67640 271144
rect 67640 271124 67692 271144
rect 67692 271124 67694 271144
rect 67638 271088 67694 271124
rect 67730 269592 67786 269648
rect 67638 269456 67694 269512
rect 67454 268776 67510 268832
rect 67362 245656 67418 245712
rect 67730 268368 67786 268424
rect 67730 266872 67786 266928
rect 67638 266736 67694 266792
rect 67730 265512 67786 265568
rect 67638 265376 67694 265432
rect 67638 264868 67640 264888
rect 67640 264868 67692 264888
rect 67692 264868 67694 264888
rect 67638 264832 67694 264868
rect 67730 262792 67786 262848
rect 67638 262268 67694 262304
rect 67638 262248 67640 262268
rect 67640 262248 67692 262268
rect 67692 262248 67694 262268
rect 67730 261432 67786 261488
rect 67638 260788 67640 260808
rect 67640 260788 67692 260808
rect 67692 260788 67694 260808
rect 67638 260752 67694 260788
rect 67638 259528 67694 259584
rect 67730 258576 67786 258632
rect 67638 258188 67694 258224
rect 67638 258168 67640 258188
rect 67640 258168 67692 258188
rect 67692 258168 67694 258188
rect 67730 257216 67786 257272
rect 67638 256828 67694 256864
rect 67638 256808 67640 256828
rect 67640 256808 67692 256828
rect 67692 256808 67694 256828
rect 67638 255856 67694 255912
rect 67730 255332 67786 255368
rect 67730 255312 67732 255332
rect 67732 255312 67784 255332
rect 67784 255312 67786 255332
rect 67638 255212 67640 255232
rect 67640 255212 67692 255232
rect 67692 255212 67694 255232
rect 67638 255176 67694 255212
rect 67638 254532 67640 254552
rect 67640 254532 67692 254552
rect 67692 254532 67694 254552
rect 67638 254496 67694 254532
rect 68098 252592 68154 252648
rect 67638 251776 67694 251832
rect 67730 250416 67786 250472
rect 67638 249872 67694 249928
rect 67730 249056 67786 249112
rect 67638 248532 67694 248568
rect 67638 248512 67640 248532
rect 67640 248512 67692 248532
rect 67692 248512 67694 248532
rect 67730 247696 67786 247752
rect 67638 247152 67694 247208
rect 67638 244568 67694 244624
rect 67730 243616 67786 243672
rect 67638 243208 67694 243264
rect 68190 241576 68246 241632
rect 67638 240896 67694 240952
rect 69846 296792 69902 296848
rect 73894 339360 73950 339416
rect 73894 338000 73950 338056
rect 74446 338000 74502 338056
rect 73342 335960 73398 336016
rect 71042 292304 71098 292360
rect 75918 339632 75974 339688
rect 77114 339632 77170 339688
rect 75918 312432 75974 312488
rect 75826 294344 75882 294400
rect 77298 299512 77354 299568
rect 78034 337320 78090 337376
rect 80978 330384 81034 330440
rect 79230 302232 79286 302288
rect 77942 294208 77998 294264
rect 79414 293120 79470 293176
rect 80978 296928 81034 296984
rect 88982 309712 89038 309768
rect 89994 295432 90050 295488
rect 94226 307128 94282 307184
rect 95790 294072 95846 294128
rect 104806 339360 104862 339416
rect 104806 338816 104862 338872
rect 107382 339224 107438 339280
rect 107566 339224 107622 339280
rect 113194 339768 113250 339824
rect 108394 301552 108450 301608
rect 111890 292712 111946 292768
rect 114466 295296 114522 295352
rect 117226 485732 117228 485752
rect 117228 485732 117280 485752
rect 117280 485732 117282 485752
rect 117226 485696 117282 485732
rect 116214 383560 116270 383616
rect 116122 369960 116178 370016
rect 117502 397976 117558 398032
rect 117318 387640 117374 387696
rect 117318 376080 117374 376136
rect 117410 363160 117466 363216
rect 117318 357040 117374 357096
rect 118974 454028 119030 454064
rect 118974 454008 118976 454028
rect 118976 454008 119028 454028
rect 119028 454008 119030 454028
rect 119342 454008 119398 454064
rect 120354 438912 120410 438968
rect 117686 384920 117742 384976
rect 118606 384920 118662 384976
rect 118606 382220 118662 382256
rect 118606 382200 118608 382220
rect 118608 382200 118660 382220
rect 118660 382200 118662 382220
rect 118606 381556 118608 381576
rect 118608 381556 118660 381576
rect 118660 381556 118662 381576
rect 118606 381520 118662 381556
rect 118606 380840 118662 380896
rect 118514 379516 118516 379536
rect 118516 379516 118568 379536
rect 118568 379516 118570 379536
rect 118514 379480 118570 379516
rect 118606 378836 118608 378856
rect 118608 378836 118660 378856
rect 118660 378836 118662 378856
rect 118606 378800 118662 378836
rect 117870 378156 117872 378176
rect 117872 378156 117924 378176
rect 117924 378156 117926 378176
rect 117870 378120 117926 378156
rect 118606 376796 118608 376816
rect 118608 376796 118660 376816
rect 118660 376796 118662 376816
rect 118606 376760 118662 376796
rect 118606 375420 118662 375456
rect 118606 375400 118608 375420
rect 118608 375400 118660 375420
rect 118660 375400 118662 375420
rect 118146 374040 118202 374096
rect 118330 373360 118386 373416
rect 118514 372680 118570 372736
rect 118146 371320 118202 371376
rect 118146 369960 118202 370016
rect 118606 368600 118662 368656
rect 118606 367920 118662 367976
rect 118606 367260 118662 367296
rect 118606 367240 118608 367260
rect 118608 367240 118660 367260
rect 118660 367240 118662 367260
rect 118606 365880 118662 365936
rect 118514 365200 118570 365256
rect 118606 364520 118662 364576
rect 117502 355680 117558 355736
rect 117502 354320 117558 354376
rect 117502 352960 117558 353016
rect 118606 362480 118662 362536
rect 118606 361800 118662 361856
rect 118054 361120 118110 361176
rect 118606 359760 118662 359816
rect 117962 359080 118018 359136
rect 118606 358400 118662 358456
rect 118238 357040 118294 357096
rect 118606 356360 118662 356416
rect 118606 353640 118662 353696
rect 117686 351600 117742 351656
rect 118606 351600 118662 351656
rect 118054 350920 118110 350976
rect 117502 350240 117558 350296
rect 117410 348880 117466 348936
rect 118514 348880 118570 348936
rect 117962 348200 118018 348256
rect 118606 347520 118662 347576
rect 118514 346160 118570 346216
rect 117870 344800 117926 344856
rect 118054 342080 118110 342136
rect 116122 340040 116178 340096
rect 117962 340040 118018 340096
rect 118606 345480 118662 345536
rect 118606 343440 118662 343496
rect 118606 342760 118662 342816
rect 118606 340756 118608 340776
rect 118608 340756 118660 340776
rect 118660 340756 118662 340776
rect 118606 340720 118662 340756
rect 115294 292576 115350 292632
rect 115754 292576 115810 292632
rect 118330 298288 118386 298344
rect 119434 375944 119490 376000
rect 119526 368328 119582 368384
rect 119342 360848 119398 360904
rect 118790 355680 118846 355736
rect 119342 338000 119398 338056
rect 119066 292032 119122 292088
rect 117962 291896 118018 291952
rect 69846 290808 69902 290864
rect 69202 282104 69258 282160
rect 68926 263608 68982 263664
rect 68834 239400 68890 239456
rect 67638 234504 67694 234560
rect 69018 253136 69074 253192
rect 69110 251232 69166 251288
rect 120906 284316 120908 284336
rect 120908 284316 120960 284336
rect 120960 284316 120962 284336
rect 120906 284280 120962 284316
rect 121274 257100 121330 257136
rect 121274 257080 121276 257100
rect 121276 257080 121328 257100
rect 121328 257080 121330 257100
rect 120078 250960 120134 251016
rect 69202 244976 69258 245032
rect 69846 242256 69902 242312
rect 70398 216008 70454 216064
rect 68926 199280 68982 199336
rect 74538 185544 74594 185600
rect 76562 237224 76618 237280
rect 76562 220088 76618 220144
rect 77390 208936 77446 208992
rect 86130 237904 86186 237960
rect 87050 215872 87106 215928
rect 84290 192480 84346 192536
rect 91282 234368 91338 234424
rect 95790 235728 95846 235784
rect 78678 182824 78734 182880
rect 98366 238584 98422 238640
rect 98642 235728 98698 235784
rect 103610 222808 103666 222864
rect 97354 176976 97410 177032
rect 107382 235864 107438 235920
rect 106278 212472 106334 212528
rect 104806 177656 104862 177712
rect 106186 177656 106242 177712
rect 108946 177656 109002 177712
rect 100666 176704 100722 176760
rect 102046 176724 102102 176760
rect 102046 176704 102048 176724
rect 102048 176704 102100 176724
rect 102100 176704 102102 176724
rect 103426 176704 103482 176760
rect 113822 237224 113878 237280
rect 113822 236000 113878 236056
rect 114466 236000 114522 236056
rect 114650 219272 114706 219328
rect 119342 206216 119398 206272
rect 121642 439456 121698 439512
rect 123114 576000 123170 576056
rect 122838 490456 122894 490512
rect 122102 439456 122158 439512
rect 121550 388320 121606 388376
rect 122010 329740 122012 329760
rect 122012 329740 122064 329760
rect 122064 329740 122066 329760
rect 122010 329704 122066 329740
rect 123206 483676 123262 483712
rect 123206 483656 123208 483676
rect 123208 483656 123260 483676
rect 123260 483656 123262 483676
rect 121550 291796 121552 291816
rect 121552 291796 121604 291816
rect 121604 291796 121606 291816
rect 121550 291760 121606 291796
rect 121642 291080 121698 291136
rect 121550 290400 121606 290456
rect 121826 295976 121882 296032
rect 121734 289720 121790 289776
rect 121642 289040 121698 289096
rect 121550 287680 121606 287736
rect 121550 287000 121606 287056
rect 121642 286356 121644 286376
rect 121644 286356 121696 286376
rect 121696 286356 121698 286376
rect 121642 286320 121698 286356
rect 121458 285640 121514 285696
rect 121458 284960 121514 285016
rect 121458 282940 121514 282976
rect 121458 282920 121460 282940
rect 121460 282920 121512 282940
rect 121512 282920 121514 282940
rect 121458 281580 121514 281616
rect 121458 281560 121460 281580
rect 121460 281560 121512 281580
rect 121512 281560 121514 281580
rect 121458 280220 121514 280256
rect 121458 280200 121460 280220
rect 121460 280200 121512 280220
rect 121512 280200 121514 280220
rect 121550 279520 121606 279576
rect 121458 278840 121514 278896
rect 121550 278160 121606 278216
rect 121458 277500 121514 277536
rect 121458 277480 121460 277500
rect 121460 277480 121512 277500
rect 121512 277480 121514 277500
rect 121642 276256 121698 276312
rect 121458 276140 121514 276176
rect 121458 276120 121460 276140
rect 121460 276120 121512 276140
rect 121512 276120 121514 276140
rect 121550 275440 121606 275496
rect 121458 274760 121514 274816
rect 121458 273400 121514 273456
rect 121458 272720 121514 272776
rect 121458 272040 121514 272096
rect 121458 271360 121514 271416
rect 121458 270000 121514 270056
rect 121550 269320 121606 269376
rect 121458 268640 121514 268696
rect 121918 275984 121974 276040
rect 123114 378936 123170 378992
rect 122286 288360 122342 288416
rect 122102 274080 122158 274136
rect 121918 272448 121974 272504
rect 121550 267960 121606 268016
rect 121642 267280 121698 267336
rect 121550 266600 121606 266656
rect 121642 265920 121698 265976
rect 121550 265240 121606 265296
rect 121642 263880 121698 263936
rect 126150 572736 126206 572792
rect 125690 484336 125746 484392
rect 121550 263200 121606 263256
rect 121550 262520 121606 262576
rect 121642 261840 121698 261896
rect 121550 261160 121606 261216
rect 121550 260480 121606 260536
rect 121550 259800 121606 259856
rect 121550 258440 121606 258496
rect 121458 257760 121514 257816
rect 121734 259120 121790 259176
rect 121458 256400 121514 256456
rect 121458 254360 121514 254416
rect 121458 253000 121514 253056
rect 121458 251640 121514 251696
rect 121458 250280 121514 250336
rect 121458 248920 121514 248976
rect 121642 255040 121698 255096
rect 121642 253680 121698 253736
rect 122746 255720 122802 255776
rect 121734 252320 121790 252376
rect 121642 249600 121698 249656
rect 121458 248240 121514 248296
rect 121366 247560 121422 247616
rect 121550 246880 121606 246936
rect 121458 246200 121514 246256
rect 121550 245520 121606 245576
rect 121458 244840 121514 244896
rect 121550 244160 121606 244216
rect 121458 242820 121514 242856
rect 121458 242800 121460 242820
rect 121460 242800 121512 242820
rect 121512 242800 121514 242820
rect 121550 242120 121606 242176
rect 122102 243480 122158 243536
rect 121642 241440 121698 241496
rect 121458 240760 121514 240816
rect 122746 240760 122802 240816
rect 122102 240080 122158 240136
rect 124494 379636 124550 379672
rect 124494 379616 124496 379636
rect 124496 379616 124548 379636
rect 124548 379616 124550 379636
rect 127346 496032 127402 496088
rect 125598 328344 125654 328400
rect 124310 301416 124366 301472
rect 124310 264560 124366 264616
rect 124310 262792 124366 262848
rect 126334 295432 126390 295488
rect 127530 386960 127586 387016
rect 129922 553968 129978 554024
rect 128542 445068 128544 445088
rect 128544 445068 128596 445088
rect 128596 445068 128598 445088
rect 128542 445032 128598 445068
rect 129738 493312 129794 493368
rect 130382 537920 130438 537976
rect 130382 461080 130438 461136
rect 128818 335280 128874 335336
rect 129738 292712 129794 292768
rect 130106 342916 130162 342952
rect 130106 342896 130108 342916
rect 130108 342896 130160 342916
rect 130160 342896 130162 342916
rect 132498 391992 132554 392048
rect 131118 293120 131174 293176
rect 132774 468424 132830 468480
rect 132774 400832 132830 400888
rect 132498 282784 132554 282840
rect 133786 282784 133842 282840
rect 133786 282104 133842 282160
rect 134062 353640 134118 353696
rect 136546 388320 136602 388376
rect 138018 460944 138074 461000
rect 137282 336096 137338 336152
rect 141146 490456 141202 490512
rect 141146 387912 141202 387968
rect 364982 701664 365038 701720
rect 140870 234368 140926 234424
rect 139398 212472 139454 212528
rect 139398 211792 139454 211848
rect 133142 198056 133198 198112
rect 112258 176840 112314 176896
rect 109774 176704 109830 176760
rect 116950 177656 117006 177712
rect 115846 177112 115902 177168
rect 119526 177656 119582 177712
rect 122010 177656 122066 177712
rect 120998 177112 121054 177168
rect 143630 219272 143686 219328
rect 143630 218592 143686 218648
rect 146942 291896 146998 291952
rect 149150 451288 149206 451344
rect 147954 298288 148010 298344
rect 149150 334600 149206 334656
rect 151818 480256 151874 480312
rect 152002 468424 152058 468480
rect 147586 188264 147642 188320
rect 336002 405728 336058 405784
rect 166262 400288 166318 400344
rect 153106 370504 153162 370560
rect 155314 197920 155370 197976
rect 162214 292576 162270 292632
rect 129646 177656 129702 177712
rect 131026 177656 131082 177712
rect 132406 177656 132462 177712
rect 133142 177112 133198 177168
rect 110694 176740 110696 176760
rect 110696 176740 110748 176760
rect 110748 176740 110750 176760
rect 110694 176704 110750 176740
rect 114374 176704 114430 176760
rect 118422 176704 118478 176760
rect 124494 176704 124550 176760
rect 125782 176704 125838 176760
rect 127070 176704 127126 176760
rect 134430 176704 134486 176760
rect 148230 176704 148286 176760
rect 109406 175888 109462 175944
rect 98366 175344 98422 175400
rect 135718 175480 135774 175536
rect 128174 175344 128230 175400
rect 158902 175344 158958 175400
rect 113178 174936 113234 174992
rect 123114 174936 123170 174992
rect 166262 178608 166318 178664
rect 169022 237904 169078 237960
rect 167090 171536 167146 171592
rect 66166 129240 66222 129296
rect 66074 128016 66130 128072
rect 65154 126248 65210 126304
rect 65982 102312 66038 102368
rect 66074 94832 66130 94888
rect 67638 125160 67694 125216
rect 67546 123528 67602 123584
rect 67362 122576 67418 122632
rect 66166 93744 66222 93800
rect 67454 120808 67510 120864
rect 67362 91024 67418 91080
rect 67730 100680 67786 100736
rect 93858 94696 93914 94752
rect 106646 94696 106702 94752
rect 118238 94696 118294 94752
rect 120630 94696 120686 94752
rect 114374 93608 114430 93664
rect 113822 93472 113878 93528
rect 103426 93200 103482 93256
rect 110142 93200 110198 93256
rect 129462 93472 129518 93528
rect 74814 92384 74870 92440
rect 84382 92384 84438 92440
rect 88982 92420 88984 92440
rect 88984 92420 89036 92440
rect 89036 92420 89038 92440
rect 88982 92384 89038 92420
rect 98182 92384 98238 92440
rect 100574 91704 100630 91760
rect 102874 91704 102930 91760
rect 97814 91296 97870 91352
rect 99194 91296 99250 91352
rect 85854 91160 85910 91216
rect 86866 91160 86922 91216
rect 88062 91160 88118 91216
rect 90638 91160 90694 91216
rect 92294 91160 92350 91216
rect 93766 91160 93822 91216
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 97906 91160 97962 91216
rect 97814 81368 97870 81424
rect 99286 91160 99342 91216
rect 101954 91432 102010 91488
rect 101862 91296 101918 91352
rect 100666 91160 100722 91216
rect 102046 91160 102102 91216
rect 101954 85448 102010 85504
rect 105910 92384 105966 92440
rect 104714 91296 104770 91352
rect 104806 91160 104862 91216
rect 103426 82728 103482 82784
rect 108946 91296 109002 91352
rect 106094 91160 106150 91216
rect 107198 91160 107254 91216
rect 108854 91160 108910 91216
rect 104806 81232 104862 81288
rect 111614 92384 111670 92440
rect 115846 92384 115902 92440
rect 110326 91296 110382 91352
rect 110234 91160 110290 91216
rect 110786 91160 110842 91216
rect 124586 92384 124642 92440
rect 125966 92384 126022 92440
rect 126518 92384 126574 92440
rect 121090 91840 121146 91896
rect 115846 91568 115902 91624
rect 113086 91296 113142 91352
rect 112994 91160 113050 91216
rect 110786 88168 110842 88224
rect 115754 91160 115810 91216
rect 117134 91296 117190 91352
rect 117226 91160 117282 91216
rect 118238 91160 118294 91216
rect 119986 91160 120042 91216
rect 122746 91296 122802 91352
rect 124034 91296 124090 91352
rect 122654 91160 122710 91216
rect 121090 89664 121146 89720
rect 117226 82592 117282 82648
rect 122838 91160 122894 91216
rect 124126 91160 124182 91216
rect 125414 91160 125470 91216
rect 151726 93608 151782 93664
rect 133142 92384 133198 92440
rect 136086 92384 136142 92440
rect 151542 92384 151598 92440
rect 152094 92384 152150 92440
rect 132406 91568 132462 91624
rect 126886 91160 126942 91216
rect 128174 91160 128230 91216
rect 131026 91160 131082 91216
rect 135074 91160 135130 91216
rect 151634 91160 151690 91216
rect 166538 92248 166594 92304
rect 167918 111732 167920 111752
rect 167920 111732 167972 111752
rect 167972 111732 167974 111752
rect 167918 111696 167974 111732
rect 168102 110064 168158 110120
rect 167918 108704 167974 108760
rect 66718 1944 66774 2000
rect 78678 50224 78734 50280
rect 120078 25472 120134 25528
rect 119894 14456 119950 14512
rect 174634 92112 174690 92168
rect 178682 299512 178738 299568
rect 180062 178608 180118 178664
rect 182914 70216 182970 70272
rect 182178 69536 182234 69592
rect 182914 69536 182970 69592
rect 188434 295296 188490 295352
rect 192574 93744 192630 93800
rect 199474 181328 199530 181384
rect 199474 93744 199530 93800
rect 203614 180104 203670 180160
rect 205086 94832 205142 94888
rect 209134 301416 209190 301472
rect 213182 294344 213238 294400
rect 211802 186904 211858 186960
rect 213274 177248 213330 177304
rect 213918 175752 213974 175808
rect 213918 175072 213974 175128
rect 214010 174664 214066 174720
rect 213918 173712 213974 173768
rect 214010 173304 214066 173360
rect 213918 172352 213974 172408
rect 214102 171944 214158 172000
rect 214010 170856 214066 170912
rect 213918 170720 213974 170776
rect 213918 169652 213974 169688
rect 213918 169632 213920 169652
rect 213920 169632 213972 169652
rect 213972 169632 213974 169652
rect 214010 169360 214066 169416
rect 213918 168292 213974 168328
rect 213918 168272 213920 168292
rect 213920 168272 213972 168292
rect 213972 168272 213974 168292
rect 214010 168000 214066 168056
rect 214102 166932 214158 166968
rect 214102 166912 214104 166932
rect 214104 166912 214156 166932
rect 214156 166912 214158 166932
rect 213918 166096 213974 166152
rect 213918 165280 213974 165336
rect 214010 164736 214066 164792
rect 213918 164092 213920 164112
rect 213920 164092 213972 164112
rect 213972 164092 213974 164112
rect 213918 164056 213974 164092
rect 214010 163376 214066 163432
rect 214654 166640 214710 166696
rect 214562 162696 214618 162752
rect 213918 162016 213974 162072
rect 214746 161200 214802 161256
rect 213918 160012 213920 160032
rect 213920 160012 213972 160032
rect 213972 160012 213974 160032
rect 213918 159976 213974 160012
rect 214010 159432 214066 159488
rect 213918 158652 213920 158672
rect 213920 158652 213972 158672
rect 213972 158652 213974 158672
rect 213918 158616 213974 158652
rect 213366 158072 213422 158128
rect 214010 157936 214066 157992
rect 214010 157256 214066 157312
rect 213918 156848 213974 156904
rect 213918 155896 213974 155952
rect 214010 155488 214066 155544
rect 214010 153856 214066 153912
rect 213918 153448 213974 153504
rect 213918 152632 213974 152688
rect 214010 152224 214066 152280
rect 213918 151952 213974 152008
rect 214010 150592 214066 150648
rect 213918 150048 213974 150104
rect 213918 148688 213974 148744
rect 214654 150728 214710 150784
rect 214562 149504 214618 149560
rect 213918 148008 213974 148064
rect 213918 146648 213974 146704
rect 214102 146376 214158 146432
rect 214010 145288 214066 145344
rect 213918 144880 213974 144936
rect 213918 143928 213974 143984
rect 214010 143520 214066 143576
rect 213274 142704 213330 142760
rect 213182 94968 213238 95024
rect 213918 142180 213974 142216
rect 213918 142160 213920 142180
rect 213920 142160 213972 142180
rect 213972 142160 213974 142180
rect 214010 141344 214066 141400
rect 213918 140936 213974 140992
rect 213918 139984 213974 140040
rect 213918 138760 213974 138816
rect 213366 138080 213422 138136
rect 214562 136720 214618 136776
rect 214010 136040 214066 136096
rect 213918 135380 213974 135416
rect 213918 135360 213920 135380
rect 213920 135360 213972 135380
rect 213972 135360 213974 135380
rect 213918 134000 213974 134056
rect 214010 132776 214066 132832
rect 213918 132524 213974 132560
rect 213918 132504 213920 132524
rect 213920 132504 213972 132524
rect 213972 132504 213974 132524
rect 213918 131416 213974 131472
rect 214010 128832 214066 128888
rect 213918 128444 213974 128480
rect 213918 128424 213920 128444
rect 213920 128424 213972 128444
rect 213972 128424 213974 128444
rect 214010 126112 214066 126168
rect 213918 125704 213974 125760
rect 214010 124752 214066 124808
rect 213918 124344 213974 124400
rect 214010 123528 214066 123584
rect 213918 122868 213974 122904
rect 213918 122848 213920 122868
rect 213920 122848 213972 122868
rect 213972 122848 213974 122868
rect 214010 122168 214066 122224
rect 213918 121760 213974 121816
rect 214010 120808 214066 120864
rect 213918 120148 213974 120184
rect 213918 120128 213920 120148
rect 213920 120128 213972 120148
rect 213972 120128 213974 120148
rect 214010 119584 214066 119640
rect 213918 118904 213974 118960
rect 214102 118804 214104 118824
rect 214104 118804 214156 118824
rect 214156 118804 214158 118824
rect 214102 118768 214158 118804
rect 214010 117544 214066 117600
rect 213918 117272 213974 117328
rect 214010 116184 214066 116240
rect 213918 115912 213974 115968
rect 214010 114960 214066 115016
rect 213918 114588 213920 114608
rect 213920 114588 213972 114608
rect 213972 114588 213974 114608
rect 213918 114552 213974 114588
rect 214010 113600 214066 113656
rect 213918 113228 213920 113248
rect 213920 113228 213972 113248
rect 213972 113228 213974 113248
rect 213918 113192 213974 113228
rect 214010 112240 214066 112296
rect 213918 111868 213920 111888
rect 213920 111868 213972 111888
rect 213972 111868 213974 111888
rect 213918 111832 213974 111868
rect 214010 110880 214066 110936
rect 213918 110492 213974 110528
rect 213918 110472 213920 110492
rect 213920 110472 213972 110492
rect 213972 110472 213974 110492
rect 214010 109656 214066 109712
rect 213918 109248 213974 109304
rect 214010 108296 214066 108352
rect 213918 107888 213974 107944
rect 214010 106936 214066 106992
rect 213918 106528 213974 106584
rect 213458 105712 213514 105768
rect 214010 105304 214066 105360
rect 213918 105032 213974 105088
rect 214010 103944 214066 104000
rect 213918 103672 213974 103728
rect 213918 102584 213974 102640
rect 213918 100816 213974 100872
rect 214010 99728 214066 99784
rect 213918 99476 213974 99512
rect 213918 99456 213920 99476
rect 213920 99456 213972 99476
rect 213972 99456 213974 99476
rect 214010 98368 214066 98424
rect 213918 97996 213920 98016
rect 213920 97996 213972 98016
rect 213972 97996 213974 98016
rect 213918 97960 213974 97996
rect 213918 97008 213974 97064
rect 213918 95784 213974 95840
rect 214654 135496 214710 135552
rect 214746 127472 214802 127528
rect 214838 101088 214894 101144
rect 214562 90344 214618 90400
rect 214930 96600 214986 96656
rect 218702 178608 218758 178664
rect 221554 177792 221610 177848
rect 224314 189624 224370 189680
rect 226982 177384 227038 177440
rect 227074 176296 227130 176352
rect 229098 176296 229154 176352
rect 227718 175788 227720 175808
rect 227720 175788 227772 175808
rect 227772 175788 227774 175808
rect 227718 175752 227774 175788
rect 229098 174256 229154 174312
rect 229190 161472 229246 161528
rect 229558 173712 229614 173768
rect 229466 172760 229522 172816
rect 229374 171808 229430 171864
rect 229282 146784 229338 146840
rect 230478 158616 230534 158672
rect 230110 157392 230166 157448
rect 229926 143384 229982 143440
rect 229742 142432 229798 142488
rect 230478 150592 230534 150648
rect 231398 173304 231454 173360
rect 231766 172372 231822 172408
rect 231766 172352 231768 172372
rect 231768 172352 231820 172372
rect 231820 172352 231822 172372
rect 231674 171400 231730 171456
rect 231674 170892 231676 170912
rect 231676 170892 231728 170912
rect 231728 170892 231730 170912
rect 231674 170856 231730 170892
rect 231766 170448 231822 170504
rect 231766 169904 231822 169960
rect 231766 169532 231768 169552
rect 231768 169532 231820 169552
rect 231820 169532 231822 169552
rect 231766 169496 231822 169532
rect 231674 168952 231730 169008
rect 231398 168544 231454 168600
rect 231766 168000 231822 168056
rect 231214 167048 231270 167104
rect 231766 166640 231822 166696
rect 231490 166096 231546 166152
rect 231582 165688 231638 165744
rect 231030 165144 231086 165200
rect 231122 164328 231178 164384
rect 231766 163784 231822 163840
rect 231674 163376 231730 163432
rect 231490 162832 231546 162888
rect 231950 162424 232006 162480
rect 231766 161880 231822 161936
rect 231306 160928 231362 160984
rect 231766 160520 231822 160576
rect 231582 159976 231638 160032
rect 231030 159568 231086 159624
rect 231766 159024 231822 159080
rect 231214 158072 231270 158128
rect 231766 157664 231822 157720
rect 231766 157120 231822 157176
rect 231122 156712 231178 156768
rect 230938 156168 230994 156224
rect 231490 154808 231546 154864
rect 230754 147736 230810 147792
rect 230846 145832 230902 145888
rect 230662 140664 230718 140720
rect 230110 137808 230166 137864
rect 230754 135360 230810 135416
rect 230570 134000 230626 134056
rect 230662 132096 230718 132152
rect 232042 155760 232098 155816
rect 231766 155216 231822 155272
rect 231766 154264 231822 154320
rect 231674 153856 231730 153912
rect 231766 152904 231822 152960
rect 231582 151952 231638 152008
rect 231766 151544 231822 151600
rect 231674 151000 231730 151056
rect 231766 149640 231822 149696
rect 231674 149096 231730 149152
rect 231306 148144 231362 148200
rect 231766 146240 231822 146296
rect 231398 145288 231454 145344
rect 231766 144336 231822 144392
rect 231766 143964 231768 143984
rect 231768 143964 231820 143984
rect 231820 143964 231822 143984
rect 231766 143928 231822 143964
rect 231766 142976 231822 143032
rect 231766 141616 231822 141672
rect 231490 141072 231546 141128
rect 231306 139748 231308 139768
rect 231308 139748 231360 139768
rect 231360 139748 231362 139768
rect 231306 139712 231362 139748
rect 231306 139168 231362 139224
rect 231766 138760 231822 138816
rect 231490 138252 231492 138272
rect 231492 138252 231544 138272
rect 231544 138252 231546 138272
rect 231490 138216 231546 138252
rect 231398 137264 231454 137320
rect 231398 135904 231454 135960
rect 231766 136856 231822 136912
rect 231766 134952 231822 135008
rect 231674 134408 231730 134464
rect 231766 133456 231822 133512
rect 231674 133048 231730 133104
rect 231582 132504 231638 132560
rect 231674 131552 231730 131608
rect 231766 131144 231822 131200
rect 231766 130600 231822 130656
rect 231398 130192 231454 130248
rect 231306 129784 231362 129840
rect 231398 128832 231454 128888
rect 231214 127336 231270 127392
rect 231122 125976 231178 126032
rect 231306 125024 231362 125080
rect 231766 129240 231822 129296
rect 231766 128288 231822 128344
rect 231674 127880 231730 127936
rect 231766 126928 231822 126984
rect 231674 126384 231730 126440
rect 231582 125432 231638 125488
rect 231766 124752 231822 124808
rect 231674 124480 231730 124536
rect 231306 123528 231362 123584
rect 231122 120672 231178 120728
rect 231490 123120 231546 123176
rect 231582 122612 231584 122632
rect 231584 122612 231636 122632
rect 231636 122612 231638 122632
rect 231582 122576 231638 122612
rect 231490 121624 231546 121680
rect 231490 120264 231546 120320
rect 231306 119720 231362 119776
rect 231122 117952 231178 118008
rect 230662 115504 230718 115560
rect 230570 114552 230626 114608
rect 231122 114144 231178 114200
rect 230570 113192 230626 113248
rect 230662 109384 230718 109440
rect 230570 107888 230626 107944
rect 231214 112240 231270 112296
rect 231122 103264 231178 103320
rect 230570 102720 230626 102776
rect 230018 98912 230074 98968
rect 230478 97960 230534 98016
rect 230938 97552 230994 97608
rect 230478 97008 230534 97064
rect 230570 95648 230626 95704
rect 231398 119312 231454 119368
rect 231490 117408 231546 117464
rect 231490 116456 231546 116512
rect 231766 124072 231822 124128
rect 231766 122168 231822 122224
rect 231766 121216 231822 121272
rect 231766 118904 231822 118960
rect 231766 118360 231822 118416
rect 231674 116048 231730 116104
rect 231674 115096 231730 115152
rect 231766 113600 231822 113656
rect 231766 112648 231822 112704
rect 231766 111288 231822 111344
rect 231490 110744 231546 110800
rect 231766 110372 231768 110392
rect 231768 110372 231820 110392
rect 231820 110372 231822 110392
rect 231766 110336 231822 110372
rect 231766 109792 231822 109848
rect 231766 108840 231822 108896
rect 231674 108432 231730 108488
rect 231766 107480 231822 107536
rect 231674 107072 231730 107128
rect 231766 106528 231822 106584
rect 231766 106120 231822 106176
rect 231674 105168 231730 105224
rect 231674 104660 231676 104680
rect 231676 104660 231728 104680
rect 231728 104660 231730 104680
rect 231674 104624 231730 104660
rect 231766 104216 231822 104272
rect 231490 103672 231546 103728
rect 231490 101768 231546 101824
rect 231582 101360 231638 101416
rect 231766 100816 231822 100872
rect 231674 100408 231730 100464
rect 231398 99864 231454 99920
rect 231766 99456 231822 99512
rect 231306 98504 231362 98560
rect 231766 96600 231822 96656
rect 238758 168272 238814 168328
rect 237378 154536 237434 154592
rect 240414 43580 240470 43616
rect 240414 43560 240416 43580
rect 240416 43560 240468 43580
rect 240468 43560 240470 43580
rect 241886 35164 241888 35184
rect 241888 35164 241940 35184
rect 241940 35164 241942 35184
rect 241886 35128 241942 35164
rect 241334 11736 241390 11792
rect 240506 3440 240562 3496
rect 241334 3440 241390 3496
rect 241702 3440 241758 3496
rect 244278 46300 244334 46336
rect 244278 46280 244280 46300
rect 244280 46280 244332 46300
rect 244332 46280 244334 46300
rect 245750 22652 245752 22672
rect 245752 22652 245804 22672
rect 245804 22652 245806 22672
rect 245750 22616 245806 22652
rect 242806 11736 242862 11792
rect 242806 3440 242862 3496
rect 245106 11736 245162 11792
rect 248510 48320 248566 48376
rect 248510 37884 248512 37904
rect 248512 37884 248564 37904
rect 248564 37884 248566 37904
rect 248510 37848 248566 37884
rect 246946 11736 247002 11792
rect 249706 15544 249762 15600
rect 246394 3440 246450 3496
rect 246946 3440 247002 3496
rect 247590 3440 247646 3496
rect 248786 3440 248842 3496
rect 249706 3440 249762 3496
rect 253110 142704 253166 142760
rect 252926 24268 252982 24304
rect 252926 24248 252928 24268
rect 252928 24248 252980 24268
rect 252980 24248 252982 24268
rect 255318 39364 255374 39400
rect 255318 39344 255320 39364
rect 255320 39344 255372 39364
rect 255372 39344 255374 39364
rect 253846 11736 253902 11792
rect 251270 8220 251326 8256
rect 251270 8200 251272 8220
rect 251272 8200 251324 8220
rect 251324 8200 251326 8220
rect 260102 177248 260158 177304
rect 256330 11736 256386 11792
rect 258446 10940 258502 10976
rect 258446 10920 258448 10940
rect 258448 10920 258500 10940
rect 258500 10920 258502 10940
rect 260378 146376 260434 146432
rect 258262 3440 258318 3496
rect 259366 3440 259422 3496
rect 260930 136584 260986 136640
rect 261114 136176 261170 136232
rect 261390 97824 261446 97880
rect 261850 146104 261906 146160
rect 264426 175344 264482 175400
rect 263046 164872 263102 164928
rect 262954 137400 263010 137456
rect 264242 165008 264298 165064
rect 264334 145288 264390 145344
rect 263138 122576 263194 122632
rect 264242 121216 264298 121272
rect 265898 174936 265954 174992
rect 265346 174120 265402 174176
rect 265806 173984 265862 174040
rect 265990 174528 266046 174584
rect 265254 173168 265310 173224
rect 265346 172760 265402 172816
rect 265806 172488 265862 172544
rect 265070 171944 265126 172000
rect 265162 171536 265218 171592
rect 265346 171128 265402 171184
rect 265254 170176 265310 170232
rect 265438 170584 265494 170640
rect 265622 169788 265678 169824
rect 265622 169768 265624 169788
rect 265624 169768 265676 169788
rect 265676 169768 265678 169788
rect 265898 169360 265954 169416
rect 265438 168952 265494 169008
rect 265346 168544 265402 168600
rect 265254 167592 265310 167648
rect 265162 167048 265218 167104
rect 265806 168408 265862 168464
rect 265530 167184 265586 167240
rect 265622 166368 265678 166424
rect 265898 165960 265954 166016
rect 265806 165724 265808 165744
rect 265808 165724 265860 165744
rect 265860 165724 265862 165744
rect 265806 165688 265862 165724
rect 265990 163784 266046 163840
rect 265622 163376 265678 163432
rect 265530 162968 265586 163024
rect 265438 162832 265494 162888
rect 264518 161200 264574 161256
rect 265346 160792 265402 160848
rect 265162 157392 265218 157448
rect 265714 162016 265770 162072
rect 265806 161608 265862 161664
rect 265622 160384 265678 160440
rect 265806 160132 265862 160168
rect 265806 160112 265808 160132
rect 265808 160112 265860 160132
rect 265860 160112 265862 160132
rect 265898 159432 265954 159488
rect 265806 159024 265862 159080
rect 265714 158772 265770 158808
rect 265714 158752 265716 158772
rect 265716 158752 265768 158772
rect 265768 158752 265770 158772
rect 265714 158208 265770 158264
rect 265622 157800 265678 157856
rect 265530 156848 265586 156904
rect 265898 156440 265954 156496
rect 265990 156032 266046 156088
rect 265530 155624 265586 155680
rect 265254 149640 265310 149696
rect 265438 148280 265494 148336
rect 265070 147872 265126 147928
rect 265070 146920 265126 146976
rect 265438 146512 265494 146568
rect 264426 141480 264482 141536
rect 264426 138216 264482 138272
rect 264426 137808 264482 137864
rect 264426 135904 264482 135960
rect 264426 128152 264482 128208
rect 264426 126792 264482 126848
rect 264426 124616 264482 124672
rect 264242 112104 264298 112160
rect 264334 110880 264390 110936
rect 264610 140528 264666 140584
rect 265254 139712 265310 139768
rect 265806 155216 265862 155272
rect 265990 154672 266046 154728
rect 265714 154536 265770 154592
rect 265898 153856 265954 153912
rect 265806 153448 265862 153504
rect 265806 153176 265862 153232
rect 266082 152632 266138 152688
rect 265806 152360 265862 152416
rect 265990 152088 266046 152144
rect 265806 151836 265862 151872
rect 265806 151816 265808 151836
rect 265808 151816 265860 151836
rect 265860 151816 265862 151836
rect 265898 151272 265954 151328
rect 265806 150864 265862 150920
rect 265898 150048 265954 150104
rect 265806 149096 265862 149152
rect 265714 148688 265770 148744
rect 265714 147056 265770 147112
rect 265898 145696 265954 145752
rect 265806 144880 265862 144936
rect 265530 144472 265586 144528
rect 265714 143928 265770 143984
rect 266174 146648 266230 146704
rect 265806 143556 265808 143576
rect 265808 143556 265860 143576
rect 265860 143556 265862 143576
rect 265806 143520 265862 143556
rect 266082 143112 266138 143168
rect 265530 142704 265586 142760
rect 265622 142296 265678 142352
rect 265714 142160 265770 142216
rect 265806 140936 265862 140992
rect 265898 140120 265954 140176
rect 265438 138760 265494 138816
rect 265162 138352 265218 138408
rect 265530 133864 265586 133920
rect 265438 131180 265440 131200
rect 265440 131180 265492 131200
rect 265492 131180 265494 131200
rect 265438 131144 265494 131180
rect 265254 130192 265310 130248
rect 265806 135360 265862 135416
rect 265806 134544 265862 134600
rect 265714 134136 265770 134192
rect 265898 133184 265954 133240
rect 266082 136992 266138 137048
rect 265714 132776 265770 132832
rect 265806 132504 265862 132560
rect 265714 131552 265770 131608
rect 265714 128560 265770 128616
rect 265622 120808 265678 120864
rect 265530 120400 265586 120456
rect 265714 120164 265716 120184
rect 265716 120164 265768 120184
rect 265768 120164 265770 120184
rect 265714 120128 265770 120164
rect 265622 119448 265678 119504
rect 265714 118788 265770 118824
rect 265714 118768 265716 118788
rect 265716 118768 265768 118788
rect 265768 118768 265770 118788
rect 265346 117816 265402 117872
rect 265714 117428 265770 117464
rect 265714 117408 265716 117428
rect 265716 117408 265768 117428
rect 265768 117408 265770 117428
rect 265622 117272 265678 117328
rect 265254 115232 265310 115288
rect 265254 113872 265310 113928
rect 265162 109656 265218 109712
rect 265530 109248 265586 109304
rect 265162 108704 265218 108760
rect 265530 106664 265586 106720
rect 265530 105712 265586 105768
rect 264518 104488 264574 104544
rect 265162 102720 265218 102776
rect 264610 101904 264666 101960
rect 265346 101360 265402 101416
rect 265530 100816 265586 100872
rect 265530 99492 265532 99512
rect 265532 99492 265584 99512
rect 265584 99492 265586 99512
rect 265530 99456 265586 99492
rect 265714 116048 265770 116104
rect 265714 114688 265770 114744
rect 265714 113464 265770 113520
rect 265714 113212 265770 113248
rect 265714 113192 265716 113212
rect 265716 113192 265768 113212
rect 265768 113192 265770 113212
rect 265714 111852 265770 111888
rect 265714 111832 265716 111852
rect 265716 111832 265768 111852
rect 265768 111832 265770 111852
rect 265714 110492 265770 110528
rect 265714 110472 265716 110492
rect 265716 110472 265768 110492
rect 265768 110472 265770 110492
rect 265714 110064 265770 110120
rect 265714 107908 265770 107944
rect 265714 107888 265716 107908
rect 265716 107888 265768 107908
rect 265768 107888 265770 107908
rect 265714 107616 265770 107672
rect 265714 106528 265770 106584
rect 265714 105304 265770 105360
rect 265714 103944 265770 104000
rect 265714 102312 265770 102368
rect 265714 100952 265770 101008
rect 265714 100136 265770 100192
rect 265622 98368 265678 98424
rect 264610 98232 264666 98288
rect 264610 97416 264666 97472
rect 265622 97008 265678 97064
rect 265530 95648 265586 95704
rect 265898 131960 265954 132016
rect 265898 127200 265954 127256
rect 265898 125976 265954 126032
rect 265898 124228 265954 124264
rect 265898 124208 265900 124228
rect 265900 124208 265952 124228
rect 265952 124208 265954 124228
rect 265990 123800 266046 123856
rect 265898 123392 265954 123448
rect 265898 122984 265954 123040
rect 265990 122032 266046 122088
rect 265898 121624 265954 121680
rect 265990 118224 266046 118280
rect 266082 116864 266138 116920
rect 265990 116456 266046 116512
rect 265990 114824 266046 114880
rect 265990 111288 266046 111344
rect 265990 108296 266046 108352
rect 265990 104932 265992 104952
rect 265992 104932 266044 104952
rect 266044 104932 266046 104952
rect 265990 104896 266046 104932
rect 265990 104080 266046 104136
rect 266082 103128 266138 103184
rect 265990 99728 266046 99784
rect 266082 98776 266138 98832
rect 264978 3848 265034 3904
rect 269946 178608 270002 178664
rect 276662 177384 276718 177440
rect 278318 175752 278374 175808
rect 279330 175752 279386 175808
rect 279514 175752 279570 175808
rect 279422 175208 279478 175264
rect 279330 174392 279386 174448
rect 282918 298152 282974 298208
rect 281630 196560 281686 196616
rect 281538 172352 281594 172408
rect 281630 168544 281686 168600
rect 280342 156304 280398 156360
rect 281538 152360 281594 152416
rect 280250 147736 280306 147792
rect 280158 136312 280214 136368
rect 281630 130872 281686 130928
rect 281630 130056 281686 130112
rect 281630 127744 281686 127800
rect 267278 125024 267334 125080
rect 281630 120128 281686 120184
rect 281630 114008 281686 114064
rect 280250 113192 280306 113248
rect 280158 108568 280214 108624
rect 279330 96600 279386 96656
rect 279330 95104 279386 95160
rect 281538 107752 281594 107808
rect 280342 104760 280398 104816
rect 281538 102448 281594 102504
rect 282826 170856 282882 170912
rect 282734 170040 282790 170096
rect 281906 169360 281962 169416
rect 281906 167728 281962 167784
rect 282366 167048 282422 167104
rect 282090 166232 282146 166288
rect 282366 165416 282422 165472
rect 282090 164736 282146 164792
rect 282826 163920 282882 163976
rect 282182 163104 282238 163160
rect 282090 162424 282146 162480
rect 282826 161608 282882 161664
rect 282826 160792 282882 160848
rect 282734 160112 282790 160168
rect 282090 159296 282146 159352
rect 282826 158480 282882 158536
rect 282734 157800 282790 157856
rect 282090 156984 282146 157040
rect 282090 155488 282146 155544
rect 282366 154672 282422 154728
rect 281906 153992 281962 154048
rect 282458 153176 282514 153232
rect 281906 151716 281908 151736
rect 281908 151716 281960 151736
rect 281960 151716 281962 151736
rect 281906 151680 281962 151716
rect 282274 150864 282330 150920
rect 282826 150048 282882 150104
rect 282734 149368 282790 149424
rect 282826 148552 282882 148608
rect 282826 147056 282882 147112
rect 282826 146260 282882 146296
rect 282826 146240 282828 146260
rect 282828 146240 282880 146260
rect 282880 146240 282882 146260
rect 282734 145424 282790 145480
rect 282826 144780 282828 144800
rect 282828 144780 282880 144800
rect 282880 144780 282882 144800
rect 282826 144744 282882 144780
rect 282734 143928 282790 143984
rect 282090 143112 282146 143168
rect 282826 142468 282828 142488
rect 282828 142468 282880 142488
rect 282880 142468 282882 142488
rect 282826 142432 282882 142468
rect 282826 141616 282882 141672
rect 282734 140800 282790 140856
rect 282826 140120 282882 140176
rect 282826 139324 282882 139360
rect 282826 139304 282828 139324
rect 282828 139304 282880 139324
rect 282880 139304 282882 139324
rect 282734 138488 282790 138544
rect 282826 137808 282882 137864
rect 282274 136992 282330 137048
rect 282366 135496 282422 135552
rect 282826 134680 282882 134736
rect 282734 134000 282790 134056
rect 281998 133184 282054 133240
rect 282274 132368 282330 132424
rect 282826 131688 282882 131744
rect 282826 128560 282882 128616
rect 282274 127064 282330 127120
rect 282826 126248 282882 126304
rect 282826 125432 282882 125488
rect 282182 123120 282238 123176
rect 282826 121624 282882 121680
rect 281906 120808 281962 120864
rect 282090 119312 282146 119368
rect 282826 118496 282882 118552
rect 282458 117816 282514 117872
rect 282550 116320 282606 116376
rect 282826 115504 282882 115560
rect 282550 114688 282606 114744
rect 282090 112376 282146 112432
rect 282826 110880 282882 110936
rect 282274 109384 282330 109440
rect 282826 107072 282882 107128
rect 283010 122440 283066 122496
rect 281998 103944 282054 104000
rect 282826 101632 282882 101688
rect 281722 100816 281778 100872
rect 281722 100136 281778 100192
rect 281906 97824 281962 97880
rect 293222 306992 293278 307048
rect 286598 3984 286654 4040
rect 298098 86944 298154 87000
rect 299662 66852 299664 66872
rect 299664 66852 299716 66872
rect 299716 66852 299718 66872
rect 299662 66816 299718 66852
rect 294142 31068 294198 31104
rect 294142 31048 294144 31068
rect 294144 31048 294196 31068
rect 294196 31048 294198 31068
rect 296074 3440 296130 3496
rect 300766 3440 300822 3496
rect 306746 8200 306802 8256
rect 305550 3440 305606 3496
rect 309230 49036 309232 49056
rect 309232 49036 309284 49056
rect 309284 49036 309286 49056
rect 309230 49000 309286 49036
rect 316774 338680 316830 338736
rect 310242 11736 310298 11792
rect 331954 93744 332010 93800
rect 332598 68856 332654 68912
rect 333242 68856 333298 68912
rect 338118 401648 338174 401704
rect 336278 202136 336334 202192
rect 338302 134408 338358 134464
rect 338302 134000 338358 134056
rect 349802 381792 349858 381848
rect 344282 188264 344338 188320
rect 344926 139984 344982 140040
rect 346306 145832 346362 145888
rect 346582 352552 346638 352608
rect 347042 169632 347098 169688
rect 346858 166268 346860 166288
rect 346860 166268 346912 166288
rect 346912 166268 346914 166288
rect 346858 166232 346914 166268
rect 346674 162832 346730 162888
rect 347042 156068 347044 156088
rect 347044 156068 347096 156088
rect 347096 156068 347098 156088
rect 347042 156032 347098 156068
rect 346674 154400 346730 154456
rect 346582 152632 346638 152688
rect 346674 151000 346730 151056
rect 346674 147600 346730 147656
rect 346490 145832 346546 145888
rect 346674 144200 346730 144256
rect 346582 142568 346638 142624
rect 346490 140800 346546 140856
rect 347134 139168 347190 139224
rect 346674 137400 346730 137456
rect 347042 118768 347098 118824
rect 347502 174664 347558 174720
rect 347502 173032 347558 173088
rect 347502 171264 347558 171320
rect 347502 167864 347558 167920
rect 347502 164464 347558 164520
rect 347502 161064 347558 161120
rect 347502 159432 347558 159488
rect 347502 157800 347558 157856
rect 347502 149232 347558 149288
rect 347502 135768 347558 135824
rect 347410 132368 347466 132424
rect 347686 128424 347742 128480
rect 347962 127336 348018 127392
rect 347686 125568 347742 125624
rect 347318 117136 347374 117192
rect 347502 115368 347558 115424
rect 347042 110372 347044 110392
rect 347044 110372 347096 110392
rect 347096 110372 347098 110392
rect 347042 110336 347098 110372
rect 347502 108704 347558 108760
rect 347502 106936 347558 106992
rect 347042 103536 347098 103592
rect 347226 101904 347282 101960
rect 347502 100136 347558 100192
rect 347502 96872 347558 96928
rect 348882 127336 348938 127392
rect 348974 123936 349030 123992
rect 349158 131008 349214 131064
rect 349158 130600 349214 130656
rect 349066 122712 349122 122768
rect 343638 47504 343694 47560
rect 359462 226888 359518 226944
rect 376758 234504 376814 234560
rect 377402 234504 377458 234560
rect 397458 702480 397514 702536
rect 394698 190984 394754 191040
rect 425702 176024 425758 176080
rect 427818 175228 427874 175264
rect 427818 175208 427820 175228
rect 427820 175208 427872 175228
rect 427872 175208 427874 175228
rect 427910 166912 427966 166968
rect 349986 128424 350042 128480
rect 388442 90344 388498 90400
rect 390650 93744 390706 93800
rect 427634 95920 427690 95976
rect 428002 165688 428058 165744
rect 430762 231104 430818 231160
rect 429198 173304 429254 173360
rect 429106 166096 429162 166152
rect 428462 133728 428518 133784
rect 428094 126248 428150 126304
rect 428094 99320 428150 99376
rect 428186 98232 428242 98288
rect 429382 172216 429438 172272
rect 429382 171128 429438 171184
rect 429290 168816 429346 168872
rect 429290 167728 429346 167784
rect 429382 140800 429438 140856
rect 430578 173168 430634 173224
rect 430670 169904 430726 169960
rect 430670 165008 430726 165064
rect 430578 163920 430634 163976
rect 430578 162424 430634 162480
rect 430578 161880 430634 161936
rect 430578 160928 430634 160984
rect 430578 159704 430634 159760
rect 430578 158480 430634 158536
rect 430578 157120 430634 157176
rect 430578 155624 430634 155680
rect 430578 154128 430634 154184
rect 430578 152768 430634 152824
rect 430578 151544 430634 151600
rect 430578 150048 430634 150104
rect 430578 148552 430634 148608
rect 430578 145968 430634 146024
rect 430578 144472 430634 144528
rect 430578 142180 430634 142216
rect 430578 142160 430580 142180
rect 430580 142160 430632 142180
rect 430632 142160 430634 142180
rect 430578 140528 430634 140584
rect 429474 138896 429530 138952
rect 429750 138896 429806 138952
rect 430578 137672 430634 137728
rect 430578 136312 430634 136368
rect 430578 134952 430634 135008
rect 430578 133728 430634 133784
rect 430578 132096 430634 132152
rect 430578 129376 430634 129432
rect 430578 125024 430634 125080
rect 430578 123800 430634 123856
rect 430578 122576 430634 122632
rect 430578 121388 430580 121408
rect 430580 121388 430632 121408
rect 430632 121388 430634 121408
rect 430578 121352 430634 121388
rect 430578 120536 430634 120592
rect 430578 119448 430634 119504
rect 430578 118088 430634 118144
rect 430578 117000 430634 117056
rect 430578 115776 430634 115832
rect 430578 114144 430634 114200
rect 430578 111424 430634 111480
rect 430578 108996 430634 109032
rect 430578 108976 430580 108996
rect 430580 108976 430632 108996
rect 430632 108976 430634 108996
rect 430578 107072 430634 107128
rect 430578 105848 430634 105904
rect 430578 104624 430634 104680
rect 430578 103436 430580 103456
rect 430580 103436 430632 103456
rect 430632 103436 430634 103456
rect 430578 103400 430634 103436
rect 430578 101496 430634 101552
rect 430578 97824 430634 97880
rect 430854 155352 430910 155408
rect 430854 149776 430910 149832
rect 430854 144064 430910 144120
rect 430854 137400 430910 137456
rect 430854 131824 430910 131880
rect 430854 113872 430910 113928
rect 430762 112648 430818 112704
rect 431866 110336 431922 110392
rect 432050 169904 432106 169960
rect 430762 102720 430818 102776
rect 432142 147464 432198 147520
rect 440422 175888 440478 175944
rect 580262 697176 580318 697232
rect 579618 683848 579674 683904
rect 579986 670692 579988 670712
rect 579988 670692 580040 670712
rect 580040 670692 580042 670712
rect 579986 670656 580042 670692
rect 580170 630808 580226 630864
rect 580354 644000 580410 644056
rect 580354 620200 580410 620256
rect 580354 617480 580410 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 579802 524456 579858 524512
rect 580170 511264 580226 511320
rect 580906 491272 580962 491328
rect 580906 484608 580962 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580906 431568 580962 431624
rect 580262 428440 580318 428496
rect 580262 418240 580318 418296
rect 579618 404912 579674 404968
rect 580262 378392 580318 378448
rect 579802 365064 579858 365120
rect 579618 351872 579674 351928
rect 580262 325216 580318 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580262 272176 580318 272232
rect 580170 258848 580226 258904
rect 579986 245520 580042 245576
rect 580170 232328 580226 232384
rect 580170 219000 580226 219056
rect 580170 205672 580226 205728
rect 580906 192480 580962 192536
rect 580262 188264 580318 188320
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 582378 152632 582434 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580354 112784 580410 112840
rect 580262 59608 580318 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect 115054 702476 115060 702540
rect 115124 702538 115130 702540
rect 397453 702538 397519 702541
rect 115124 702536 397519 702538
rect 115124 702480 397458 702536
rect 397514 702480 397519 702536
rect 115124 702478 397519 702480
rect 115124 702476 115130 702478
rect 397453 702475 397519 702478
rect 364977 701722 365043 701725
rect 436134 701722 436140 701724
rect 364977 701720 436140 701722
rect 364977 701664 364982 701720
rect 365038 701664 436140 701720
rect 364977 701662 436140 701664
rect 364977 701659 365043 701662
rect 436134 701660 436140 701662
rect 436204 701660 436210 701724
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 579613 683906 579679 683909
rect 583520 683906 584960 683996
rect 579613 683904 584960 683906
rect 579613 683848 579618 683904
rect 579674 683848 584960 683904
rect 579613 683846 584960 683848
rect 579613 683843 579679 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 579981 670714 580047 670717
rect 583520 670714 584960 670804
rect 579981 670712 584960 670714
rect 579981 670656 579986 670712
rect 580042 670656 584960 670712
rect 579981 670654 584960 670656
rect 579981 670651 580047 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580349 644058 580415 644061
rect 583520 644058 584960 644148
rect 580349 644056 584960 644058
rect 580349 644000 580354 644056
rect 580410 644000 584960 644056
rect 580349 643998 584960 644000
rect 580349 643995 580415 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 111558 620196 111564 620260
rect 111628 620258 111634 620260
rect 580349 620258 580415 620261
rect 111628 620256 580415 620258
rect 111628 620200 580354 620256
rect 580410 620200 580415 620256
rect 111628 620198 580415 620200
rect 111628 620196 111634 620198
rect 580349 620195 580415 620198
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580349 617538 580415 617541
rect 583520 617538 584960 617628
rect 580349 617536 584960 617538
rect 580349 617480 580354 617536
rect 580410 617480 584960 617536
rect 580349 617478 584960 617480
rect 580349 617475 580415 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect 88241 584082 88307 584085
rect 106917 584082 106983 584085
rect 88241 584080 106983 584082
rect 88241 584024 88246 584080
rect 88302 584024 106922 584080
rect 106978 584024 106983 584080
rect 88241 584022 106983 584024
rect 88241 584019 88307 584022
rect 106917 584019 106983 584022
rect 50889 583946 50955 583949
rect 75085 583946 75151 583949
rect 50889 583944 75151 583946
rect 50889 583888 50894 583944
rect 50950 583888 75090 583944
rect 75146 583888 75151 583944
rect 50889 583886 75151 583888
rect 50889 583883 50955 583886
rect 75085 583883 75151 583886
rect 88977 583946 89043 583949
rect 111793 583946 111859 583949
rect 88977 583944 111859 583946
rect 88977 583888 88982 583944
rect 89038 583888 111798 583944
rect 111854 583888 111859 583944
rect 88977 583886 111859 583888
rect 88977 583883 89043 583886
rect 111793 583883 111859 583886
rect 57697 583810 57763 583813
rect 81433 583810 81499 583813
rect 81801 583810 81867 583813
rect 57697 583808 81867 583810
rect 57697 583752 57702 583808
rect 57758 583752 81438 583808
rect 81494 583752 81806 583808
rect 81862 583752 81867 583808
rect 57697 583750 81867 583752
rect 57697 583747 57763 583750
rect 81433 583747 81499 583750
rect 81801 583747 81867 583750
rect 91369 583810 91435 583813
rect 124254 583810 124260 583812
rect 91369 583808 124260 583810
rect 91369 583752 91374 583808
rect 91430 583752 124260 583808
rect 91369 583750 124260 583752
rect 91369 583747 91435 583750
rect 124254 583748 124260 583750
rect 124324 583748 124330 583812
rect 101857 582450 101923 582453
rect 118734 582450 118740 582452
rect 101857 582448 118740 582450
rect 101857 582392 101862 582448
rect 101918 582392 118740 582448
rect 101857 582390 118740 582392
rect 101857 582387 101923 582390
rect 118734 582388 118740 582390
rect 118804 582388 118810 582452
rect 100569 581770 100635 581773
rect 109125 581770 109191 581773
rect 100569 581768 109191 581770
rect 100569 581712 100574 581768
rect 100630 581712 109130 581768
rect 109186 581712 109191 581768
rect 100569 581710 109191 581712
rect 100569 581707 100635 581710
rect 109125 581707 109191 581710
rect 67633 581362 67699 581365
rect 70166 581362 70226 581468
rect 67633 581360 70226 581362
rect 67633 581304 67638 581360
rect 67694 581304 70226 581360
rect 67633 581302 70226 581304
rect 67633 581299 67699 581302
rect 108941 580818 109007 580821
rect 105892 580816 109007 580818
rect 67817 580682 67883 580685
rect 68553 580682 68619 580685
rect 70166 580682 70226 580788
rect 105892 580760 108946 580816
rect 109002 580760 109007 580816
rect 105892 580758 109007 580760
rect 108941 580755 109007 580758
rect 67817 580680 70226 580682
rect 67817 580624 67822 580680
rect 67878 580624 68558 580680
rect 68614 580624 70226 580680
rect 67817 580622 70226 580624
rect 67817 580619 67883 580622
rect 68553 580619 68619 580622
rect 108849 580138 108915 580141
rect 105892 580136 108915 580138
rect -960 580002 480 580092
rect 105892 580080 108854 580136
rect 108910 580080 108915 580136
rect 105892 580078 108915 580080
rect 108849 580075 108915 580078
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 108389 579458 108455 579461
rect 105892 579456 108455 579458
rect 67357 579186 67423 579189
rect 70166 579186 70226 579428
rect 105892 579400 108394 579456
rect 108450 579400 108455 579456
rect 105892 579398 108455 579400
rect 108389 579395 108455 579398
rect 67357 579184 70226 579186
rect 67357 579128 67362 579184
rect 67418 579128 70226 579184
rect 67357 579126 70226 579128
rect 67357 579123 67423 579126
rect 108941 578778 109007 578781
rect 105892 578776 109007 578778
rect 67633 578506 67699 578509
rect 70166 578506 70226 578748
rect 105892 578720 108946 578776
rect 109002 578720 109007 578776
rect 105892 578718 109007 578720
rect 108941 578715 109007 578718
rect 67633 578504 70226 578506
rect 67633 578448 67638 578504
rect 67694 578448 70226 578504
rect 67633 578446 70226 578448
rect 67633 578443 67699 578446
rect 108941 578098 109007 578101
rect 105892 578096 109007 578098
rect 68185 577826 68251 577829
rect 70166 577826 70226 578068
rect 105892 578040 108946 578096
rect 109002 578040 109007 578096
rect 105892 578038 109007 578040
rect 108941 578035 109007 578038
rect 68185 577824 70226 577826
rect 68185 577768 68190 577824
rect 68246 577768 70226 577824
rect 68185 577766 70226 577768
rect 68185 577763 68251 577766
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 108849 577554 108915 577557
rect 105892 577552 108915 577554
rect 105892 577496 108854 577552
rect 108910 577496 108915 577552
rect 583520 577540 584960 577630
rect 105892 577494 108915 577496
rect 108849 577491 108915 577494
rect 67541 577146 67607 577149
rect 70166 577146 70226 577388
rect 67541 577144 70226 577146
rect 67541 577088 67546 577144
rect 67602 577088 70226 577144
rect 67541 577086 70226 577088
rect 67541 577083 67607 577086
rect 108481 576738 108547 576741
rect 105892 576736 108547 576738
rect 68737 576466 68803 576469
rect 70166 576466 70226 576708
rect 105892 576680 108486 576736
rect 108542 576680 108547 576736
rect 105892 576678 108547 576680
rect 108481 576675 108547 576678
rect 68737 576464 70226 576466
rect 68737 576408 68742 576464
rect 68798 576408 70226 576464
rect 68737 576406 70226 576408
rect 68737 576403 68803 576406
rect 108941 576194 109007 576197
rect 105892 576192 109007 576194
rect 105892 576136 108946 576192
rect 109002 576136 109007 576192
rect 105892 576134 109007 576136
rect 108941 576131 109007 576134
rect 123109 576058 123175 576061
rect 123334 576058 123340 576060
rect 123109 576056 123340 576058
rect 67633 575786 67699 575789
rect 70166 575786 70226 576028
rect 123109 576000 123114 576056
rect 123170 576000 123340 576056
rect 123109 575998 123340 576000
rect 123109 575995 123175 575998
rect 123334 575996 123340 575998
rect 123404 575996 123410 576060
rect 67633 575784 70226 575786
rect 67633 575728 67638 575784
rect 67694 575728 70226 575784
rect 67633 575726 70226 575728
rect 67633 575723 67699 575726
rect 70166 575106 70226 575348
rect 64830 575046 70226 575106
rect 64638 574228 64644 574292
rect 64708 574290 64714 574292
rect 64830 574290 64890 575046
rect 106365 574698 106431 574701
rect 105892 574696 106431 574698
rect 67633 574426 67699 574429
rect 70166 574426 70226 574668
rect 105892 574640 106370 574696
rect 106426 574640 106431 574696
rect 105892 574638 106431 574640
rect 106365 574635 106431 574638
rect 67633 574424 70226 574426
rect 67633 574368 67638 574424
rect 67694 574368 70226 574424
rect 67633 574366 70226 574368
rect 67633 574363 67699 574366
rect 64708 574230 64890 574290
rect 64708 574228 64714 574230
rect 108941 574018 109007 574021
rect 105892 574016 109007 574018
rect 67725 573474 67791 573477
rect 70166 573474 70226 573988
rect 105892 573960 108946 574016
rect 109002 573960 109007 574016
rect 105892 573958 109007 573960
rect 108941 573955 109007 573958
rect 67725 573472 70226 573474
rect 67725 573416 67730 573472
rect 67786 573416 70226 573472
rect 67725 573414 70226 573416
rect 67725 573411 67791 573414
rect 107653 573338 107719 573341
rect 105892 573336 107719 573338
rect 105892 573280 107658 573336
rect 107714 573280 107719 573336
rect 105892 573278 107719 573280
rect 107653 573275 107719 573278
rect 67633 573066 67699 573069
rect 67633 573064 70410 573066
rect 67633 573008 67638 573064
rect 67694 573008 70410 573064
rect 67633 573006 70410 573008
rect 67633 573003 67699 573006
rect 70350 572764 70410 573006
rect 106181 572794 106247 572797
rect 126145 572796 126211 572797
rect 126094 572794 126100 572796
rect 105892 572792 106247 572794
rect 105892 572736 106186 572792
rect 106242 572736 106247 572792
rect 105892 572734 106247 572736
rect 126054 572734 126100 572794
rect 126164 572792 126211 572796
rect 126206 572736 126211 572792
rect 106181 572731 106247 572734
rect 126094 572732 126100 572734
rect 126164 572732 126211 572736
rect 126145 572731 126211 572732
rect 108941 571978 109007 571981
rect 105892 571976 109007 571978
rect 67909 571842 67975 571845
rect 68645 571842 68711 571845
rect 70166 571842 70226 571948
rect 105892 571920 108946 571976
rect 109002 571920 109007 571976
rect 105892 571918 109007 571920
rect 108941 571915 109007 571918
rect 67909 571840 70226 571842
rect 67909 571784 67914 571840
rect 67970 571784 68650 571840
rect 68706 571784 70226 571840
rect 67909 571782 70226 571784
rect 67909 571779 67975 571782
rect 68645 571779 68711 571782
rect 67817 571706 67883 571709
rect 68461 571706 68527 571709
rect 67817 571704 70226 571706
rect 67817 571648 67822 571704
rect 67878 571648 68466 571704
rect 68522 571648 70226 571704
rect 67817 571646 70226 571648
rect 67817 571643 67883 571646
rect 68461 571643 68527 571646
rect 70166 571404 70226 571646
rect 107837 571434 107903 571437
rect 105892 571432 107903 571434
rect 105892 571376 107842 571432
rect 107898 571376 107903 571432
rect 105892 571374 107903 571376
rect 107837 571371 107903 571374
rect 108849 570618 108915 570621
rect 105892 570616 108915 570618
rect 66110 570284 66116 570348
rect 66180 570346 66186 570348
rect 70166 570346 70226 570588
rect 105892 570560 108854 570616
rect 108910 570560 108915 570616
rect 105892 570558 108915 570560
rect 108849 570555 108915 570558
rect 66180 570286 70226 570346
rect 66180 570284 66186 570286
rect 67633 570074 67699 570077
rect 108941 570074 109007 570077
rect 67633 570072 70042 570074
rect 67633 570016 67638 570072
rect 67694 570016 70042 570072
rect 67633 570014 70042 570016
rect 105892 570072 109007 570074
rect 105892 570016 108946 570072
rect 109002 570016 109007 570072
rect 105892 570014 109007 570016
rect 67633 570011 67699 570014
rect 69982 569802 70042 570014
rect 108941 570011 109007 570014
rect 70166 569802 70226 569908
rect 69982 569742 70226 569802
rect 108941 569258 109007 569261
rect 105892 569256 109007 569258
rect 67633 568986 67699 568989
rect 70166 568986 70226 569228
rect 105892 569200 108946 569256
rect 109002 569200 109007 569256
rect 105892 569198 109007 569200
rect 108941 569195 109007 569198
rect 67633 568984 70226 568986
rect 67633 568928 67638 568984
rect 67694 568928 70226 568984
rect 67633 568926 70226 568928
rect 67633 568923 67699 568926
rect 67725 568714 67791 568717
rect 67725 568712 70042 568714
rect 67725 568656 67730 568712
rect 67786 568656 70042 568712
rect 67725 568654 70042 568656
rect 67725 568651 67791 568654
rect 69982 568442 70042 568654
rect 70166 568442 70226 568548
rect 69982 568382 70226 568442
rect 108941 567898 109007 567901
rect 105892 567896 109007 567898
rect 67725 567626 67791 567629
rect 70166 567626 70226 567868
rect 105892 567840 108946 567896
rect 109002 567840 109007 567896
rect 105892 567838 109007 567840
rect 108941 567835 109007 567838
rect 67725 567624 70226 567626
rect 67725 567568 67730 567624
rect 67786 567568 70226 567624
rect 67725 567566 70226 567568
rect 67725 567563 67791 567566
rect 67633 567218 67699 567221
rect 108941 567218 109007 567221
rect 67633 567216 70042 567218
rect 67633 567160 67638 567216
rect 67694 567210 70042 567216
rect 105892 567216 109007 567218
rect 67694 567160 70226 567210
rect 67633 567158 70226 567160
rect 105892 567160 108946 567216
rect 109002 567160 109007 567216
rect 105892 567158 109007 567160
rect 67633 567155 67699 567158
rect 69982 567150 70226 567158
rect 108941 567155 109007 567158
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 108389 566538 108455 566541
rect 105892 566536 108455 566538
rect 105892 566480 108394 566536
rect 108450 566480 108455 566536
rect 105892 566478 108455 566480
rect 108389 566475 108455 566478
rect 70166 565892 70226 565964
rect 67633 565858 67699 565861
rect 69982 565858 70226 565892
rect 108941 565858 109007 565861
rect 67633 565856 70226 565858
rect 67633 565800 67638 565856
rect 67694 565832 70226 565856
rect 105892 565856 109007 565858
rect 67694 565800 70042 565832
rect 67633 565798 70042 565800
rect 105892 565800 108946 565856
rect 109002 565800 109007 565856
rect 105892 565798 109007 565800
rect 67633 565795 67699 565798
rect 108941 565795 109007 565798
rect 108941 565178 109007 565181
rect 105892 565176 109007 565178
rect 67633 564906 67699 564909
rect 70166 564906 70226 565148
rect 105892 565120 108946 565176
rect 109002 565120 109007 565176
rect 105892 565118 109007 565120
rect 108941 565115 109007 565118
rect 67633 564904 70226 564906
rect 67633 564848 67638 564904
rect 67694 564848 70226 564904
rect 67633 564846 70226 564848
rect 67633 564843 67699 564846
rect 67265 564498 67331 564501
rect 106406 564498 106412 564500
rect 67265 564496 70042 564498
rect 67265 564440 67270 564496
rect 67326 564440 70042 564496
rect 67265 564438 70042 564440
rect 67265 564435 67331 564438
rect 69982 564362 70042 564438
rect 70166 564362 70226 564468
rect 105892 564438 106412 564498
rect 106406 564436 106412 564438
rect 106476 564436 106482 564500
rect 69982 564302 70226 564362
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect 108389 563954 108455 563957
rect 105892 563952 108455 563954
rect 105892 563896 108394 563952
rect 108450 563896 108455 563952
rect 105892 563894 108455 563896
rect 108389 563891 108455 563894
rect 67725 563546 67791 563549
rect 70166 563546 70226 563788
rect 67725 563544 70226 563546
rect 67725 563488 67730 563544
rect 67786 563488 70226 563544
rect 67725 563486 70226 563488
rect 67725 563483 67791 563486
rect 67633 563138 67699 563141
rect 107694 563138 107700 563140
rect 67633 563136 70042 563138
rect 67633 563080 67638 563136
rect 67694 563080 70042 563136
rect 67633 563078 70042 563080
rect 67633 563075 67699 563078
rect 69982 563002 70042 563078
rect 70166 563002 70226 563108
rect 105892 563078 107700 563138
rect 107694 563076 107700 563078
rect 107764 563076 107770 563140
rect 69982 562942 70226 563002
rect 108941 562458 109007 562461
rect 105892 562456 109007 562458
rect 67633 562322 67699 562325
rect 70166 562322 70226 562428
rect 105892 562400 108946 562456
rect 109002 562400 109007 562456
rect 105892 562398 109007 562400
rect 108941 562395 109007 562398
rect 67633 562320 70226 562322
rect 67633 562264 67638 562320
rect 67694 562264 70226 562320
rect 67633 562262 70226 562264
rect 67633 562259 67699 562262
rect 67633 562186 67699 562189
rect 67633 562184 70410 562186
rect 67633 562128 67638 562184
rect 67694 562128 70410 562184
rect 67633 562126 70410 562128
rect 67633 562123 67699 562126
rect 70350 561884 70410 562126
rect 108941 561098 109007 561101
rect 105892 561096 109007 561098
rect 67725 560826 67791 560829
rect 70166 560826 70226 561068
rect 105892 561040 108946 561096
rect 109002 561040 109007 561096
rect 105892 561038 109007 561040
rect 108941 561035 109007 561038
rect 67725 560824 70226 560826
rect 67725 560768 67730 560824
rect 67786 560768 70226 560824
rect 67725 560766 70226 560768
rect 67725 560763 67791 560766
rect 67633 560418 67699 560421
rect 106273 560418 106339 560421
rect 108205 560418 108271 560421
rect 67633 560416 70042 560418
rect 67633 560360 67638 560416
rect 67694 560360 70042 560416
rect 105892 560416 108271 560418
rect 67633 560358 70042 560360
rect 67633 560355 67699 560358
rect 69982 560282 70042 560358
rect 70166 560282 70226 560388
rect 105892 560360 106278 560416
rect 106334 560360 108210 560416
rect 108266 560360 108271 560416
rect 105892 560358 108271 560360
rect 106273 560355 106339 560358
rect 108205 560355 108271 560358
rect 69982 560222 70226 560282
rect 108849 559738 108915 559741
rect 105892 559736 108915 559738
rect 105892 559680 108854 559736
rect 108910 559680 108915 559736
rect 105892 559678 108915 559680
rect 108849 559675 108915 559678
rect 67633 559466 67699 559469
rect 67633 559464 70410 559466
rect 67633 559408 67638 559464
rect 67694 559408 70410 559464
rect 67633 559406 70410 559408
rect 67633 559403 67699 559406
rect 70350 559164 70410 559406
rect 108941 559058 109007 559061
rect 105892 559056 109007 559058
rect 105892 559000 108946 559056
rect 109002 559000 109007 559056
rect 105892 558998 109007 559000
rect 108941 558995 109007 558998
rect 68829 558922 68895 558925
rect 68829 558920 70226 558922
rect 68829 558864 68834 558920
rect 68890 558864 70226 558920
rect 68829 558862 70226 558864
rect 68829 558859 68895 558862
rect 70166 558484 70226 558862
rect 108941 558378 109007 558381
rect 105892 558376 109007 558378
rect 105892 558320 108946 558376
rect 109002 558320 109007 558376
rect 105892 558318 109007 558320
rect 108941 558315 109007 558318
rect 107745 557698 107811 557701
rect 105892 557696 107811 557698
rect 62982 557500 62988 557564
rect 63052 557562 63058 557564
rect 70166 557562 70226 557668
rect 105892 557640 107750 557696
rect 107806 557640 107811 557696
rect 105892 557638 107811 557640
rect 107745 557635 107811 557638
rect 63052 557502 70226 557562
rect 63052 557500 63058 557502
rect 68277 557426 68343 557429
rect 69974 557426 69980 557428
rect 68277 557424 69980 557426
rect 68277 557368 68282 557424
rect 68338 557368 69980 557424
rect 68277 557366 69980 557368
rect 68277 557363 68343 557366
rect 69974 557364 69980 557366
rect 70044 557364 70050 557428
rect 108941 557018 109007 557021
rect 105892 557016 109007 557018
rect 67725 556746 67791 556749
rect 70166 556746 70226 556988
rect 105892 556960 108946 557016
rect 109002 556960 109007 557016
rect 105892 556958 109007 556960
rect 108941 556955 109007 556958
rect 67725 556744 70226 556746
rect 67725 556688 67730 556744
rect 67786 556688 70226 556744
rect 67725 556686 70226 556688
rect 67725 556683 67791 556686
rect 107653 556338 107719 556341
rect 105892 556336 107719 556338
rect 67633 556202 67699 556205
rect 70166 556202 70226 556308
rect 105892 556280 107658 556336
rect 107714 556280 107719 556336
rect 105892 556278 107719 556280
rect 107653 556275 107719 556278
rect 67633 556200 70226 556202
rect 67633 556144 67638 556200
rect 67694 556144 70226 556200
rect 67633 556142 70226 556144
rect 67633 556139 67699 556142
rect 108849 555794 108915 555797
rect 105892 555792 108915 555794
rect 105892 555736 108854 555792
rect 108910 555736 108915 555792
rect 105892 555734 108915 555736
rect 108849 555731 108915 555734
rect 67725 555386 67791 555389
rect 70166 555386 70226 555628
rect 67725 555384 70226 555386
rect 67725 555328 67730 555384
rect 67786 555328 70226 555384
rect 67725 555326 70226 555328
rect 67725 555323 67791 555326
rect 67633 554842 67699 554845
rect 70166 554842 70226 554948
rect 67633 554840 70226 554842
rect 67633 554784 67638 554840
rect 67694 554784 70226 554840
rect 67633 554782 70226 554784
rect 67633 554779 67699 554782
rect 108941 554298 109007 554301
rect 105892 554296 109007 554298
rect -960 553890 480 553980
rect 68870 553964 68876 554028
rect 68940 554026 68946 554028
rect 70166 554026 70226 554268
rect 105892 554240 108946 554296
rect 109002 554240 109007 554296
rect 105892 554238 109007 554240
rect 108941 554235 109007 554238
rect 111558 554026 111564 554028
rect 68940 553966 70226 554026
rect 105862 553966 111564 554026
rect 68940 553964 68946 553966
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 105862 553724 105922 553966
rect 111558 553964 111564 553966
rect 111628 554026 111634 554028
rect 129917 554026 129983 554029
rect 111628 554024 129983 554026
rect 111628 553968 129922 554024
rect 129978 553968 129983 554024
rect 111628 553966 129983 553968
rect 111628 553964 111634 553966
rect 129917 553963 129983 553966
rect 67633 553482 67699 553485
rect 70166 553482 70226 553588
rect 67633 553480 70226 553482
rect 67633 553424 67638 553480
rect 67694 553424 70226 553480
rect 67633 553422 70226 553424
rect 67633 553419 67699 553422
rect 108113 552938 108179 552941
rect 105892 552936 108179 552938
rect 105892 552880 108118 552936
rect 108174 552880 108179 552936
rect 105892 552878 108179 552880
rect 108113 552875 108179 552878
rect 106038 552604 106044 552668
rect 106108 552666 106114 552668
rect 107837 552666 107903 552669
rect 106108 552664 107903 552666
rect 106108 552608 107842 552664
rect 107898 552608 107903 552664
rect 106108 552606 107903 552608
rect 106108 552604 106114 552606
rect 107837 552603 107903 552606
rect 106774 552258 106780 552260
rect 67633 552122 67699 552125
rect 70166 552122 70226 552228
rect 105892 552198 106780 552258
rect 106774 552196 106780 552198
rect 106844 552196 106850 552260
rect 67633 552120 70226 552122
rect 67633 552064 67638 552120
rect 67694 552064 70226 552120
rect 67633 552062 70226 552064
rect 67633 552059 67699 552062
rect 107009 551578 107075 551581
rect 105892 551576 107075 551578
rect 67633 551306 67699 551309
rect 70166 551306 70226 551548
rect 105892 551520 107014 551576
rect 107070 551520 107075 551576
rect 105892 551518 107075 551520
rect 107009 551515 107075 551518
rect 67633 551304 70226 551306
rect 67633 551248 67638 551304
rect 67694 551248 70226 551304
rect 67633 551246 70226 551248
rect 67633 551243 67699 551246
rect 583520 551020 584960 551260
rect 108941 550898 109007 550901
rect 105892 550896 109007 550898
rect 68921 550762 68987 550765
rect 70166 550762 70226 550868
rect 105892 550840 108946 550896
rect 109002 550840 109007 550896
rect 105892 550838 109007 550840
rect 108941 550835 109007 550838
rect 68921 550760 70226 550762
rect 68921 550704 68926 550760
rect 68982 550704 70226 550760
rect 68921 550702 70226 550704
rect 68921 550699 68987 550702
rect 108849 550218 108915 550221
rect 105892 550216 108915 550218
rect 67725 549946 67791 549949
rect 70166 549946 70226 550188
rect 105892 550160 108854 550216
rect 108910 550160 108915 550216
rect 105892 550158 108915 550160
rect 108849 550155 108915 550158
rect 67725 549944 70226 549946
rect 67725 549888 67730 549944
rect 67786 549888 70226 549944
rect 67725 549886 70226 549888
rect 67725 549883 67791 549886
rect 108941 549538 109007 549541
rect 105892 549536 109007 549538
rect 67633 549402 67699 549405
rect 70166 549402 70226 549508
rect 105892 549480 108946 549536
rect 109002 549480 109007 549536
rect 105892 549478 109007 549480
rect 108941 549475 109007 549478
rect 67633 549400 70226 549402
rect 67633 549344 67638 549400
rect 67694 549344 70226 549400
rect 67633 549342 70226 549344
rect 67633 549339 67699 549342
rect 108941 548858 109007 548861
rect 105892 548856 109007 548858
rect 68134 548524 68140 548588
rect 68204 548586 68210 548588
rect 70166 548586 70226 548828
rect 105892 548800 108946 548856
rect 109002 548800 109007 548856
rect 105892 548798 109007 548800
rect 108941 548795 109007 548798
rect 68204 548526 70226 548586
rect 68204 548524 68210 548526
rect 67633 548042 67699 548045
rect 70166 548042 70226 548148
rect 67633 548040 70226 548042
rect 67633 547984 67638 548040
rect 67694 547984 70226 548040
rect 67633 547982 70226 547984
rect 67633 547979 67699 547982
rect 108941 547498 109007 547501
rect 105892 547496 109007 547498
rect 70166 547226 70226 547468
rect 105892 547440 108946 547496
rect 109002 547440 109007 547496
rect 105892 547438 109007 547440
rect 108941 547435 109007 547438
rect 64830 547166 70226 547226
rect 61878 546620 61884 546684
rect 61948 546682 61954 546684
rect 64830 546682 64890 547166
rect 107929 546818 107995 546821
rect 105892 546816 107995 546818
rect 61948 546622 64890 546682
rect 61948 546620 61954 546622
rect 67633 546546 67699 546549
rect 70166 546546 70226 546788
rect 105892 546760 107934 546816
rect 107990 546760 107995 546816
rect 105892 546758 107995 546760
rect 107929 546755 107995 546758
rect 67633 546544 70226 546546
rect 67633 546488 67638 546544
rect 67694 546488 70226 546544
rect 67633 546486 70226 546488
rect 67633 546483 67699 546486
rect 108941 546138 109007 546141
rect 105892 546136 109007 546138
rect 105892 546080 108946 546136
rect 109002 546080 109007 546136
rect 105892 546078 109007 546080
rect 108941 546075 109007 546078
rect 108941 545458 109007 545461
rect 105892 545456 109007 545458
rect 66662 545124 66668 545188
rect 66732 545186 66738 545188
rect 69197 545186 69263 545189
rect 70166 545186 70226 545428
rect 105892 545400 108946 545456
rect 109002 545400 109007 545456
rect 105892 545398 109007 545400
rect 108941 545395 109007 545398
rect 66732 545184 70226 545186
rect 66732 545128 69202 545184
rect 69258 545128 70226 545184
rect 66732 545126 70226 545128
rect 66732 545124 66738 545126
rect 69197 545123 69263 545126
rect 68829 544506 68895 544509
rect 70166 544506 70226 544748
rect 68829 544504 70226 544506
rect 68829 544448 68834 544504
rect 68890 544448 70226 544504
rect 68829 544446 70226 544448
rect 105862 544506 105922 544748
rect 111701 544506 111767 544509
rect 105862 544504 113190 544506
rect 105862 544448 111706 544504
rect 111762 544448 113190 544504
rect 105862 544446 113190 544448
rect 68829 544443 68895 544446
rect 111701 544443 111767 544446
rect 113130 544370 113190 544446
rect 115974 544370 115980 544372
rect 113130 544310 115980 544370
rect 115974 544308 115980 544310
rect 116044 544308 116050 544372
rect 67725 543962 67791 543965
rect 68277 543962 68343 543965
rect 70166 543962 70226 544068
rect 67725 543960 70226 543962
rect 67725 543904 67730 543960
rect 67786 543904 68282 543960
rect 68338 543904 70226 543960
rect 67725 543902 70226 543904
rect 67725 543899 67791 543902
rect 68277 543899 68343 543902
rect 105678 543829 105738 544068
rect 105678 543824 105787 543829
rect 105678 543768 105726 543824
rect 105782 543768 105787 543824
rect 105678 543766 105787 543768
rect 105721 543763 105787 543766
rect 108941 543418 109007 543421
rect 105892 543416 109007 543418
rect 68001 543282 68067 543285
rect 69013 543282 69079 543285
rect 70166 543282 70226 543388
rect 105892 543360 108946 543416
rect 109002 543360 109007 543416
rect 105892 543358 109007 543360
rect 108941 543355 109007 543358
rect 68001 543280 70226 543282
rect 68001 543224 68006 543280
rect 68062 543224 69018 543280
rect 69074 543224 70226 543280
rect 68001 543222 70226 543224
rect 68001 543219 68067 543222
rect 69013 543219 69079 543222
rect 108246 542738 108252 542740
rect 67633 542602 67699 542605
rect 70166 542602 70226 542708
rect 105892 542678 108252 542738
rect 108246 542676 108252 542678
rect 108316 542676 108322 542740
rect 67633 542600 70226 542602
rect 67633 542544 67638 542600
rect 67694 542544 70226 542600
rect 67633 542542 70226 542544
rect 67633 542539 67699 542542
rect 106917 542058 106983 542061
rect 105892 542056 106983 542058
rect 67725 541786 67791 541789
rect 70166 541786 70226 542028
rect 105892 542000 106922 542056
rect 106978 542000 106983 542056
rect 105892 541998 106983 542000
rect 106917 541995 106983 541998
rect 67725 541784 70226 541786
rect 67725 541728 67730 541784
rect 67786 541728 70226 541784
rect 67725 541726 70226 541728
rect 67725 541723 67791 541726
rect 67633 541242 67699 541245
rect 70166 541242 70226 541348
rect 67633 541240 70226 541242
rect 67633 541184 67638 541240
rect 67694 541184 70226 541240
rect 67633 541182 70226 541184
rect 67633 541179 67699 541182
rect -960 540684 480 540924
rect 107837 540698 107903 540701
rect 105892 540696 107903 540698
rect 105892 540668 107842 540696
rect 67633 540154 67699 540157
rect 70166 540154 70226 540668
rect 105862 540640 107842 540668
rect 107898 540640 107903 540696
rect 105862 540638 107903 540640
rect 105862 540429 105922 540638
rect 107837 540635 107903 540638
rect 105813 540424 105922 540429
rect 105813 540368 105818 540424
rect 105874 540368 105922 540424
rect 105813 540366 105922 540368
rect 105813 540363 105879 540366
rect 67633 540152 70226 540154
rect 67633 540096 67638 540152
rect 67694 540096 70226 540152
rect 67633 540094 70226 540096
rect 67633 540091 67699 540094
rect 108941 540018 109007 540021
rect 105892 540016 109007 540018
rect 105892 539960 108946 540016
rect 109002 539960 109007 540016
rect 105892 539958 109007 539960
rect 108941 539955 109007 539958
rect 80329 538114 80395 538117
rect 115054 538114 115060 538116
rect 80329 538112 115060 538114
rect 80329 538056 80334 538112
rect 80390 538056 115060 538112
rect 80329 538054 115060 538056
rect 80329 538051 80395 538054
rect 115054 538052 115060 538054
rect 115124 538052 115130 538116
rect 100937 537978 101003 537981
rect 101990 537978 101996 537980
rect 100937 537976 101996 537978
rect 100937 537920 100942 537976
rect 100998 537920 101996 537976
rect 100937 537918 101996 537920
rect 100937 537915 101003 537918
rect 101990 537916 101996 537918
rect 102060 537978 102066 537980
rect 130377 537978 130443 537981
rect 102060 537976 130443 537978
rect 102060 537920 130382 537976
rect 130438 537920 130443 537976
rect 102060 537918 130443 537920
rect 102060 537916 102066 537918
rect 130377 537915 130443 537918
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 46749 537434 46815 537437
rect 80329 537434 80395 537437
rect 46749 537432 80395 537434
rect 46749 537376 46754 537432
rect 46810 537376 80334 537432
rect 80390 537376 80395 537432
rect 46749 537374 80395 537376
rect 46749 537371 46815 537374
rect 80329 537371 80395 537374
rect 97073 536890 97139 536893
rect 98494 536890 98500 536892
rect 97073 536888 98500 536890
rect 97073 536832 97078 536888
rect 97134 536832 98500 536888
rect 97073 536830 98500 536832
rect 97073 536827 97139 536830
rect 98494 536828 98500 536830
rect 98564 536828 98570 536892
rect 92565 531994 92631 531997
rect 110638 531994 110644 531996
rect 92565 531992 110644 531994
rect 92565 531936 92570 531992
rect 92626 531936 110644 531992
rect 92565 531934 110644 531936
rect 92565 531931 92631 531934
rect 110638 531932 110644 531934
rect 110708 531932 110714 531996
rect -960 527914 480 528004
rect 3141 527914 3207 527917
rect -960 527912 3207 527914
rect -960 527856 3146 527912
rect 3202 527856 3207 527912
rect -960 527854 3207 527856
rect -960 527764 480 527854
rect 3141 527851 3207 527854
rect 579797 524514 579863 524517
rect 583520 524514 584960 524604
rect 579797 524512 584960 524514
rect 579797 524456 579802 524512
rect 579858 524456 584960 524512
rect 579797 524454 584960 524456
rect 579797 524451 579863 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 57830 498748 57836 498812
rect 57900 498810 57906 498812
rect 86125 498810 86191 498813
rect 57900 498808 86191 498810
rect 57900 498752 86130 498808
rect 86186 498752 86191 498808
rect 57900 498750 86191 498752
rect 57900 498748 57906 498750
rect 86125 498747 86191 498750
rect 583520 497844 584960 498084
rect 90357 497450 90423 497453
rect 111742 497450 111748 497452
rect 90357 497448 111748 497450
rect 90357 497392 90362 497448
rect 90418 497392 111748 497448
rect 90357 497390 111748 497392
rect 90357 497387 90423 497390
rect 111742 497388 111748 497390
rect 111812 497388 111818 497452
rect 86769 496226 86835 496229
rect 111926 496226 111932 496228
rect 86769 496224 111932 496226
rect 86769 496168 86774 496224
rect 86830 496168 111932 496224
rect 86769 496166 111932 496168
rect 86769 496163 86835 496166
rect 111926 496164 111932 496166
rect 111996 496164 112002 496228
rect 89621 496090 89687 496093
rect 124254 496090 124260 496092
rect 89621 496088 124260 496090
rect 89621 496032 89626 496088
rect 89682 496032 124260 496088
rect 89621 496030 124260 496032
rect 89621 496027 89687 496030
rect 124254 496028 124260 496030
rect 124324 496090 124330 496092
rect 127341 496090 127407 496093
rect 124324 496088 127407 496090
rect 124324 496032 127346 496088
rect 127402 496032 127407 496088
rect 124324 496030 127407 496032
rect 124324 496028 124330 496030
rect 127341 496027 127407 496030
rect 111793 494730 111859 494733
rect 118918 494730 118924 494732
rect 111793 494728 118924 494730
rect 111793 494672 111798 494728
rect 111854 494672 118924 494728
rect 111793 494670 118924 494672
rect 111793 494667 111859 494670
rect 118918 494668 118924 494670
rect 118988 494668 118994 494732
rect 54886 493308 54892 493372
rect 54956 493370 54962 493372
rect 57697 493370 57763 493373
rect 54956 493368 57763 493370
rect 54956 493312 57702 493368
rect 57758 493312 57763 493368
rect 54956 493310 57763 493312
rect 54956 493308 54962 493310
rect 57697 493307 57763 493310
rect 95785 493370 95851 493373
rect 118734 493370 118740 493372
rect 95785 493368 118740 493370
rect 95785 493312 95790 493368
rect 95846 493312 118740 493368
rect 95785 493310 118740 493312
rect 95785 493307 95851 493310
rect 118734 493308 118740 493310
rect 118804 493370 118810 493372
rect 129733 493370 129799 493373
rect 118804 493368 129799 493370
rect 118804 493312 129738 493368
rect 129794 493312 129799 493368
rect 118804 493310 129799 493312
rect 118804 493308 118810 493310
rect 129733 493307 129799 493310
rect 57646 492628 57652 492692
rect 57716 492690 57722 492692
rect 58617 492690 58683 492693
rect 57716 492688 58683 492690
rect 57716 492632 58622 492688
rect 58678 492632 58683 492688
rect 57716 492630 58683 492632
rect 57716 492628 57722 492630
rect 58617 492627 58683 492630
rect 63493 491330 63559 491333
rect 580901 491330 580967 491333
rect 63493 491328 580967 491330
rect 63493 491272 63498 491328
rect 63554 491272 580906 491328
rect 580962 491272 580967 491328
rect 63493 491270 580967 491272
rect 63493 491267 63559 491270
rect 580901 491267 580967 491270
rect 87689 490650 87755 490653
rect 95049 490650 95115 490653
rect 100702 490650 100708 490652
rect 87689 490648 100708 490650
rect 87689 490592 87694 490648
rect 87750 490592 95054 490648
rect 95110 490592 100708 490648
rect 87689 490590 100708 490592
rect 87689 490587 87755 490590
rect 95049 490587 95115 490590
rect 100702 490588 100708 490590
rect 100772 490588 100778 490652
rect 97073 490514 97139 490517
rect 122833 490514 122899 490517
rect 141141 490514 141207 490517
rect 97073 490512 141207 490514
rect 97073 490456 97078 490512
rect 97134 490456 122838 490512
rect 122894 490456 141146 490512
rect 141202 490456 141207 490512
rect 97073 490454 141207 490456
rect 97073 490451 97139 490454
rect 122833 490451 122899 490454
rect 141141 490451 141207 490454
rect 69749 489970 69815 489973
rect 69749 489968 70226 489970
rect 69749 489912 69754 489968
rect 69810 489912 70226 489968
rect 69749 489910 70226 489912
rect 69749 489907 69815 489910
rect 70166 489804 70226 489910
rect 48078 489092 48084 489156
rect 48148 489154 48154 489156
rect 69841 489154 69907 489157
rect 48148 489152 69907 489154
rect 48148 489096 69846 489152
rect 69902 489096 69907 489152
rect 48148 489094 69907 489096
rect 48148 489092 48154 489094
rect 69841 489091 69907 489094
rect -960 488596 480 488836
rect 99790 488746 99850 488988
rect 103421 488746 103487 488749
rect 99790 488744 103487 488746
rect 99790 488688 103426 488744
rect 103482 488688 103487 488744
rect 99790 488686 103487 488688
rect 103421 488683 103487 488686
rect 102869 488610 102935 488613
rect 99790 488608 102935 488610
rect 99790 488552 102874 488608
rect 102930 488552 102935 488608
rect 99790 488550 102935 488552
rect 99790 488444 99850 488550
rect 102869 488547 102935 488550
rect 67633 487930 67699 487933
rect 70166 487930 70226 488308
rect 103329 488066 103395 488069
rect 67633 487928 70226 487930
rect 67633 487872 67638 487928
rect 67694 487872 70226 487928
rect 67633 487870 70226 487872
rect 99790 488064 103395 488066
rect 99790 488008 103334 488064
rect 103390 488008 103395 488064
rect 99790 488006 103395 488008
rect 67633 487867 67699 487870
rect 99790 487764 99850 488006
rect 103329 488003 103395 488006
rect 67633 487250 67699 487253
rect 70166 487250 70226 487628
rect 67633 487248 70226 487250
rect 67633 487192 67638 487248
rect 67694 487192 70226 487248
rect 67633 487190 70226 487192
rect 67633 487187 67699 487190
rect 99322 487188 99328 487252
rect 99392 487250 99398 487252
rect 103605 487250 103671 487253
rect 114369 487252 114435 487253
rect 114318 487250 114324 487252
rect 99392 487248 103671 487250
rect 99392 487192 103610 487248
rect 103666 487192 103671 487248
rect 99392 487190 103671 487192
rect 114278 487190 114324 487250
rect 114388 487248 114435 487252
rect 114430 487192 114435 487248
rect 99392 487188 99398 487190
rect 103605 487187 103671 487190
rect 114318 487188 114324 487190
rect 114388 487188 114435 487192
rect 114369 487187 114435 487188
rect 67633 486570 67699 486573
rect 70166 486570 70226 486948
rect 67633 486568 70226 486570
rect 67633 486512 67638 486568
rect 67694 486512 70226 486568
rect 67633 486510 70226 486512
rect 99606 486570 99666 486948
rect 103329 486570 103395 486573
rect 99606 486568 103395 486570
rect 99606 486512 103334 486568
rect 103390 486512 103395 486568
rect 99606 486510 103395 486512
rect 67633 486507 67699 486510
rect 103329 486507 103395 486510
rect 68093 486026 68159 486029
rect 69197 486026 69263 486029
rect 70350 486026 70410 486268
rect 68093 486024 70410 486026
rect 68093 485968 68098 486024
rect 68154 485968 69202 486024
rect 69258 485968 70410 486024
rect 68093 485966 70410 485968
rect 99606 486026 99666 486268
rect 103421 486026 103487 486029
rect 99606 486024 103487 486026
rect 99606 485968 103426 486024
rect 103482 485968 103487 486024
rect 99606 485966 103487 485968
rect 68093 485963 68159 485966
rect 69197 485963 69263 485966
rect 103421 485963 103487 485966
rect 117221 485754 117287 485757
rect 124438 485754 124444 485756
rect 117221 485752 124444 485754
rect 117221 485696 117226 485752
rect 117282 485696 124444 485752
rect 117221 485694 124444 485696
rect 117221 485691 117287 485694
rect 124438 485692 124444 485694
rect 124508 485692 124514 485756
rect 67633 485210 67699 485213
rect 70166 485210 70226 485588
rect 99606 485346 99666 485588
rect 102225 485346 102291 485349
rect 99606 485344 102291 485346
rect 99606 485288 102230 485344
rect 102286 485288 102291 485344
rect 99606 485286 102291 485288
rect 102225 485283 102291 485286
rect 67633 485208 70226 485210
rect 67633 485152 67638 485208
rect 67694 485152 70226 485208
rect 67633 485150 70226 485152
rect 67633 485147 67699 485150
rect 68369 484666 68435 484669
rect 70166 484666 70226 484908
rect 70526 484666 70532 484668
rect 68369 484664 70532 484666
rect 68369 484608 68374 484664
rect 68430 484608 70532 484664
rect 68369 484606 70532 484608
rect 68369 484603 68435 484606
rect 70526 484604 70532 484606
rect 70596 484604 70602 484668
rect 99790 484666 99850 484908
rect 102225 484666 102291 484669
rect 99790 484664 102291 484666
rect 99790 484608 102230 484664
rect 102286 484608 102291 484664
rect 99790 484606 102291 484608
rect 102225 484603 102291 484606
rect 580901 484666 580967 484669
rect 583520 484666 584960 484756
rect 580901 484664 584960 484666
rect 580901 484608 580906 484664
rect 580962 484608 584960 484664
rect 580901 484606 584960 484608
rect 580901 484603 580967 484606
rect 583520 484516 584960 484606
rect 125685 484394 125751 484397
rect 126094 484394 126100 484396
rect 125685 484392 126100 484394
rect 125685 484336 125690 484392
rect 125746 484336 126100 484392
rect 125685 484334 126100 484336
rect 125685 484331 125751 484334
rect 126094 484332 126100 484334
rect 126164 484332 126170 484396
rect 70166 483578 70226 484228
rect 102225 483850 102291 483853
rect 99790 483848 102291 483850
rect 99790 483792 102230 483848
rect 102286 483792 102291 483848
rect 99790 483790 102291 483792
rect 99790 483684 99850 483790
rect 102225 483787 102291 483790
rect 123201 483714 123267 483717
rect 123334 483714 123340 483716
rect 123201 483712 123340 483714
rect 123201 483656 123206 483712
rect 123262 483656 123340 483712
rect 123201 483654 123340 483656
rect 123201 483651 123267 483654
rect 123334 483652 123340 483654
rect 123404 483652 123410 483716
rect 60690 483518 70226 483578
rect 58566 482972 58572 483036
rect 58636 483034 58642 483036
rect 60690 483034 60750 483518
rect 58636 482974 60750 483034
rect 69982 483110 70226 483170
rect 58636 482972 58642 482974
rect 53741 482898 53807 482901
rect 58574 482898 58634 482972
rect 53741 482896 58634 482898
rect 53741 482840 53746 482896
rect 53802 482840 58634 482896
rect 53741 482838 58634 482840
rect 69105 482898 69171 482901
rect 69982 482898 70042 483110
rect 70166 483004 70226 483110
rect 69105 482896 70042 482898
rect 69105 482840 69110 482896
rect 69166 482840 70042 482896
rect 69105 482838 70042 482840
rect 53741 482835 53807 482838
rect 69105 482835 69171 482838
rect 67633 482626 67699 482629
rect 99606 482626 99666 482868
rect 102317 482626 102383 482629
rect 67633 482624 70226 482626
rect 67633 482568 67638 482624
rect 67694 482568 70226 482624
rect 67633 482566 70226 482568
rect 99606 482624 102383 482626
rect 99606 482568 102322 482624
rect 102378 482568 102383 482624
rect 99606 482566 102383 482568
rect 67633 482563 67699 482566
rect 70166 482324 70226 482566
rect 102317 482563 102383 482566
rect 102225 482490 102291 482493
rect 99790 482488 102291 482490
rect 99790 482432 102230 482488
rect 102286 482432 102291 482488
rect 99790 482430 102291 482432
rect 99790 482324 99850 482430
rect 102225 482427 102291 482430
rect 99790 481750 100034 481810
rect 99790 481644 99850 481750
rect 99974 481538 100034 481750
rect 102225 481538 102291 481541
rect 99974 481536 102291 481538
rect 67633 481130 67699 481133
rect 70166 481130 70226 481508
rect 99974 481480 102230 481536
rect 102286 481480 102291 481536
rect 99974 481478 102291 481480
rect 102225 481475 102291 481478
rect 104893 481538 104959 481541
rect 106038 481538 106044 481540
rect 104893 481536 106044 481538
rect 104893 481480 104898 481536
rect 104954 481480 106044 481536
rect 104893 481478 106044 481480
rect 104893 481475 104959 481478
rect 106038 481476 106044 481478
rect 106108 481476 106114 481540
rect 102317 481266 102383 481269
rect 67633 481128 70226 481130
rect 67633 481072 67638 481128
rect 67694 481072 70226 481128
rect 67633 481070 70226 481072
rect 99790 481264 102383 481266
rect 99790 481208 102322 481264
rect 102378 481208 102383 481264
rect 99790 481206 102383 481208
rect 67633 481067 67699 481070
rect 99790 480964 99850 481206
rect 102317 481203 102383 481206
rect 53598 480796 53604 480860
rect 53668 480858 53674 480860
rect 59261 480858 59327 480861
rect 53668 480856 59327 480858
rect 53668 480800 59266 480856
rect 59322 480800 59327 480856
rect 53668 480798 59327 480800
rect 53668 480796 53674 480798
rect 59261 480795 59327 480798
rect 65926 480524 65932 480588
rect 65996 480586 66002 480588
rect 67357 480586 67423 480589
rect 70350 480586 70410 480828
rect 65996 480584 70410 480586
rect 65996 480528 67362 480584
rect 67418 480528 70410 480584
rect 65996 480526 70410 480528
rect 65996 480524 66002 480526
rect 67357 480523 67423 480526
rect 104893 480314 104959 480317
rect 151813 480314 151879 480317
rect 104893 480312 151879 480314
rect 99790 480210 100034 480270
rect 104893 480256 104898 480312
rect 104954 480256 151818 480312
rect 151874 480256 151879 480312
rect 104893 480254 151879 480256
rect 104893 480251 104959 480254
rect 151813 480251 151879 480254
rect 99790 480148 99850 480210
rect 99974 480178 100034 480210
rect 101949 480178 102015 480181
rect 99974 480176 102015 480178
rect 67541 479906 67607 479909
rect 70350 479906 70410 480148
rect 99974 480120 101954 480176
rect 102010 480120 102015 480176
rect 99974 480118 102015 480120
rect 101949 480115 102015 480118
rect 102225 479906 102291 479909
rect 67541 479904 70410 479906
rect 67541 479848 67546 479904
rect 67602 479848 70410 479904
rect 67541 479846 70410 479848
rect 99790 479904 102291 479906
rect 99790 479848 102230 479904
rect 102286 479848 102291 479904
rect 99790 479846 102291 479848
rect 67541 479843 67607 479846
rect 68369 479770 68435 479773
rect 68369 479768 70226 479770
rect 68369 479712 68374 479768
rect 68430 479712 70226 479768
rect 68369 479710 70226 479712
rect 68369 479707 68435 479710
rect 70166 479604 70226 479710
rect 99790 479604 99850 479846
rect 102225 479843 102291 479846
rect 113081 479498 113147 479501
rect 117998 479498 118004 479500
rect 113081 479496 118004 479498
rect 113081 479440 113086 479496
rect 113142 479440 118004 479496
rect 113081 479438 118004 479440
rect 113081 479435 113147 479438
rect 117998 479436 118004 479438
rect 118068 479436 118074 479500
rect 61510 478484 61516 478548
rect 61580 478546 61586 478548
rect 67449 478546 67515 478549
rect 70350 478546 70410 478788
rect 61580 478544 70410 478546
rect 61580 478488 67454 478544
rect 67510 478488 70410 478544
rect 61580 478486 70410 478488
rect 61580 478484 61586 478486
rect 67449 478483 67515 478486
rect 99790 477730 99850 478108
rect 102869 477730 102935 477733
rect 99790 477728 102935 477730
rect 99790 477672 102874 477728
rect 102930 477672 102935 477728
rect 99790 477670 102935 477672
rect 102869 477667 102935 477670
rect 64638 477396 64644 477460
rect 64708 477458 64714 477460
rect 66897 477458 66963 477461
rect 64708 477456 66963 477458
rect 64708 477400 66902 477456
rect 66958 477400 66963 477456
rect 64708 477398 66963 477400
rect 64708 477396 64714 477398
rect 66897 477395 66963 477398
rect 68645 477186 68711 477189
rect 70350 477186 70410 477428
rect 68645 477184 70410 477186
rect 68645 477128 68650 477184
rect 68706 477128 70410 477184
rect 68645 477126 70410 477128
rect 99790 477186 99850 477428
rect 102409 477186 102475 477189
rect 99790 477184 102475 477186
rect 99790 477128 102414 477184
rect 102470 477128 102475 477184
rect 99790 477126 102475 477128
rect 68645 477123 68711 477126
rect 102409 477123 102475 477126
rect 67633 477050 67699 477053
rect 102225 477050 102291 477053
rect 67633 477048 70226 477050
rect 67633 476992 67638 477048
rect 67694 476992 70226 477048
rect 67633 476990 70226 476992
rect 67633 476987 67699 476990
rect 70166 476884 70226 476990
rect 99790 477048 102291 477050
rect 99790 476992 102230 477048
rect 102286 476992 102291 477048
rect 99790 476990 102291 476992
rect 99790 476884 99850 476990
rect 102225 476987 102291 476990
rect 66897 476506 66963 476509
rect 102317 476506 102383 476509
rect 66897 476504 70410 476506
rect 66897 476448 66902 476504
rect 66958 476448 70410 476504
rect 66897 476446 70410 476448
rect 66897 476443 66963 476446
rect 70350 476204 70410 476446
rect 99790 476504 102383 476506
rect 99790 476448 102322 476504
rect 102378 476448 102383 476504
rect 99790 476446 102383 476448
rect 99790 476204 99850 476446
rect 102317 476443 102383 476446
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 67633 475690 67699 475693
rect 102225 475690 102291 475693
rect 67633 475688 70226 475690
rect 67633 475632 67638 475688
rect 67694 475632 70226 475688
rect 67633 475630 70226 475632
rect 67633 475627 67699 475630
rect 70166 475524 70226 475630
rect 99790 475688 102291 475690
rect 99790 475632 102230 475688
rect 102286 475632 102291 475688
rect 99790 475630 102291 475632
rect 99790 475524 99850 475630
rect 102225 475627 102291 475630
rect 67725 475146 67791 475149
rect 102317 475146 102383 475149
rect 67725 475144 70226 475146
rect 67725 475088 67730 475144
rect 67786 475088 70226 475144
rect 67725 475086 70226 475088
rect 67725 475083 67791 475086
rect 70166 474844 70226 475086
rect 99790 475144 102383 475146
rect 99790 475088 102322 475144
rect 102378 475088 102383 475144
rect 99790 475086 102383 475088
rect 99790 474844 99850 475086
rect 102317 475083 102383 475086
rect 67633 474330 67699 474333
rect 102225 474330 102291 474333
rect 67633 474328 70226 474330
rect 67633 474272 67638 474328
rect 67694 474272 70226 474328
rect 67633 474270 70226 474272
rect 67633 474267 67699 474270
rect 70166 474164 70226 474270
rect 99790 474328 102291 474330
rect 99790 474272 102230 474328
rect 102286 474272 102291 474328
rect 99790 474270 102291 474272
rect 99790 474164 99850 474270
rect 102225 474267 102291 474270
rect 103421 474058 103487 474061
rect 106406 474058 106412 474060
rect 103421 474056 106412 474058
rect 103421 474000 103426 474056
rect 103482 474000 106412 474056
rect 103421 473998 106412 474000
rect 103421 473995 103487 473998
rect 106406 473996 106412 473998
rect 106476 473996 106482 474060
rect 67633 473650 67699 473653
rect 67633 473648 70226 473650
rect 67633 473592 67638 473648
rect 67694 473592 70226 473648
rect 67633 473590 70226 473592
rect 67633 473587 67699 473590
rect 70166 473484 70226 473590
rect 102225 472970 102291 472973
rect 99790 472968 102291 472970
rect 99790 472912 102230 472968
rect 102286 472912 102291 472968
rect 99790 472910 102291 472912
rect 99790 472804 99850 472910
rect 102225 472907 102291 472910
rect 67633 472562 67699 472565
rect 67633 472560 70226 472562
rect 67633 472504 67638 472560
rect 67694 472504 70226 472560
rect 67633 472502 70226 472504
rect 67633 472499 67699 472502
rect 70166 472124 70226 472502
rect 102317 472426 102383 472429
rect 99790 472424 102383 472426
rect 99790 472368 102322 472424
rect 102378 472368 102383 472424
rect 99790 472366 102383 472368
rect 99790 472124 99850 472366
rect 102317 472363 102383 472366
rect 107694 471820 107700 471884
rect 107764 471882 107770 471884
rect 108297 471882 108363 471885
rect 107764 471880 108363 471882
rect 107764 471824 108302 471880
rect 108358 471824 108363 471880
rect 107764 471822 108363 471824
rect 107764 471820 107770 471822
rect 108297 471819 108363 471822
rect 66110 471548 66116 471612
rect 66180 471610 66186 471612
rect 102225 471610 102291 471613
rect 66180 471550 70226 471610
rect 66180 471548 66186 471550
rect 70166 471444 70226 471550
rect 99790 471608 102291 471610
rect 99790 471552 102230 471608
rect 102286 471552 102291 471608
rect 99790 471550 102291 471552
rect 99790 471444 99850 471550
rect 102225 471547 102291 471550
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 67633 471066 67699 471069
rect 108297 471066 108363 471069
rect 67633 471064 70226 471066
rect 67633 471008 67638 471064
rect 67694 471008 70226 471064
rect 67633 471006 70226 471008
rect 67633 471003 67699 471006
rect 60590 470732 60596 470796
rect 60660 470794 60666 470796
rect 66110 470794 66116 470796
rect 60660 470734 66116 470794
rect 60660 470732 60666 470734
rect 66110 470732 66116 470734
rect 66180 470732 66186 470796
rect 70166 470764 70226 471006
rect 99790 471064 108363 471066
rect 99790 471008 108302 471064
rect 108358 471008 108363 471064
rect 99790 471006 108363 471008
rect 99790 470764 99850 471006
rect 108297 471003 108363 471006
rect 67541 470250 67607 470253
rect 102777 470250 102843 470253
rect 67541 470248 70226 470250
rect 67541 470192 67546 470248
rect 67602 470192 70226 470248
rect 67541 470190 70226 470192
rect 67541 470187 67607 470190
rect 70166 470084 70226 470190
rect 99790 470248 102843 470250
rect 99790 470192 102782 470248
rect 102838 470192 102843 470248
rect 99790 470190 102843 470192
rect 99790 470084 99850 470190
rect 102777 470187 102843 470190
rect 67633 469706 67699 469709
rect 67633 469704 70226 469706
rect 67633 469648 67638 469704
rect 67694 469648 70226 469704
rect 67633 469646 70226 469648
rect 67633 469643 67699 469646
rect 70166 469404 70226 469646
rect 102225 469570 102291 469573
rect 99790 469568 102291 469570
rect 99790 469512 102230 469568
rect 102286 469512 102291 469568
rect 99790 469510 102291 469512
rect 99790 469404 99850 469510
rect 102225 469507 102291 469510
rect 60457 469162 60523 469165
rect 60457 469160 64890 469162
rect 60457 469104 60462 469160
rect 60518 469104 64890 469160
rect 60457 469102 64890 469104
rect 60457 469099 60523 469102
rect 64830 469026 64890 469102
rect 103513 469026 103579 469029
rect 64830 468966 70226 469026
rect 70166 468724 70226 468966
rect 99790 469024 103579 469026
rect 99790 468968 103518 469024
rect 103574 468968 103579 469024
rect 99790 468966 103579 468968
rect 99790 468724 99850 468966
rect 103513 468963 103579 468966
rect 104750 468420 104756 468484
rect 104820 468482 104826 468484
rect 132769 468482 132835 468485
rect 151997 468482 152063 468485
rect 104820 468480 152063 468482
rect 104820 468424 132774 468480
rect 132830 468424 152002 468480
rect 152058 468424 152063 468480
rect 104820 468422 152063 468424
rect 104820 468420 104826 468422
rect 132769 468419 132835 468422
rect 151997 468419 152063 468422
rect 67633 468210 67699 468213
rect 67633 468208 70226 468210
rect 67633 468152 67638 468208
rect 67694 468152 70226 468208
rect 67633 468150 70226 468152
rect 67633 468147 67699 468150
rect 70166 468044 70226 468150
rect 59118 467876 59124 467940
rect 59188 467938 59194 467940
rect 60457 467938 60523 467941
rect 59188 467936 60523 467938
rect 59188 467880 60462 467936
rect 60518 467880 60523 467936
rect 59188 467878 60523 467880
rect 59188 467876 59194 467878
rect 60457 467875 60523 467878
rect 67633 466850 67699 466853
rect 99790 466850 99850 467228
rect 102225 466850 102291 466853
rect 67633 466848 70226 466850
rect 67633 466792 67638 466848
rect 67694 466792 70226 466848
rect 67633 466790 70226 466792
rect 99790 466848 102291 466850
rect 99790 466792 102230 466848
rect 102286 466792 102291 466848
rect 99790 466790 102291 466792
rect 67633 466787 67699 466790
rect 70166 466684 70226 466790
rect 102225 466787 102291 466790
rect 104750 466578 104756 466580
rect 64454 466380 64460 466444
rect 64524 466442 64530 466444
rect 67265 466442 67331 466445
rect 67449 466442 67515 466445
rect 64524 466440 67515 466442
rect 64524 466384 67270 466440
rect 67326 466384 67454 466440
rect 67510 466384 67515 466440
rect 64524 466382 67515 466384
rect 64524 466380 64530 466382
rect 67265 466379 67331 466382
rect 67449 466379 67515 466382
rect 99606 466306 99666 466548
rect 100158 466518 104756 466578
rect 100158 466306 100218 466518
rect 104750 466516 104756 466518
rect 104820 466516 104826 466580
rect 99606 466246 100218 466306
rect 64822 466108 64828 466172
rect 64892 466170 64898 466172
rect 65609 466170 65675 466173
rect 64892 466168 65675 466170
rect 64892 466112 65614 466168
rect 65670 466112 65675 466168
rect 64892 466110 65675 466112
rect 64892 466108 64898 466110
rect 65609 466107 65675 466110
rect 67633 466170 67699 466173
rect 102225 466170 102291 466173
rect 67633 466168 70226 466170
rect 67633 466112 67638 466168
rect 67694 466112 70226 466168
rect 67633 466110 70226 466112
rect 67633 466107 67699 466110
rect 70166 466004 70226 466110
rect 99790 466168 102291 466170
rect 99790 466112 102230 466168
rect 102286 466112 102291 466168
rect 99790 466110 102291 466112
rect 99790 466004 99850 466110
rect 102225 466107 102291 466110
rect 108481 465762 108547 465765
rect 110638 465762 110644 465764
rect 108481 465760 110644 465762
rect 108481 465704 108486 465760
rect 108542 465704 110644 465760
rect 108481 465702 110644 465704
rect 108481 465699 108547 465702
rect 110638 465700 110644 465702
rect 110708 465700 110714 465764
rect 67449 465626 67515 465629
rect 67449 465624 70410 465626
rect 67449 465568 67454 465624
rect 67510 465568 70410 465624
rect 67449 465566 70410 465568
rect 67449 465563 67515 465566
rect 70350 465324 70410 465566
rect 102317 465490 102383 465493
rect 99790 465488 102383 465490
rect 99790 465432 102322 465488
rect 102378 465432 102383 465488
rect 99790 465430 102383 465432
rect 99790 465324 99850 465430
rect 102317 465427 102383 465430
rect 103513 464946 103579 464949
rect 99790 464944 103579 464946
rect 99790 464888 103518 464944
rect 103574 464888 103579 464944
rect 99790 464886 103579 464888
rect 67633 464810 67699 464813
rect 67633 464808 70226 464810
rect 67633 464752 67638 464808
rect 67694 464752 70226 464808
rect 67633 464750 70226 464752
rect 67633 464747 67699 464750
rect 70166 464644 70226 464750
rect 99790 464644 99850 464886
rect 103513 464883 103579 464886
rect 67725 464266 67791 464269
rect 67725 464264 70410 464266
rect 67725 464208 67730 464264
rect 67786 464208 70410 464264
rect 67725 464206 70410 464208
rect 67725 464203 67791 464206
rect 70350 463964 70410 464206
rect 104014 464130 104020 464132
rect 99790 464070 104020 464130
rect 99790 463964 99850 464070
rect 104014 464068 104020 464070
rect 104084 464130 104090 464132
rect 104709 464130 104775 464133
rect 104084 464128 104775 464130
rect 104084 464072 104714 464128
rect 104770 464072 104775 464128
rect 104084 464070 104775 464072
rect 104084 464068 104090 464070
rect 104709 464067 104775 464070
rect 67633 462906 67699 462909
rect 70350 462906 70410 463148
rect 67633 462904 70410 462906
rect 67633 462848 67638 462904
rect 67694 462848 70410 462904
rect 67633 462846 70410 462848
rect 99606 462906 99666 463148
rect 102225 462906 102291 462909
rect 99606 462904 102291 462906
rect 99606 462848 102230 462904
rect 102286 462848 102291 462904
rect 99606 462846 102291 462848
rect 67633 462843 67699 462846
rect 102225 462843 102291 462846
rect 67633 462770 67699 462773
rect 67633 462768 70226 462770
rect -960 462634 480 462724
rect 67633 462712 67638 462768
rect 67694 462712 70226 462768
rect 67633 462710 70226 462712
rect 67633 462707 67699 462710
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect 70166 462604 70226 462710
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 106641 462226 106707 462229
rect 106774 462226 106780 462228
rect 106641 462224 106780 462226
rect 106641 462168 106646 462224
rect 106702 462168 106780 462224
rect 106641 462166 106780 462168
rect 106641 462163 106707 462166
rect 106774 462164 106780 462166
rect 106844 462164 106850 462228
rect 102225 462090 102291 462093
rect 99790 462088 102291 462090
rect 99790 462032 102230 462088
rect 102286 462032 102291 462088
rect 99790 462030 102291 462032
rect 99790 461924 99850 462030
rect 102225 462027 102291 462030
rect 102317 461546 102383 461549
rect 99790 461544 102383 461546
rect 99790 461488 102322 461544
rect 102378 461488 102383 461544
rect 99790 461486 102383 461488
rect 67633 461410 67699 461413
rect 67633 461408 70226 461410
rect 67633 461352 67638 461408
rect 67694 461352 70226 461408
rect 67633 461350 70226 461352
rect 67633 461347 67699 461350
rect 70166 461244 70226 461350
rect 99790 461244 99850 461486
rect 102317 461483 102383 461486
rect 130377 461138 130443 461141
rect 133822 461138 133828 461140
rect 130377 461136 133828 461138
rect 130377 461080 130382 461136
rect 130438 461080 133828 461136
rect 130377 461078 133828 461080
rect 130377 461075 130443 461078
rect 133822 461076 133828 461078
rect 133892 461076 133898 461140
rect 106641 461002 106707 461005
rect 138013 461002 138079 461005
rect 106641 461000 138079 461002
rect 106641 460944 106646 461000
rect 106702 460944 138018 461000
rect 138074 460944 138079 461000
rect 106641 460942 138079 460944
rect 106641 460939 106707 460942
rect 138013 460939 138079 460942
rect 64689 460866 64755 460869
rect 64822 460866 64828 460868
rect 64689 460864 64828 460866
rect 64689 460808 64694 460864
rect 64750 460808 64828 460864
rect 64689 460806 64828 460808
rect 64689 460803 64755 460806
rect 64822 460804 64828 460806
rect 64892 460804 64898 460868
rect 67633 460730 67699 460733
rect 102133 460730 102199 460733
rect 67633 460728 70226 460730
rect 67633 460672 67638 460728
rect 67694 460672 70226 460728
rect 67633 460670 70226 460672
rect 67633 460667 67699 460670
rect 70166 460564 70226 460670
rect 99790 460728 102199 460730
rect 99790 460672 102138 460728
rect 102194 460672 102199 460728
rect 99790 460670 102199 460672
rect 99790 460564 99850 460670
rect 102133 460667 102199 460670
rect 67725 460186 67791 460189
rect 102317 460186 102383 460189
rect 67725 460184 70226 460186
rect 67725 460128 67730 460184
rect 67786 460128 70226 460184
rect 67725 460126 70226 460128
rect 67725 460123 67791 460126
rect 70166 459884 70226 460126
rect 99790 460184 102383 460186
rect 99790 460128 102322 460184
rect 102378 460128 102383 460184
rect 99790 460126 102383 460128
rect 99790 459884 99850 460126
rect 102317 460123 102383 460126
rect 67633 459370 67699 459373
rect 102133 459370 102199 459373
rect 67633 459368 70226 459370
rect 67633 459312 67638 459368
rect 67694 459312 70226 459368
rect 67633 459310 70226 459312
rect 67633 459307 67699 459310
rect 70166 459204 70226 459310
rect 99790 459368 102199 459370
rect 99790 459312 102138 459368
rect 102194 459312 102199 459368
rect 99790 459310 102199 459312
rect 99790 459204 99850 459310
rect 102133 459307 102199 459310
rect 32949 458826 33015 458829
rect 62982 458826 62988 458828
rect 32949 458824 62988 458826
rect 32949 458768 32954 458824
rect 33010 458768 62988 458824
rect 32949 458766 62988 458768
rect 32949 458763 33015 458766
rect 62982 458764 62988 458766
rect 63052 458826 63058 458828
rect 63052 458766 70226 458826
rect 63052 458764 63058 458766
rect 70166 458524 70226 458766
rect 102133 458690 102199 458693
rect 99790 458688 102199 458690
rect 99790 458632 102138 458688
rect 102194 458632 102199 458688
rect 99790 458630 102199 458632
rect 99790 458524 99850 458630
rect 102133 458627 102199 458630
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 102317 458010 102383 458013
rect 99790 458008 102383 458010
rect 99790 457952 102322 458008
rect 102378 457952 102383 458008
rect 583520 457996 584960 458086
rect 99790 457950 102383 457952
rect 99790 457844 99850 457950
rect 102317 457947 102383 457950
rect 67725 457330 67791 457333
rect 70166 457330 70226 457708
rect 67725 457328 70226 457330
rect 67725 457272 67730 457328
rect 67786 457272 70226 457328
rect 67725 457270 70226 457272
rect 67725 457267 67791 457270
rect 67633 456922 67699 456925
rect 67633 456920 69858 456922
rect 67633 456864 67638 456920
rect 67694 456864 69858 456920
rect 67633 456862 69858 456864
rect 67633 456859 67699 456862
rect 69798 456786 69858 456862
rect 70350 456786 70410 457028
rect 69798 456726 70410 456786
rect 102133 456650 102199 456653
rect 99790 456648 102199 456650
rect 99790 456592 102138 456648
rect 102194 456592 102199 456648
rect 99790 456590 102199 456592
rect 99790 456484 99850 456590
rect 102133 456587 102199 456590
rect 103513 456106 103579 456109
rect 99790 456104 103579 456106
rect 99790 456048 103518 456104
rect 103574 456048 103579 456104
rect 99790 456046 103579 456048
rect 67633 455970 67699 455973
rect 67633 455968 70226 455970
rect 67633 455912 67638 455968
rect 67694 455912 70226 455968
rect 67633 455910 70226 455912
rect 67633 455907 67699 455910
rect 70166 455804 70226 455910
rect 99790 455804 99850 456046
rect 103513 456043 103579 456046
rect 42701 454746 42767 454749
rect 67633 454746 67699 454749
rect 70166 454746 70226 454988
rect 42701 454744 64890 454746
rect 42701 454688 42706 454744
rect 42762 454688 64890 454744
rect 42701 454686 64890 454688
rect 42701 454683 42767 454686
rect 64830 454610 64890 454686
rect 67633 454744 70226 454746
rect 67633 454688 67638 454744
rect 67694 454688 70226 454744
rect 67633 454686 70226 454688
rect 99790 454746 99850 454988
rect 102133 454746 102199 454749
rect 99790 454744 102199 454746
rect 99790 454688 102138 454744
rect 102194 454688 102199 454744
rect 99790 454686 102199 454688
rect 67633 454683 67699 454686
rect 102133 454683 102199 454686
rect 68870 454610 68876 454612
rect 64830 454550 68876 454610
rect 68870 454548 68876 454550
rect 68940 454610 68946 454612
rect 102869 454610 102935 454613
rect 103329 454610 103395 454613
rect 68940 454550 70226 454610
rect 68940 454548 68946 454550
rect 70166 454444 70226 454550
rect 99790 454608 103395 454610
rect 99790 454552 102874 454608
rect 102930 454552 103334 454608
rect 103390 454552 103395 454608
rect 99790 454550 103395 454552
rect 99790 454444 99850 454550
rect 102869 454547 102935 454550
rect 103329 454547 103395 454550
rect 118969 454066 119035 454069
rect 119337 454066 119403 454069
rect 129774 454066 129780 454068
rect 118969 454064 129780 454066
rect 118969 454008 118974 454064
rect 119030 454008 119342 454064
rect 119398 454008 129780 454064
rect 118969 454006 129780 454008
rect 118969 454003 119035 454006
rect 119337 454003 119403 454006
rect 129774 454004 129780 454006
rect 129844 454004 129850 454068
rect 57697 453932 57763 453933
rect 57646 453930 57652 453932
rect 57606 453870 57652 453930
rect 57716 453928 57763 453932
rect 102133 453930 102199 453933
rect 57758 453872 57763 453928
rect 57646 453868 57652 453870
rect 57716 453868 57763 453872
rect 57697 453867 57763 453868
rect 99790 453928 102199 453930
rect 99790 453872 102138 453928
rect 102194 453872 102199 453928
rect 99790 453870 102199 453872
rect 99790 453764 99850 453870
rect 102133 453867 102199 453870
rect 67633 453386 67699 453389
rect 70350 453386 70410 453628
rect 102317 453386 102383 453389
rect 67633 453384 70410 453386
rect 67633 453328 67638 453384
rect 67694 453328 70410 453384
rect 67633 453326 70410 453328
rect 99790 453384 102383 453386
rect 99790 453328 102322 453384
rect 102378 453328 102383 453384
rect 99790 453326 102383 453328
rect 67633 453323 67699 453326
rect 67725 453250 67791 453253
rect 67725 453248 70226 453250
rect 67725 453192 67730 453248
rect 67786 453192 70226 453248
rect 67725 453190 70226 453192
rect 67725 453187 67791 453190
rect 70166 453084 70226 453190
rect 99790 453084 99850 453326
rect 102317 453323 102383 453326
rect 69054 451964 69060 452028
rect 69124 452026 69130 452028
rect 70166 452026 70226 452268
rect 69124 451966 70226 452026
rect 99790 452026 99850 452268
rect 102133 452026 102199 452029
rect 115933 452028 115999 452029
rect 115933 452026 115980 452028
rect 99790 452024 102199 452026
rect 99790 451968 102138 452024
rect 102194 451968 102199 452024
rect 99790 451966 102199 451968
rect 115888 452024 115980 452026
rect 115888 451968 115938 452024
rect 115888 451966 115980 451968
rect 69124 451964 69130 451966
rect 102133 451963 102199 451966
rect 115933 451964 115980 451966
rect 116044 451964 116050 452028
rect 115933 451963 115999 451964
rect 68921 451890 68987 451893
rect 68921 451888 70226 451890
rect 68921 451832 68926 451888
rect 68982 451832 70226 451888
rect 68921 451830 70226 451832
rect 68921 451827 68987 451830
rect 70166 451724 70226 451830
rect 64689 451482 64755 451485
rect 64822 451482 64828 451484
rect 64689 451480 64828 451482
rect 64689 451424 64694 451480
rect 64750 451424 64828 451480
rect 64689 451422 64828 451424
rect 64689 451419 64755 451422
rect 64822 451420 64828 451422
rect 64892 451420 64898 451484
rect 69054 451346 69060 451348
rect 62622 451286 69060 451346
rect 35709 451210 35775 451213
rect 62622 451212 62682 451286
rect 69054 451284 69060 451286
rect 69124 451284 69130 451348
rect 108982 451284 108988 451348
rect 109052 451346 109058 451348
rect 149145 451346 149211 451349
rect 109052 451344 149211 451346
rect 109052 451288 149150 451344
rect 149206 451288 149211 451344
rect 109052 451286 149211 451288
rect 109052 451284 109058 451286
rect 149145 451283 149211 451286
rect 64781 451212 64847 451213
rect 62614 451210 62620 451212
rect 35709 451208 62620 451210
rect 35709 451152 35714 451208
rect 35770 451152 62620 451208
rect 35709 451150 62620 451152
rect 35709 451147 35775 451150
rect 62614 451148 62620 451150
rect 62684 451148 62690 451212
rect 64781 451210 64828 451212
rect 64736 451208 64828 451210
rect 64892 451210 64898 451212
rect 101949 451210 102015 451213
rect 64736 451152 64786 451208
rect 64736 451150 64828 451152
rect 64781 451148 64828 451150
rect 64892 451150 64974 451210
rect 99790 451208 102015 451210
rect 99790 451152 101954 451208
rect 102010 451152 102015 451208
rect 99790 451150 102015 451152
rect 64892 451148 64898 451150
rect 64781 451147 64847 451148
rect 99790 451044 99850 451150
rect 101949 451147 102015 451150
rect 102501 450666 102567 450669
rect 99790 450664 102567 450666
rect 99790 450608 102506 450664
rect 102562 450608 102567 450664
rect 99790 450606 102567 450608
rect 99790 450364 99850 450606
rect 102501 450603 102567 450606
rect 105353 450530 105419 450533
rect 108982 450530 108988 450532
rect 105353 450528 108988 450530
rect 105353 450472 105358 450528
rect 105414 450472 108988 450528
rect 105353 450470 108988 450472
rect 105353 450467 105419 450470
rect 108982 450468 108988 450470
rect 109052 450468 109058 450532
rect 68134 450122 68140 450124
rect 64830 450062 68140 450122
rect 49417 449986 49483 449989
rect 64830 449986 64890 450062
rect 68134 450060 68140 450062
rect 68204 450060 68210 450124
rect 49417 449984 64890 449986
rect 49417 449928 49422 449984
rect 49478 449928 64890 449984
rect 49417 449926 64890 449928
rect 67633 449986 67699 449989
rect 70166 449986 70226 450228
rect 67633 449984 70226 449986
rect 67633 449928 67638 449984
rect 67694 449928 70226 449984
rect 67633 449926 70226 449928
rect 49417 449923 49483 449926
rect 67633 449923 67699 449926
rect 102133 449850 102199 449853
rect 99790 449848 102199 449850
rect 99790 449792 102138 449848
rect 102194 449792 102199 449848
rect 99790 449790 102199 449792
rect 99790 449684 99850 449790
rect 102133 449787 102199 449790
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 67633 449170 67699 449173
rect 70166 449170 70226 449548
rect 102317 449306 102383 449309
rect 67633 449168 70226 449170
rect 67633 449112 67638 449168
rect 67694 449112 70226 449168
rect 67633 449110 70226 449112
rect 99790 449304 102383 449306
rect 99790 449248 102322 449304
rect 102378 449248 102383 449304
rect 99790 449246 102383 449248
rect 67633 449107 67699 449110
rect 99790 449004 99850 449246
rect 102317 449243 102383 449246
rect 68134 448564 68140 448628
rect 68204 448626 68210 448628
rect 70350 448626 70410 448868
rect 68204 448566 70410 448626
rect 68204 448564 68210 448566
rect 67633 447810 67699 447813
rect 70166 447810 70226 448188
rect 99606 447946 99666 448188
rect 102317 447946 102383 447949
rect 99606 447944 102383 447946
rect 99606 447888 102322 447944
rect 102378 447888 102383 447944
rect 99606 447886 102383 447888
rect 102317 447883 102383 447886
rect 102133 447810 102199 447813
rect 67633 447808 70226 447810
rect 67633 447752 67638 447808
rect 67694 447752 70226 447808
rect 67633 447750 70226 447752
rect 99790 447808 102199 447810
rect 99790 447752 102138 447808
rect 102194 447752 102199 447808
rect 99790 447750 102199 447752
rect 67633 447747 67699 447750
rect 99790 447644 99850 447750
rect 102133 447747 102199 447750
rect 61878 447340 61884 447404
rect 61948 447402 61954 447404
rect 63217 447402 63283 447405
rect 61948 447400 64890 447402
rect 61948 447344 63222 447400
rect 63278 447344 64890 447400
rect 61948 447342 64890 447344
rect 61948 447340 61954 447342
rect 63217 447339 63283 447342
rect 64830 447266 64890 447342
rect 70350 447266 70410 447508
rect 64830 447206 70410 447266
rect 105721 447266 105787 447269
rect 111926 447266 111932 447268
rect 105721 447264 111932 447266
rect 105721 447208 105726 447264
rect 105782 447208 111932 447264
rect 105721 447206 111932 447208
rect 105721 447203 105787 447206
rect 111926 447204 111932 447206
rect 111996 447204 112002 447268
rect 64781 447132 64847 447133
rect 64781 447128 64828 447132
rect 64892 447130 64898 447132
rect 64781 447072 64786 447128
rect 64781 447068 64828 447072
rect 64892 447070 64938 447130
rect 64892 447068 64898 447070
rect 64781 447067 64847 447068
rect 67633 446586 67699 446589
rect 70166 446586 70226 446828
rect 67633 446584 70226 446586
rect 67633 446528 67638 446584
rect 67694 446528 70226 446584
rect 67633 446526 70226 446528
rect 99606 446586 99666 446828
rect 101029 446586 101095 446589
rect 99606 446584 101095 446586
rect 99606 446528 101034 446584
rect 101090 446528 101095 446584
rect 99606 446526 101095 446528
rect 67633 446523 67699 446526
rect 101029 446523 101095 446526
rect 48129 446450 48195 446453
rect 66662 446450 66668 446452
rect 48129 446448 66668 446450
rect 48129 446392 48134 446448
rect 48190 446392 66668 446448
rect 48129 446390 66668 446392
rect 48129 446387 48195 446390
rect 66662 446388 66668 446390
rect 66732 446450 66738 446452
rect 66732 446390 70226 446450
rect 66732 446388 66738 446390
rect 70166 446284 70226 446390
rect 61745 445772 61811 445773
rect 61694 445770 61700 445772
rect 61654 445710 61700 445770
rect 61764 445768 61811 445772
rect 102317 445770 102383 445773
rect 61806 445712 61811 445768
rect 61694 445708 61700 445710
rect 61764 445708 61811 445712
rect 61745 445707 61811 445708
rect 99790 445768 102383 445770
rect 99790 445712 102322 445768
rect 102378 445712 102383 445768
rect 99790 445710 102383 445712
rect 99790 445604 99850 445710
rect 102317 445707 102383 445710
rect 102133 445226 102199 445229
rect 99790 445224 102199 445226
rect 99790 445168 102138 445224
rect 102194 445168 102199 445224
rect 99790 445166 102199 445168
rect 67633 445090 67699 445093
rect 68737 445090 68803 445093
rect 67633 445088 70226 445090
rect 67633 445032 67638 445088
rect 67694 445032 68742 445088
rect 68798 445032 70226 445088
rect 67633 445030 70226 445032
rect 67633 445027 67699 445030
rect 68737 445027 68803 445030
rect 70166 444924 70226 445030
rect 99790 444924 99850 445166
rect 102133 445163 102199 445166
rect 128537 445090 128603 445093
rect 128854 445090 128860 445092
rect 128537 445088 128860 445090
rect 128537 445032 128542 445088
rect 128598 445032 128860 445088
rect 128537 445030 128860 445032
rect 128537 445027 128603 445030
rect 128854 445028 128860 445030
rect 128924 445028 128930 445092
rect 583520 444668 584960 444908
rect 67633 443866 67699 443869
rect 68277 443866 68343 443869
rect 70350 443866 70410 444108
rect 67633 443864 70410 443866
rect 67633 443808 67638 443864
rect 67694 443808 68282 443864
rect 68338 443808 70410 443864
rect 67633 443806 70410 443808
rect 99606 443866 99666 444108
rect 102317 443866 102383 443869
rect 99606 443864 102383 443866
rect 99606 443808 102322 443864
rect 102378 443808 102383 443864
rect 99606 443806 102383 443808
rect 67633 443803 67699 443806
rect 68277 443803 68343 443806
rect 102317 443803 102383 443806
rect 99373 443730 99439 443733
rect 102133 443730 102199 443733
rect 99373 443728 102199 443730
rect 99373 443672 99378 443728
rect 99434 443672 102138 443728
rect 102194 443672 102199 443728
rect 99373 443670 102199 443672
rect 99373 443667 99439 443670
rect 99790 443564 99850 443670
rect 102133 443667 102199 443670
rect 66253 443050 66319 443053
rect 66662 443050 66668 443052
rect 66253 443048 66668 443050
rect 66253 442992 66258 443048
rect 66314 442992 66668 443048
rect 66253 442990 66668 442992
rect 66253 442987 66319 442990
rect 66662 442988 66668 442990
rect 66732 443050 66738 443052
rect 70166 443050 70226 443428
rect 66732 442990 70226 443050
rect 66732 442988 66738 442990
rect 67725 442778 67791 442781
rect 67725 442776 70380 442778
rect 67725 442720 67730 442776
rect 67786 442720 70380 442776
rect 67725 442718 70380 442720
rect 67725 442715 67791 442718
rect 58566 442444 58572 442508
rect 58636 442506 58642 442508
rect 58636 442446 60750 442506
rect 58636 442444 58642 442446
rect 60690 442370 60750 442446
rect 70342 442370 70348 442372
rect 60690 442310 70348 442370
rect 70342 442308 70348 442310
rect 70412 442308 70418 442372
rect 99790 442370 99850 442748
rect 99925 442506 99991 442509
rect 113173 442506 113239 442509
rect 99925 442504 113239 442506
rect 99925 442448 99930 442504
rect 99986 442448 113178 442504
rect 113234 442448 113239 442504
rect 99925 442446 113239 442448
rect 99925 442443 99991 442446
rect 113173 442443 113239 442446
rect 102133 442370 102199 442373
rect 99790 442368 102199 442370
rect 99790 442312 102138 442368
rect 102194 442312 102199 442368
rect 99790 442310 102199 442312
rect 102133 442307 102199 442310
rect 120022 442234 120028 442236
rect 103470 442174 120028 442234
rect 67633 441826 67699 441829
rect 70350 441826 70410 442068
rect 67633 441824 70410 441826
rect 67633 441768 67638 441824
rect 67694 441768 70410 441824
rect 67633 441766 70410 441768
rect 99606 441826 99666 442068
rect 101990 441900 101996 441964
rect 102060 441962 102066 441964
rect 103470 441962 103530 442174
rect 120022 442172 120028 442174
rect 120092 442172 120098 442236
rect 102060 441902 103530 441962
rect 102060 441900 102066 441902
rect 101998 441826 102058 441900
rect 99606 441766 102058 441826
rect 67633 441763 67699 441766
rect 67633 441146 67699 441149
rect 70350 441146 70410 441388
rect 67633 441144 70410 441146
rect 67633 441088 67638 441144
rect 67694 441088 70410 441144
rect 67633 441086 70410 441088
rect 99606 441146 99666 441388
rect 100753 441146 100819 441149
rect 99606 441144 100819 441146
rect 99606 441088 100758 441144
rect 100814 441088 100819 441144
rect 99606 441086 100819 441088
rect 67633 441083 67699 441086
rect 100753 441083 100819 441086
rect 67633 441010 67699 441013
rect 67633 441008 70226 441010
rect 67633 440952 67638 441008
rect 67694 440952 70226 441008
rect 67633 440950 70226 440952
rect 67633 440947 67699 440950
rect 70166 440844 70226 440950
rect 99790 440194 100034 440228
rect 100845 440194 100911 440197
rect 99790 440192 100911 440194
rect 99790 440168 100850 440192
rect 99790 440164 99850 440168
rect 99974 440136 100850 440168
rect 100906 440136 100911 440192
rect 99974 440134 100911 440136
rect 100845 440131 100911 440134
rect 121637 439514 121703 439517
rect 122097 439514 122163 439517
rect 125726 439514 125732 439516
rect 121637 439512 125732 439514
rect 121637 439456 121642 439512
rect 121698 439456 122102 439512
rect 122158 439456 125732 439512
rect 121637 439454 125732 439456
rect 121637 439451 121703 439454
rect 122097 439451 122163 439454
rect 125726 439452 125732 439454
rect 125796 439452 125802 439516
rect 65926 438908 65932 438972
rect 65996 438970 66002 438972
rect 71037 438970 71103 438973
rect 65996 438968 71103 438970
rect 65996 438912 71042 438968
rect 71098 438912 71103 438968
rect 65996 438910 71103 438912
rect 65996 438908 66002 438910
rect 71037 438907 71103 438910
rect 99649 438970 99715 438973
rect 120349 438970 120415 438973
rect 121678 438970 121684 438972
rect 99649 438968 121684 438970
rect 99649 438912 99654 438968
rect 99710 438912 120354 438968
rect 120410 438912 121684 438968
rect 99649 438910 121684 438912
rect 99649 438907 99715 438910
rect 120349 438907 120415 438910
rect 121678 438908 121684 438910
rect 121748 438908 121754 438972
rect 84193 438698 84259 438701
rect 84837 438698 84903 438701
rect 111742 438698 111748 438700
rect 84193 438696 111748 438698
rect 84193 438640 84198 438696
rect 84254 438640 84842 438696
rect 84898 438640 111748 438696
rect 84193 438638 111748 438640
rect 84193 438635 84259 438638
rect 84837 438635 84903 438638
rect 111742 438636 111748 438638
rect 111812 438636 111818 438700
rect 57881 438154 57947 438157
rect 75177 438154 75243 438157
rect 57881 438152 75243 438154
rect 57881 438096 57886 438152
rect 57942 438096 75182 438152
rect 75238 438096 75243 438152
rect 57881 438094 75243 438096
rect 57881 438091 57947 438094
rect 75177 438091 75243 438094
rect 97073 437882 97139 437885
rect 98494 437882 98500 437884
rect 97073 437880 98500 437882
rect 97073 437824 97078 437880
rect 97134 437824 98500 437880
rect 97073 437822 98500 437824
rect 97073 437819 97139 437822
rect 98494 437820 98500 437822
rect 98564 437820 98570 437884
rect 64413 437610 64479 437613
rect 64822 437610 64828 437612
rect 64413 437608 64828 437610
rect 64413 437552 64418 437608
rect 64474 437552 64828 437608
rect 64413 437550 64828 437552
rect 64413 437547 64479 437550
rect 64822 437548 64828 437550
rect 64892 437548 64898 437612
rect 57830 437412 57836 437476
rect 57900 437474 57906 437476
rect 84193 437474 84259 437477
rect 85021 437474 85087 437477
rect 57900 437472 85087 437474
rect 57900 437416 84198 437472
rect 84254 437416 85026 437472
rect 85082 437416 85087 437472
rect 57900 437414 85087 437416
rect 57900 437412 57906 437414
rect 84193 437411 84259 437414
rect 85021 437411 85087 437414
rect -960 436508 480 436748
rect 69105 436522 69171 436525
rect 69238 436522 69244 436524
rect 69105 436520 69244 436522
rect 69105 436464 69110 436520
rect 69166 436464 69244 436520
rect 69105 436462 69244 436464
rect 69105 436459 69171 436462
rect 69238 436460 69244 436462
rect 69308 436460 69314 436524
rect 70393 436116 70459 436117
rect 70342 436114 70348 436116
rect 70302 436054 70348 436114
rect 70412 436112 70459 436116
rect 70454 436056 70459 436112
rect 70342 436052 70348 436054
rect 70412 436052 70459 436056
rect 70393 436051 70459 436052
rect 48078 434556 48084 434620
rect 48148 434618 48154 434620
rect 77293 434618 77359 434621
rect 48148 434616 77359 434618
rect 48148 434560 77298 434616
rect 77354 434560 77359 434616
rect 48148 434558 77359 434560
rect 48148 434556 48154 434558
rect 77293 434555 77359 434558
rect 64413 432034 64479 432037
rect 64822 432034 64828 432036
rect 64413 432032 64828 432034
rect 64413 431976 64418 432032
rect 64474 431976 64828 432032
rect 64413 431974 64828 431976
rect 64413 431971 64479 431974
rect 64822 431972 64828 431974
rect 64892 431972 64898 432036
rect 64505 431898 64571 431901
rect 64822 431898 64828 431900
rect 64505 431896 64828 431898
rect 64505 431840 64510 431896
rect 64566 431840 64828 431896
rect 64505 431838 64828 431840
rect 64505 431835 64571 431838
rect 64822 431836 64828 431838
rect 64892 431836 64898 431900
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect 69054 428436 69060 428500
rect 69124 428498 69130 428500
rect 580257 428498 580323 428501
rect 69124 428496 580323 428498
rect 69124 428440 580262 428496
rect 580318 428440 580323 428496
rect 69124 428438 580323 428440
rect 69124 428436 69130 428438
rect 580257 428435 580323 428438
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 64505 422378 64571 422381
rect 64822 422378 64828 422380
rect 64505 422376 64828 422378
rect 64505 422320 64510 422376
rect 64566 422320 64828 422376
rect 64505 422318 64828 422320
rect 64505 422315 64571 422318
rect 64822 422316 64828 422318
rect 64892 422316 64898 422380
rect 580257 418298 580323 418301
rect 583520 418298 584960 418388
rect 580257 418296 584960 418298
rect 580257 418240 580262 418296
rect 580318 418240 584960 418296
rect 580257 418238 584960 418240
rect 580257 418235 580323 418238
rect 583520 418148 584960 418238
rect 64505 412586 64571 412589
rect 64822 412586 64828 412588
rect 64505 412584 64828 412586
rect 64505 412528 64510 412584
rect 64566 412528 64828 412584
rect 64505 412526 64828 412528
rect 64505 412523 64571 412526
rect 64822 412524 64828 412526
rect 64892 412524 64898 412588
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 58985 407010 59051 407013
rect 59118 407010 59124 407012
rect 58985 407008 59124 407010
rect 58985 406952 58990 407008
rect 59046 406952 59124 407008
rect 58985 406950 59124 406952
rect 58985 406947 59051 406950
rect 59118 406948 59124 406950
rect 59188 406948 59194 407012
rect 58985 405786 59051 405789
rect 335997 405786 336063 405789
rect 58985 405784 336063 405786
rect 58985 405728 58990 405784
rect 59046 405728 336002 405784
rect 336058 405728 336063 405784
rect 58985 405726 336063 405728
rect 58985 405723 59051 405726
rect 335997 405723 336063 405726
rect 579613 404970 579679 404973
rect 583520 404970 584960 405060
rect 579613 404968 584960 404970
rect 579613 404912 579618 404968
rect 579674 404912 584960 404968
rect 579613 404910 584960 404912
rect 579613 404907 579679 404910
rect 583520 404820 584960 404910
rect 64505 403066 64571 403069
rect 64822 403066 64828 403068
rect 64505 403064 64828 403066
rect 64505 403008 64510 403064
rect 64566 403008 64828 403064
rect 64505 403006 64828 403008
rect 64505 403003 64571 403006
rect 64822 403004 64828 403006
rect 64892 403004 64898 403068
rect 61510 402188 61516 402252
rect 61580 402250 61586 402252
rect 61580 402190 64890 402250
rect 61580 402188 61586 402190
rect 64830 401706 64890 402190
rect 68829 401706 68895 401709
rect 338113 401706 338179 401709
rect 64830 401704 338179 401706
rect 64830 401648 68834 401704
rect 68890 401648 338118 401704
rect 338174 401648 338179 401704
rect 64830 401646 338179 401648
rect 68829 401643 68895 401646
rect 338113 401643 338179 401646
rect 94497 401026 94563 401029
rect 121862 401026 121868 401028
rect 94497 401024 121868 401026
rect 94497 400968 94502 401024
rect 94558 400968 121868 401024
rect 94497 400966 121868 400968
rect 94497 400963 94563 400966
rect 121862 400964 121868 400966
rect 121932 400964 121938 401028
rect 98494 400828 98500 400892
rect 98564 400890 98570 400892
rect 132769 400890 132835 400893
rect 98564 400888 132835 400890
rect 98564 400832 132774 400888
rect 132830 400832 132835 400888
rect 98564 400830 132835 400832
rect 98564 400828 98570 400830
rect 132769 400827 132835 400830
rect 64505 400348 64571 400349
rect 64454 400346 64460 400348
rect 64378 400286 64460 400346
rect 64524 400346 64571 400348
rect 166257 400346 166323 400349
rect 64524 400344 166323 400346
rect 64566 400288 166262 400344
rect 166318 400288 166323 400344
rect 64454 400284 64460 400286
rect 64524 400286 166323 400288
rect 64524 400284 64571 400286
rect 64505 400283 64571 400284
rect 166257 400283 166323 400286
rect 104014 397972 104020 398036
rect 104084 398034 104090 398036
rect 117497 398034 117563 398037
rect 104084 398032 117563 398034
rect 104084 397976 117502 398032
rect 117558 397976 117563 398032
rect 104084 397974 117563 397976
rect 104084 397972 104090 397974
rect 117497 397971 117563 397974
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 106917 395314 106983 395317
rect 118734 395314 118740 395316
rect 106917 395312 118740 395314
rect 106917 395256 106922 395312
rect 106978 395256 118740 395312
rect 106917 395254 118740 395256
rect 106917 395251 106983 395254
rect 118734 395252 118740 395254
rect 118804 395252 118810 395316
rect 41321 392594 41387 392597
rect 82997 392594 83063 392597
rect 41321 392592 84210 392594
rect 41321 392536 41326 392592
rect 41382 392536 83002 392592
rect 83058 392536 84210 392592
rect 41321 392534 84210 392536
rect 41321 392531 41387 392534
rect 82997 392531 83063 392534
rect 84150 392050 84210 392534
rect 132493 392050 132559 392053
rect 84150 392048 132559 392050
rect 84150 391992 132498 392048
rect 132554 391992 132559 392048
rect 84150 391990 132559 391992
rect 132493 391987 132559 391990
rect 583520 391628 584960 391868
rect 103329 391234 103395 391237
rect 115422 391234 115428 391236
rect 103329 391232 115428 391234
rect 103329 391176 103334 391232
rect 103390 391176 115428 391232
rect 103329 391174 115428 391176
rect 103329 391171 103395 391174
rect 115422 391172 115428 391174
rect 115492 391172 115498 391236
rect 103421 390010 103487 390013
rect 116158 390010 116164 390012
rect 103421 390008 116164 390010
rect 103421 389952 103426 390008
rect 103482 389952 116164 390008
rect 103421 389950 116164 389952
rect 103421 389947 103487 389950
rect 116158 389948 116164 389950
rect 116228 389948 116234 390012
rect 96153 389874 96219 389877
rect 118918 389874 118924 389876
rect 96153 389872 118924 389874
rect 96153 389816 96158 389872
rect 96214 389816 118924 389872
rect 96153 389814 118924 389816
rect 96153 389811 96219 389814
rect 118918 389812 118924 389814
rect 118988 389874 118994 389876
rect 124254 389874 124260 389876
rect 118988 389814 124260 389874
rect 118988 389812 118994 389814
rect 124254 389812 124260 389814
rect 124324 389812 124330 389876
rect 114277 389332 114343 389333
rect 114277 389330 114324 389332
rect 114232 389328 114324 389330
rect 114232 389272 114282 389328
rect 114232 389270 114324 389272
rect 114277 389268 114324 389270
rect 114388 389268 114394 389332
rect 114277 389267 114343 389268
rect 100702 388860 100708 388924
rect 100772 388922 100778 388924
rect 101397 388922 101463 388925
rect 100772 388920 101463 388922
rect 100772 388864 101402 388920
rect 101458 388864 101463 388920
rect 100772 388862 101463 388864
rect 100772 388860 100778 388862
rect 101397 388859 101463 388862
rect 106181 388514 106247 388517
rect 119286 388514 119292 388516
rect 106181 388512 119292 388514
rect 106181 388456 106186 388512
rect 106242 388456 119292 388512
rect 106181 388454 119292 388456
rect 106181 388451 106247 388454
rect 119286 388452 119292 388454
rect 119356 388452 119362 388516
rect 58525 388380 58591 388381
rect 53598 388316 53604 388380
rect 53668 388378 53674 388380
rect 58525 388378 58572 388380
rect 53668 388376 58572 388378
rect 58636 388378 58642 388380
rect 108757 388378 108823 388381
rect 121545 388378 121611 388381
rect 53668 388320 58530 388376
rect 53668 388318 58572 388320
rect 53668 388316 53674 388318
rect 58525 388316 58572 388318
rect 58636 388318 58718 388378
rect 108757 388376 121611 388378
rect 108757 388320 108762 388376
rect 108818 388320 121550 388376
rect 121606 388320 121611 388376
rect 108757 388318 121611 388320
rect 58636 388316 58642 388318
rect 58525 388315 58591 388316
rect 108757 388315 108823 388318
rect 121545 388315 121611 388318
rect 136541 388378 136607 388381
rect 305494 388378 305500 388380
rect 136541 388376 305500 388378
rect 136541 388320 136546 388376
rect 136602 388320 305500 388376
rect 136541 388318 305500 388320
rect 136541 388315 136607 388318
rect 305494 388316 305500 388318
rect 305564 388316 305570 388380
rect 70894 387908 70900 387972
rect 70964 387970 70970 387972
rect 74625 387970 74691 387973
rect 70964 387968 74691 387970
rect 70964 387912 74630 387968
rect 74686 387912 74691 387968
rect 70964 387910 74691 387912
rect 70964 387908 70970 387910
rect 74625 387907 74691 387910
rect 112805 387970 112871 387973
rect 137134 387970 137140 387972
rect 112805 387968 137140 387970
rect 112805 387912 112810 387968
rect 112866 387912 137140 387968
rect 112805 387910 137140 387912
rect 112805 387907 112871 387910
rect 137134 387908 137140 387910
rect 137204 387970 137210 387972
rect 141141 387970 141207 387973
rect 137204 387968 141207 387970
rect 137204 387912 141146 387968
rect 141202 387912 141207 387968
rect 137204 387910 141207 387912
rect 137204 387908 137210 387910
rect 141141 387907 141207 387910
rect 55070 387772 55076 387836
rect 55140 387834 55146 387836
rect 56593 387834 56659 387837
rect 78029 387834 78095 387837
rect 55140 387832 78095 387834
rect 55140 387776 56598 387832
rect 56654 387776 78034 387832
rect 78090 387776 78095 387832
rect 55140 387774 78095 387776
rect 55140 387772 55146 387774
rect 56593 387771 56659 387774
rect 78029 387771 78095 387774
rect 117313 387700 117379 387701
rect 117262 387698 117268 387700
rect 117222 387638 117268 387698
rect 117332 387696 117379 387700
rect 117374 387640 117379 387696
rect 117262 387636 117268 387638
rect 117332 387636 117379 387640
rect 117313 387635 117379 387636
rect 50838 387092 50844 387156
rect 50908 387154 50914 387156
rect 51901 387154 51967 387157
rect 52361 387154 52427 387157
rect 50908 387152 52427 387154
rect 50908 387096 51906 387152
rect 51962 387096 52366 387152
rect 52422 387096 52427 387152
rect 50908 387094 52427 387096
rect 50908 387092 50914 387094
rect 51901 387091 51967 387094
rect 52361 387091 52427 387094
rect 127525 387018 127591 387021
rect 295374 387018 295380 387020
rect 127525 387016 295380 387018
rect 127525 386960 127530 387016
rect 127586 386960 295380 387016
rect 127525 386958 295380 386960
rect 127525 386955 127591 386958
rect 295374 386956 295380 386958
rect 295444 386956 295450 387020
rect 54937 386612 55003 386613
rect 54886 386548 54892 386612
rect 54956 386610 55003 386612
rect 54956 386608 55048 386610
rect 54998 386552 55048 386608
rect 54956 386550 55048 386552
rect 54956 386548 55003 386550
rect 54937 386547 55003 386548
rect 86217 386474 86283 386477
rect 306414 386474 306420 386476
rect 86217 386472 306420 386474
rect 86217 386416 86222 386472
rect 86278 386416 306420 386472
rect 86217 386414 306420 386416
rect 86217 386411 86283 386414
rect 306414 386412 306420 386414
rect 306484 386412 306490 386476
rect 68737 386202 68803 386205
rect 68737 386200 70226 386202
rect 68737 386144 68742 386200
rect 68798 386144 70226 386200
rect 68737 386142 70226 386144
rect 68737 386139 68803 386142
rect 70166 385250 70226 386142
rect 115289 385930 115355 385933
rect 115606 385930 115612 385932
rect 115289 385928 115612 385930
rect 115289 385872 115294 385928
rect 115350 385872 115612 385928
rect 115289 385870 115612 385872
rect 115289 385867 115355 385870
rect 115606 385868 115612 385870
rect 115676 385868 115682 385932
rect 74809 385386 74875 385389
rect 268326 385386 268332 385388
rect 74809 385384 268332 385386
rect 74809 385328 74814 385384
rect 74870 385328 268332 385384
rect 74809 385326 268332 385328
rect 74809 385323 74875 385326
rect 268326 385324 268332 385326
rect 268396 385324 268402 385388
rect 123518 385250 123524 385252
rect 70166 385190 123524 385250
rect 123518 385188 123524 385190
rect 123588 385188 123594 385252
rect 117681 384978 117747 384981
rect 118601 384978 118667 384981
rect 115828 384976 118667 384978
rect 68829 384842 68895 384845
rect 70166 384842 70226 384948
rect 115828 384920 117686 384976
rect 117742 384920 118606 384976
rect 118662 384920 118667 384976
rect 115828 384918 118667 384920
rect 117681 384915 117747 384918
rect 118601 384915 118667 384918
rect 68829 384840 70226 384842
rect 68829 384784 68834 384840
rect 68890 384784 70226 384840
rect 68829 384782 70226 384784
rect 68829 384779 68895 384782
rect -960 384284 480 384524
rect 57830 384236 57836 384300
rect 57900 384298 57906 384300
rect 69238 384298 69244 384300
rect 57900 384238 69244 384298
rect 57900 384236 57906 384238
rect 69238 384236 69244 384238
rect 69308 384236 69314 384300
rect 115798 384026 115858 384268
rect 116025 384026 116091 384029
rect 115798 384024 116091 384026
rect 115798 383968 116030 384024
rect 116086 383968 116091 384024
rect 115798 383966 116091 383968
rect 116025 383963 116091 383966
rect 116209 383618 116275 383621
rect 115828 383616 116275 383618
rect 68737 383482 68803 383485
rect 70166 383482 70226 383588
rect 115828 383560 116214 383616
rect 116270 383560 116275 383616
rect 115828 383558 116275 383560
rect 116209 383555 116275 383558
rect 68737 383480 70226 383482
rect 68737 383424 68742 383480
rect 68798 383424 70226 383480
rect 68737 383422 70226 383424
rect 68737 383419 68803 383422
rect 43897 383210 43963 383213
rect 69974 383210 69980 383212
rect 43897 383208 69980 383210
rect 43897 383152 43902 383208
rect 43958 383152 69980 383208
rect 43897 383150 69980 383152
rect 43897 383147 43963 383150
rect 69974 383148 69980 383150
rect 70044 383148 70050 383212
rect 67633 382530 67699 382533
rect 70166 382530 70226 382908
rect 67633 382528 70226 382530
rect 67633 382472 67638 382528
rect 67694 382472 70226 382528
rect 67633 382470 70226 382472
rect 67633 382467 67699 382470
rect 64638 382196 64644 382260
rect 64708 382258 64714 382260
rect 118601 382258 118667 382261
rect 64708 382198 64890 382258
rect 115828 382256 118667 382258
rect 64708 382196 64714 382198
rect 64830 382122 64890 382198
rect 66897 382122 66963 382125
rect 70166 382122 70226 382228
rect 115828 382200 118606 382256
rect 118662 382200 118667 382256
rect 115828 382198 118667 382200
rect 118601 382195 118667 382198
rect 64830 382120 70226 382122
rect 64830 382064 66902 382120
rect 66958 382064 70226 382120
rect 64830 382062 70226 382064
rect 66897 382059 66963 382062
rect 115606 381788 115612 381852
rect 115676 381850 115682 381852
rect 349797 381850 349863 381853
rect 115676 381848 349863 381850
rect 115676 381792 349802 381848
rect 349858 381792 349863 381848
rect 115676 381790 349863 381792
rect 115676 381788 115682 381790
rect 349797 381787 349863 381790
rect 118601 381578 118667 381581
rect 115828 381576 118667 381578
rect 115828 381520 118606 381576
rect 118662 381520 118667 381576
rect 115828 381518 118667 381520
rect 118601 381515 118667 381518
rect 118601 380898 118667 380901
rect 115828 380896 118667 380898
rect 67633 380762 67699 380765
rect 70166 380762 70226 380868
rect 115828 380840 118606 380896
rect 118662 380840 118667 380896
rect 115828 380838 118667 380840
rect 118601 380835 118667 380838
rect 67633 380760 70226 380762
rect 67633 380704 67638 380760
rect 67694 380704 70226 380760
rect 67633 380702 70226 380704
rect 67633 380699 67699 380702
rect 67633 379810 67699 379813
rect 70166 379810 70226 380188
rect 67633 379808 70226 379810
rect 67633 379752 67638 379808
rect 67694 379752 70226 379808
rect 67633 379750 70226 379752
rect 67633 379747 67699 379750
rect 68001 379674 68067 379677
rect 124489 379676 124555 379677
rect 68870 379674 68876 379676
rect 68001 379672 68876 379674
rect 68001 379616 68006 379672
rect 68062 379616 68876 379672
rect 68001 379614 68876 379616
rect 68001 379611 68067 379614
rect 68870 379612 68876 379614
rect 68940 379674 68946 379676
rect 124438 379674 124444 379676
rect 68940 379614 70226 379674
rect 124398 379614 124444 379674
rect 124508 379672 124555 379676
rect 124550 379616 124555 379672
rect 68940 379612 68946 379614
rect 44030 379476 44036 379540
rect 44100 379538 44106 379540
rect 64454 379538 64460 379540
rect 44100 379478 64460 379538
rect 44100 379476 44106 379478
rect 64454 379476 64460 379478
rect 64524 379538 64530 379540
rect 65149 379538 65215 379541
rect 64524 379536 65215 379538
rect 64524 379480 65154 379536
rect 65210 379480 65215 379536
rect 70166 379508 70226 379614
rect 124438 379612 124444 379614
rect 124508 379612 124555 379616
rect 124489 379611 124555 379612
rect 117998 379538 118004 379540
rect 64524 379478 65215 379480
rect 115828 379478 118004 379538
rect 64524 379476 64530 379478
rect 65149 379475 65215 379478
rect 117998 379476 118004 379478
rect 118068 379538 118074 379540
rect 118509 379538 118575 379541
rect 118068 379536 118575 379538
rect 118068 379480 118514 379536
rect 118570 379480 118575 379536
rect 118068 379478 118575 379480
rect 118068 379476 118074 379478
rect 118509 379475 118575 379478
rect 123109 378994 123175 378997
rect 123334 378994 123340 378996
rect 123109 378992 123340 378994
rect 123109 378936 123114 378992
rect 123170 378936 123340 378992
rect 123109 378934 123340 378936
rect 123109 378931 123175 378934
rect 123334 378932 123340 378934
rect 123404 378932 123410 378996
rect 118601 378858 118667 378861
rect 115828 378856 118667 378858
rect 115828 378800 118606 378856
rect 118662 378800 118667 378856
rect 115828 378798 118667 378800
rect 118601 378795 118667 378798
rect 67633 378722 67699 378725
rect 67633 378720 70226 378722
rect 67633 378664 67638 378720
rect 67694 378664 70226 378720
rect 67633 378662 70226 378664
rect 67633 378659 67699 378662
rect 70166 378148 70226 378662
rect 115381 378586 115447 378589
rect 115381 378584 115858 378586
rect 115381 378528 115386 378584
rect 115442 378528 115858 378584
rect 115381 378526 115858 378528
rect 115381 378523 115447 378526
rect 115798 378178 115858 378526
rect 580257 378450 580323 378453
rect 583520 378450 584960 378540
rect 580257 378448 584960 378450
rect 580257 378392 580262 378448
rect 580318 378392 584960 378448
rect 580257 378390 584960 378392
rect 580257 378387 580323 378390
rect 583520 378300 584960 378390
rect 117865 378178 117931 378181
rect 115798 378176 117931 378178
rect 115798 378148 117870 378176
rect 115828 378120 117870 378148
rect 117926 378120 117931 378176
rect 115828 378118 117931 378120
rect 117865 378115 117931 378118
rect 60590 377980 60596 378044
rect 60660 378042 60666 378044
rect 61878 378042 61884 378044
rect 60660 377982 61884 378042
rect 60660 377980 60666 377982
rect 61878 377980 61884 377982
rect 61948 377980 61954 378044
rect 115289 377906 115355 377909
rect 115422 377906 115428 377908
rect 115289 377904 115428 377906
rect 115289 377848 115294 377904
rect 115350 377848 115428 377904
rect 115289 377846 115428 377848
rect 115289 377843 115355 377846
rect 115422 377844 115428 377846
rect 115492 377844 115498 377908
rect 67633 377090 67699 377093
rect 70166 377090 70226 377468
rect 67633 377088 70226 377090
rect 67633 377032 67638 377088
rect 67694 377032 70226 377088
rect 67633 377030 70226 377032
rect 67633 377027 67699 377030
rect 61878 376892 61884 376956
rect 61948 376954 61954 376956
rect 61948 376894 70226 376954
rect 61948 376892 61954 376894
rect 70166 376788 70226 376894
rect 118601 376818 118667 376821
rect 115828 376816 118667 376818
rect 115828 376760 118606 376816
rect 118662 376760 118667 376816
rect 115828 376758 118667 376760
rect 118601 376755 118667 376758
rect 117313 376138 117379 376141
rect 115828 376136 117379 376138
rect 115828 376080 117318 376136
rect 117374 376080 117379 376136
rect 115828 376078 117379 376080
rect 117313 376075 117379 376078
rect 67633 376002 67699 376005
rect 119429 376002 119495 376005
rect 252870 376002 252876 376004
rect 67633 376000 70226 376002
rect 67633 375944 67638 376000
rect 67694 375944 70226 376000
rect 67633 375942 70226 375944
rect 67633 375939 67699 375942
rect 70166 375428 70226 375942
rect 119429 376000 252876 376002
rect 119429 375944 119434 376000
rect 119490 375944 252876 376000
rect 119429 375942 252876 375944
rect 119429 375939 119495 375942
rect 252870 375940 252876 375942
rect 252940 375940 252946 376004
rect 118601 375458 118667 375461
rect 115828 375456 118667 375458
rect 115828 375400 118606 375456
rect 118662 375400 118667 375456
rect 115828 375398 118667 375400
rect 118601 375395 118667 375398
rect 67633 374642 67699 374645
rect 70166 374642 70226 374748
rect 67633 374640 70226 374642
rect 67633 374584 67638 374640
rect 67694 374584 70226 374640
rect 67633 374582 70226 374584
rect 67633 374579 67699 374582
rect 69105 374234 69171 374237
rect 69105 374232 70226 374234
rect 69105 374176 69110 374232
rect 69166 374176 70226 374232
rect 69105 374174 70226 374176
rect 69105 374171 69171 374174
rect 70166 374068 70226 374174
rect 118141 374098 118207 374101
rect 115828 374096 118207 374098
rect 115828 374040 118146 374096
rect 118202 374040 118207 374096
rect 115828 374038 118207 374040
rect 118141 374035 118207 374038
rect 118325 373418 118391 373421
rect 115828 373416 118391 373418
rect 115828 373360 118330 373416
rect 118386 373360 118391 373416
rect 115828 373358 118391 373360
rect 118325 373355 118391 373358
rect 67633 373282 67699 373285
rect 67633 373280 70226 373282
rect 67633 373224 67638 373280
rect 67694 373224 70226 373280
rect 67633 373222 70226 373224
rect 67633 373219 67699 373222
rect 70166 372708 70226 373222
rect 117262 372738 117268 372740
rect 115828 372678 117268 372738
rect 117262 372676 117268 372678
rect 117332 372738 117338 372740
rect 118509 372738 118575 372741
rect 117332 372736 118575 372738
rect 117332 372680 118514 372736
rect 118570 372680 118575 372736
rect 117332 372678 118575 372680
rect 117332 372676 117338 372678
rect 118509 372675 118575 372678
rect 67633 372466 67699 372469
rect 67633 372464 70226 372466
rect 67633 372408 67638 372464
rect 67694 372408 70226 372464
rect 67633 372406 70226 372408
rect 67633 372403 67699 372406
rect 70166 372028 70226 372406
rect 67449 371786 67515 371789
rect 67449 371784 70226 371786
rect 67449 371728 67454 371784
rect 67510 371728 70226 371784
rect 67449 371726 70226 371728
rect 67449 371723 67515 371726
rect -960 371378 480 371468
rect 3233 371378 3299 371381
rect -960 371376 3299 371378
rect -960 371320 3238 371376
rect 3294 371320 3299 371376
rect 70166 371348 70226 371726
rect 116158 371378 116164 371380
rect -960 371318 3299 371320
rect 115828 371318 116164 371378
rect -960 371228 480 371318
rect 3233 371315 3299 371318
rect 116158 371316 116164 371318
rect 116228 371378 116234 371380
rect 118141 371378 118207 371381
rect 116228 371376 118207 371378
rect 116228 371320 118146 371376
rect 118202 371320 118207 371376
rect 116228 371318 118207 371320
rect 116228 371316 116234 371318
rect 118141 371315 118207 371318
rect 67725 370290 67791 370293
rect 115798 370290 115858 370668
rect 153101 370562 153167 370565
rect 299606 370562 299612 370564
rect 153101 370560 299612 370562
rect 153101 370504 153106 370560
rect 153162 370504 299612 370560
rect 153101 370502 299612 370504
rect 153101 370499 153167 370502
rect 299606 370500 299612 370502
rect 299676 370500 299682 370564
rect 115933 370290 115999 370293
rect 67725 370288 70226 370290
rect 67725 370232 67730 370288
rect 67786 370232 70226 370288
rect 67725 370230 70226 370232
rect 115798 370288 115999 370290
rect 115798 370232 115938 370288
rect 115994 370232 115999 370288
rect 115798 370230 115999 370232
rect 67725 370227 67791 370230
rect 70166 369988 70226 370230
rect 115933 370227 115999 370230
rect 116117 370018 116183 370021
rect 118141 370018 118207 370021
rect 115828 370016 118207 370018
rect 115828 369960 116122 370016
rect 116178 369960 118146 370016
rect 118202 369960 118207 370016
rect 115828 369958 118207 369960
rect 116117 369955 116183 369958
rect 118141 369955 118207 369958
rect 67633 369746 67699 369749
rect 67633 369744 70226 369746
rect 67633 369688 67638 369744
rect 67694 369688 70226 369744
rect 67633 369686 70226 369688
rect 67633 369683 67699 369686
rect 70166 369308 70226 369686
rect 67633 369066 67699 369069
rect 67633 369064 70226 369066
rect 67633 369008 67638 369064
rect 67694 369008 70226 369064
rect 67633 369006 70226 369008
rect 67633 369003 67699 369006
rect 70166 368628 70226 369006
rect 118601 368658 118667 368661
rect 115828 368656 118667 368658
rect 115828 368600 118606 368656
rect 118662 368600 118667 368656
rect 115828 368598 118667 368600
rect 118601 368595 118667 368598
rect 119521 368386 119587 368389
rect 119838 368386 119844 368388
rect 119521 368384 119844 368386
rect 119521 368328 119526 368384
rect 119582 368328 119844 368384
rect 119521 368326 119844 368328
rect 119521 368323 119587 368326
rect 119838 368324 119844 368326
rect 119908 368324 119914 368388
rect 118601 367978 118667 367981
rect 115828 367976 118667 367978
rect 115828 367920 118606 367976
rect 118662 367920 118667 367976
rect 115828 367918 118667 367920
rect 118601 367915 118667 367918
rect 119286 367644 119292 367708
rect 119356 367706 119362 367708
rect 251214 367706 251220 367708
rect 119356 367646 251220 367706
rect 119356 367644 119362 367646
rect 251214 367644 251220 367646
rect 251284 367644 251290 367708
rect 67909 367434 67975 367437
rect 68737 367434 68803 367437
rect 67909 367432 70226 367434
rect 67909 367376 67914 367432
rect 67970 367376 68742 367432
rect 68798 367376 70226 367432
rect 67909 367374 70226 367376
rect 67909 367371 67975 367374
rect 68737 367371 68803 367374
rect 70166 367268 70226 367374
rect 118601 367298 118667 367301
rect 115828 367296 118667 367298
rect 115828 367240 118606 367296
rect 118662 367240 118667 367296
rect 115828 367238 118667 367240
rect 118601 367235 118667 367238
rect 67633 366482 67699 366485
rect 70166 366482 70226 366588
rect 67633 366480 70226 366482
rect 67633 366424 67638 366480
rect 67694 366424 70226 366480
rect 67633 366422 70226 366424
rect 67633 366419 67699 366422
rect 60181 365938 60247 365941
rect 60590 365938 60596 365940
rect 60181 365936 60596 365938
rect 60181 365880 60186 365936
rect 60242 365880 60596 365936
rect 60181 365878 60596 365880
rect 60181 365875 60247 365878
rect 60590 365876 60596 365878
rect 60660 365876 60666 365940
rect 118601 365938 118667 365941
rect 115828 365936 118667 365938
rect 68461 365802 68527 365805
rect 70166 365802 70226 365908
rect 115828 365880 118606 365936
rect 118662 365880 118667 365936
rect 115828 365878 118667 365880
rect 118601 365875 118667 365878
rect 68461 365800 70226 365802
rect 68461 365744 68466 365800
rect 68522 365744 70226 365800
rect 68461 365742 70226 365744
rect 68461 365739 68527 365742
rect 118509 365258 118575 365261
rect 115828 365256 118575 365258
rect 115828 365200 118514 365256
rect 118570 365200 118575 365256
rect 115828 365198 118575 365200
rect 118509 365195 118575 365198
rect 579797 365122 579863 365125
rect 583520 365122 584960 365212
rect 579797 365120 584960 365122
rect 579797 365064 579802 365120
rect 579858 365064 584960 365120
rect 579797 365062 584960 365064
rect 579797 365059 579863 365062
rect 583520 364972 584960 365062
rect 68553 364714 68619 364717
rect 68553 364712 70226 364714
rect 68553 364656 68558 364712
rect 68614 364656 70226 364712
rect 68553 364654 70226 364656
rect 68553 364651 68619 364654
rect 70166 364548 70226 364654
rect 118601 364578 118667 364581
rect 115828 364576 118667 364578
rect 115828 364520 118606 364576
rect 118662 364520 118667 364576
rect 115828 364518 118667 364520
rect 118601 364515 118667 364518
rect 67633 363762 67699 363765
rect 70166 363762 70226 363868
rect 67633 363760 70226 363762
rect 67633 363704 67638 363760
rect 67694 363704 70226 363760
rect 67633 363702 70226 363704
rect 67633 363699 67699 363702
rect 67725 363626 67791 363629
rect 67725 363624 70226 363626
rect 67725 363568 67730 363624
rect 67786 363568 70226 363624
rect 67725 363566 70226 363568
rect 67725 363563 67791 363566
rect 70166 363188 70226 363566
rect 117405 363218 117471 363221
rect 115828 363216 117471 363218
rect 115828 363160 117410 363216
rect 117466 363160 117471 363216
rect 115828 363158 117471 363160
rect 117405 363155 117471 363158
rect 118601 362538 118667 362541
rect 115828 362536 118667 362538
rect 67633 362402 67699 362405
rect 70166 362402 70226 362508
rect 115828 362480 118606 362536
rect 118662 362480 118667 362536
rect 115828 362478 118667 362480
rect 118601 362475 118667 362478
rect 67633 362400 70226 362402
rect 67633 362344 67638 362400
rect 67694 362344 70226 362400
rect 67633 362342 70226 362344
rect 67633 362339 67699 362342
rect 118601 361858 118667 361861
rect 115828 361856 118667 361858
rect 115828 361800 118606 361856
rect 118662 361800 118667 361856
rect 115828 361798 118667 361800
rect 118601 361795 118667 361798
rect 67633 361314 67699 361317
rect 67633 361312 70226 361314
rect 67633 361256 67638 361312
rect 67694 361256 70226 361312
rect 67633 361254 70226 361256
rect 67633 361251 67699 361254
rect 70166 361148 70226 361254
rect 118049 361178 118115 361181
rect 115828 361176 118115 361178
rect 115828 361120 118054 361176
rect 118110 361120 118115 361176
rect 115828 361118 118115 361120
rect 118049 361115 118115 361118
rect 119337 360906 119403 360909
rect 255262 360906 255268 360908
rect 119337 360904 255268 360906
rect 119337 360848 119342 360904
rect 119398 360848 255268 360904
rect 119337 360846 255268 360848
rect 119337 360843 119403 360846
rect 255262 360844 255268 360846
rect 255332 360844 255338 360908
rect 67633 360634 67699 360637
rect 67633 360632 70226 360634
rect 67633 360576 67638 360632
rect 67694 360576 70226 360632
rect 67633 360574 70226 360576
rect 67633 360571 67699 360574
rect 70166 360468 70226 360574
rect 118601 359818 118667 359821
rect 115828 359816 118667 359818
rect 67633 359546 67699 359549
rect 70166 359546 70226 359788
rect 115828 359760 118606 359816
rect 118662 359760 118667 359816
rect 115828 359758 118667 359760
rect 118601 359755 118667 359758
rect 67633 359544 70226 359546
rect 67633 359488 67638 359544
rect 67694 359488 70226 359544
rect 67633 359486 70226 359488
rect 67633 359483 67699 359486
rect 117957 359138 118023 359141
rect 115828 359136 118023 359138
rect 115828 359080 117962 359136
rect 118018 359080 118023 359136
rect 115828 359078 118023 359080
rect 117957 359075 118023 359078
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect 118601 358458 118667 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect 115828 358456 118667 358458
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 67633 358186 67699 358189
rect 70166 358186 70226 358428
rect 115828 358400 118606 358456
rect 118662 358400 118667 358456
rect 115828 358398 118667 358400
rect 118601 358395 118667 358398
rect 67633 358184 70226 358186
rect 67633 358128 67638 358184
rect 67694 358128 70226 358184
rect 67633 358126 70226 358128
rect 67633 358123 67699 358126
rect 67633 357506 67699 357509
rect 70166 357506 70226 357748
rect 67633 357504 70226 357506
rect 67633 357448 67638 357504
rect 67694 357448 70226 357504
rect 67633 357446 70226 357448
rect 67633 357443 67699 357446
rect 117313 357098 117379 357101
rect 118233 357098 118299 357101
rect 115828 357096 118299 357098
rect 67633 356962 67699 356965
rect 70166 356962 70226 357068
rect 115828 357040 117318 357096
rect 117374 357040 118238 357096
rect 118294 357040 118299 357096
rect 115828 357038 118299 357040
rect 117313 357035 117379 357038
rect 118233 357035 118299 357038
rect 67633 356960 70226 356962
rect 67633 356904 67638 356960
rect 67694 356904 70226 356960
rect 67633 356902 70226 356904
rect 67633 356899 67699 356902
rect 118601 356418 118667 356421
rect 115828 356416 118667 356418
rect 115828 356360 118606 356416
rect 118662 356360 118667 356416
rect 115828 356358 118667 356360
rect 118601 356355 118667 356358
rect 67633 355874 67699 355877
rect 67633 355872 70226 355874
rect 67633 355816 67638 355872
rect 67694 355816 70226 355872
rect 67633 355814 70226 355816
rect 67633 355811 67699 355814
rect 70166 355708 70226 355814
rect 117497 355738 117563 355741
rect 118785 355738 118851 355741
rect 115828 355736 118851 355738
rect 115828 355680 117502 355736
rect 117558 355680 118790 355736
rect 118846 355680 118851 355736
rect 115828 355678 118851 355680
rect 117497 355675 117563 355678
rect 118785 355675 118851 355678
rect 67633 354786 67699 354789
rect 70166 354786 70226 355028
rect 67633 354784 70226 354786
rect 67633 354728 67638 354784
rect 67694 354728 70226 354784
rect 67633 354726 70226 354728
rect 67633 354723 67699 354726
rect 117497 354378 117563 354381
rect 115828 354376 117563 354378
rect 62614 353364 62620 353428
rect 62684 353426 62690 353428
rect 67357 353426 67423 353429
rect 70166 353426 70226 354348
rect 115828 354320 117502 354376
rect 117558 354320 117563 354376
rect 115828 354318 117563 354320
rect 117497 354315 117563 354318
rect 118601 353698 118667 353701
rect 115828 353696 118667 353698
rect 115828 353640 118606 353696
rect 118662 353640 118667 353696
rect 115828 353638 118667 353640
rect 118601 353635 118667 353638
rect 133822 353636 133828 353700
rect 133892 353698 133898 353700
rect 134057 353698 134123 353701
rect 133892 353696 134123 353698
rect 133892 353640 134062 353696
rect 134118 353640 134123 353696
rect 133892 353638 134123 353640
rect 133892 353636 133898 353638
rect 134057 353635 134123 353638
rect 62684 353424 70226 353426
rect 62684 353368 67362 353424
rect 67418 353368 70226 353424
rect 62684 353366 70226 353368
rect 62684 353364 62690 353366
rect 67357 353363 67423 353366
rect 117497 353018 117563 353021
rect 115828 353016 117563 353018
rect 68553 352746 68619 352749
rect 69197 352746 69263 352749
rect 70166 352746 70226 352988
rect 115828 352960 117502 353016
rect 117558 352960 117563 353016
rect 115828 352958 117563 352960
rect 117497 352955 117563 352958
rect 68553 352744 70226 352746
rect 68553 352688 68558 352744
rect 68614 352688 69202 352744
rect 69258 352688 70226 352744
rect 68553 352686 70226 352688
rect 68553 352683 68619 352686
rect 69197 352683 69263 352686
rect 67633 352610 67699 352613
rect 67633 352608 70226 352610
rect 67633 352552 67638 352608
rect 67694 352552 70226 352608
rect 67633 352550 70226 352552
rect 67633 352547 67699 352550
rect 70166 352308 70226 352550
rect 123518 352548 123524 352612
rect 123588 352610 123594 352612
rect 346577 352610 346643 352613
rect 123588 352608 346643 352610
rect 123588 352552 346582 352608
rect 346638 352552 346643 352608
rect 123588 352550 346643 352552
rect 123588 352548 123594 352550
rect 346577 352547 346643 352550
rect 579613 351930 579679 351933
rect 583520 351930 584960 352020
rect 579613 351928 584960 351930
rect 579613 351872 579618 351928
rect 579674 351872 584960 351928
rect 579613 351870 584960 351872
rect 579613 351867 579679 351870
rect 583520 351780 584960 351870
rect 117681 351658 117747 351661
rect 118601 351658 118667 351661
rect 115828 351656 118667 351658
rect 68001 351250 68067 351253
rect 68921 351250 68987 351253
rect 70166 351250 70226 351628
rect 115828 351600 117686 351656
rect 117742 351600 118606 351656
rect 118662 351600 118667 351656
rect 115828 351598 118667 351600
rect 117681 351595 117747 351598
rect 118601 351595 118667 351598
rect 68001 351248 70226 351250
rect 68001 351192 68006 351248
rect 68062 351192 68926 351248
rect 68982 351192 70226 351248
rect 68001 351190 70226 351192
rect 68001 351187 68067 351190
rect 68921 351187 68987 351190
rect 118049 350978 118115 350981
rect 115828 350976 118115 350978
rect 115828 350920 118054 350976
rect 118110 350920 118115 350976
rect 115828 350918 118115 350920
rect 118049 350915 118115 350918
rect 117497 350298 117563 350301
rect 115828 350296 117563 350298
rect 67633 349890 67699 349893
rect 70166 349890 70226 350268
rect 115828 350240 117502 350296
rect 117558 350240 117563 350296
rect 115828 350238 117563 350240
rect 117497 350235 117563 350238
rect 67633 349888 70226 349890
rect 67633 349832 67638 349888
rect 67694 349832 70226 349888
rect 67633 349830 70226 349832
rect 67633 349827 67699 349830
rect 67633 349210 67699 349213
rect 70166 349210 70226 349588
rect 67633 349208 70226 349210
rect 67633 349152 67638 349208
rect 67694 349152 70226 349208
rect 67633 349150 70226 349152
rect 67633 349147 67699 349150
rect 117405 348938 117471 348941
rect 118509 348938 118575 348941
rect 115828 348936 118575 348938
rect 67633 348530 67699 348533
rect 70166 348530 70226 348908
rect 115828 348880 117410 348936
rect 117466 348880 118514 348936
rect 118570 348880 118575 348936
rect 115828 348878 118575 348880
rect 117405 348875 117471 348878
rect 118509 348875 118575 348878
rect 67633 348528 70226 348530
rect 67633 348472 67638 348528
rect 67694 348472 70226 348528
rect 67633 348470 70226 348472
rect 67633 348467 67699 348470
rect 117957 348258 118023 348261
rect 115828 348256 118023 348258
rect 115828 348200 117962 348256
rect 118018 348200 118023 348256
rect 115828 348198 118023 348200
rect 117957 348195 118023 348198
rect 118601 347578 118667 347581
rect 115828 347576 118667 347578
rect 68686 347380 68692 347444
rect 68756 347442 68762 347444
rect 70166 347442 70226 347548
rect 115828 347520 118606 347576
rect 118662 347520 118667 347576
rect 115828 347518 118667 347520
rect 118601 347515 118667 347518
rect 68756 347382 70226 347442
rect 68756 347380 68762 347382
rect 67633 347306 67699 347309
rect 67633 347304 70226 347306
rect 67633 347248 67638 347304
rect 67694 347248 70226 347304
rect 67633 347246 70226 347248
rect 67633 347243 67699 347246
rect 61694 346972 61700 347036
rect 61764 347034 61770 347036
rect 68686 347034 68692 347036
rect 61764 346974 68692 347034
rect 61764 346972 61770 346974
rect 68686 346972 68692 346974
rect 68756 346972 68762 347036
rect 70166 346868 70226 347246
rect 118509 346218 118575 346221
rect 115828 346216 118575 346218
rect 66662 345884 66668 345948
rect 66732 345946 66738 345948
rect 67081 345946 67147 345949
rect 66732 345944 67147 345946
rect 66732 345888 67086 345944
rect 67142 345888 67147 345944
rect 66732 345886 67147 345888
rect 66732 345884 66738 345886
rect 67081 345883 67147 345886
rect 67633 345674 67699 345677
rect 70166 345674 70226 346188
rect 115828 346160 118514 346216
rect 118570 346160 118575 346216
rect 115828 346158 118575 346160
rect 118509 346155 118575 346158
rect 67633 345672 70226 345674
rect 67633 345616 67638 345672
rect 67694 345616 70226 345672
rect 67633 345614 70226 345616
rect 67633 345611 67699 345614
rect 118601 345538 118667 345541
rect 115828 345536 118667 345538
rect -960 345402 480 345492
rect 115828 345480 118606 345536
rect 118662 345480 118667 345536
rect 115828 345478 118667 345480
rect 118601 345475 118667 345478
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 117865 344858 117931 344861
rect 115828 344856 117931 344858
rect 115828 344828 117870 344856
rect 67633 344450 67699 344453
rect 70166 344450 70226 344828
rect 115798 344800 117870 344828
rect 117926 344800 117931 344856
rect 115798 344798 117931 344800
rect 115289 344586 115355 344589
rect 115798 344586 115858 344798
rect 117865 344795 117931 344798
rect 115289 344584 115858 344586
rect 115289 344528 115294 344584
rect 115350 344528 115858 344584
rect 115289 344526 115858 344528
rect 115289 344523 115355 344526
rect 67633 344448 70226 344450
rect 67633 344392 67638 344448
rect 67694 344392 70226 344448
rect 67633 344390 70226 344392
rect 67633 344387 67699 344390
rect 68001 344314 68067 344317
rect 68001 344312 70226 344314
rect 68001 344256 68006 344312
rect 68062 344256 70226 344312
rect 68001 344254 70226 344256
rect 68001 344251 68067 344254
rect 70166 344148 70226 344254
rect 118601 343498 118667 343501
rect 115828 343496 118667 343498
rect 67633 342954 67699 342957
rect 70166 342954 70226 343468
rect 115828 343440 118606 343496
rect 118662 343440 118667 343496
rect 115828 343438 118667 343440
rect 118601 343435 118667 343438
rect 67633 342952 70226 342954
rect 67633 342896 67638 342952
rect 67694 342896 70226 342952
rect 67633 342894 70226 342896
rect 67633 342891 67699 342894
rect 129774 342892 129780 342956
rect 129844 342954 129850 342956
rect 130101 342954 130167 342957
rect 129844 342952 130167 342954
rect 129844 342896 130106 342952
rect 130162 342896 130167 342952
rect 129844 342894 130167 342896
rect 129844 342892 129850 342894
rect 130101 342891 130167 342894
rect 118601 342818 118667 342821
rect 115828 342816 118667 342818
rect 115828 342760 118606 342816
rect 118662 342760 118667 342816
rect 115828 342758 118667 342760
rect 118601 342755 118667 342758
rect 115974 342410 115980 342412
rect 115798 342350 115980 342410
rect 115798 342138 115858 342350
rect 115974 342348 115980 342350
rect 116044 342348 116050 342412
rect 118049 342138 118115 342141
rect 115798 342136 118115 342138
rect 115798 342108 118054 342136
rect 67633 341730 67699 341733
rect 70166 341730 70226 342108
rect 115828 342080 118054 342108
rect 118110 342080 118115 342136
rect 115828 342078 118115 342080
rect 118049 342075 118115 342078
rect 67633 341728 70226 341730
rect 67633 341672 67638 341728
rect 67694 341672 70226 341728
rect 67633 341670 70226 341672
rect 67633 341667 67699 341670
rect 68645 341594 68711 341597
rect 68645 341592 70226 341594
rect 68645 341536 68650 341592
rect 68706 341536 70226 341592
rect 68645 341534 70226 341536
rect 68645 341531 68711 341534
rect 70166 341050 70226 341534
rect 70526 341050 70532 341052
rect 70166 340990 70532 341050
rect 70526 340988 70532 340990
rect 70596 340988 70602 341052
rect 118601 340778 118667 340781
rect 115828 340776 118667 340778
rect 68645 340642 68711 340645
rect 70534 340642 70594 340748
rect 115828 340720 118606 340776
rect 118662 340720 118667 340776
rect 115828 340718 118667 340720
rect 118601 340715 118667 340718
rect 68645 340640 70594 340642
rect 68645 340584 68650 340640
rect 68706 340584 70594 340640
rect 68645 340582 70594 340584
rect 68645 340579 68711 340582
rect 70534 339962 70594 340582
rect 116117 340098 116183 340101
rect 117957 340098 118023 340101
rect 115828 340096 118023 340098
rect 115828 340040 116122 340096
rect 116178 340040 117962 340096
rect 118018 340040 118023 340096
rect 115828 340038 118023 340040
rect 116117 340035 116183 340038
rect 117957 340035 118023 340038
rect 71681 339962 71747 339965
rect 70534 339960 71747 339962
rect 70534 339904 71686 339960
rect 71742 339904 71747 339960
rect 70534 339902 71747 339904
rect 71681 339899 71747 339902
rect 113189 339826 113255 339829
rect 118734 339826 118740 339828
rect 113189 339824 118740 339826
rect 113189 339768 113194 339824
rect 113250 339768 118740 339824
rect 113189 339766 118740 339768
rect 113189 339763 113255 339766
rect 118734 339764 118740 339766
rect 118804 339764 118810 339828
rect 45277 339690 45343 339693
rect 75913 339690 75979 339693
rect 77109 339690 77175 339693
rect 45277 339688 77175 339690
rect 45277 339632 45282 339688
rect 45338 339632 75918 339688
rect 75974 339632 77114 339688
rect 77170 339632 77175 339688
rect 45277 339630 77175 339632
rect 45277 339627 45343 339630
rect 75913 339627 75979 339630
rect 77109 339627 77175 339630
rect 57830 339356 57836 339420
rect 57900 339418 57906 339420
rect 73889 339418 73955 339421
rect 57900 339416 73955 339418
rect 57900 339360 73894 339416
rect 73950 339360 73955 339416
rect 57900 339358 73955 339360
rect 57900 339356 57906 339358
rect 73889 339355 73955 339358
rect 104801 339418 104867 339421
rect 121678 339418 121684 339420
rect 104801 339416 121684 339418
rect 104801 339360 104806 339416
rect 104862 339360 121684 339416
rect 104801 339358 121684 339360
rect 104801 339355 104867 339358
rect 121678 339356 121684 339358
rect 121748 339356 121754 339420
rect 107377 339282 107443 339285
rect 107561 339282 107627 339285
rect 120022 339282 120028 339284
rect 107377 339280 120028 339282
rect 107377 339224 107382 339280
rect 107438 339224 107566 339280
rect 107622 339224 120028 339280
rect 107377 339222 120028 339224
rect 107377 339219 107443 339222
rect 107561 339219 107627 339222
rect 120022 339220 120028 339222
rect 120092 339220 120098 339284
rect 61694 338812 61700 338876
rect 61764 338874 61770 338876
rect 104801 338874 104867 338877
rect 61764 338872 104867 338874
rect 61764 338816 104806 338872
rect 104862 338816 104867 338872
rect 61764 338814 104867 338816
rect 61764 338812 61770 338814
rect 104801 338811 104867 338814
rect 68870 338676 68876 338740
rect 68940 338738 68946 338740
rect 316769 338738 316835 338741
rect 68940 338736 316835 338738
rect 68940 338680 316774 338736
rect 316830 338680 316835 338736
rect 68940 338678 316835 338680
rect 68940 338676 68946 338678
rect 316769 338675 316835 338678
rect 583520 338452 584960 338692
rect 53097 338058 53163 338061
rect 71313 338058 71379 338061
rect 53097 338056 71379 338058
rect 53097 338000 53102 338056
rect 53158 338000 71318 338056
rect 71374 338000 71379 338056
rect 53097 337998 71379 338000
rect 53097 337995 53163 337998
rect 71313 337995 71379 337998
rect 73889 338058 73955 338061
rect 74441 338058 74507 338061
rect 119337 338058 119403 338061
rect 73889 338056 119403 338058
rect 73889 338000 73894 338056
rect 73950 338000 74446 338056
rect 74502 338000 119342 338056
rect 119398 338000 119403 338056
rect 73889 337998 119403 338000
rect 73889 337995 73955 337998
rect 74441 337995 74507 337998
rect 119337 337995 119403 337998
rect 71313 337378 71379 337381
rect 78029 337378 78095 337381
rect 71313 337376 78095 337378
rect 71313 337320 71318 337376
rect 71374 337320 78034 337376
rect 78090 337320 78095 337376
rect 71313 337318 78095 337320
rect 71313 337315 71379 337318
rect 78029 337315 78095 337318
rect 60590 336092 60596 336156
rect 60660 336154 60666 336156
rect 137277 336154 137343 336157
rect 60660 336152 137343 336154
rect 60660 336096 137282 336152
rect 137338 336096 137343 336152
rect 60660 336094 137343 336096
rect 60660 336092 60666 336094
rect 137277 336091 137343 336094
rect 73337 336018 73403 336021
rect 258390 336018 258396 336020
rect 73337 336016 258396 336018
rect 73337 335960 73342 336016
rect 73398 335960 258396 336016
rect 73337 335958 258396 335960
rect 73337 335955 73403 335958
rect 258390 335956 258396 335958
rect 258460 335956 258466 336020
rect 128813 335340 128879 335341
rect 128813 335336 128860 335340
rect 128924 335338 128930 335340
rect 128813 335280 128818 335336
rect 128813 335276 128860 335280
rect 128924 335278 128970 335338
rect 128924 335276 128930 335278
rect 128813 335275 128879 335276
rect 149145 334658 149211 334661
rect 241830 334658 241836 334660
rect 149145 334656 241836 334658
rect 149145 334600 149150 334656
rect 149206 334600 241836 334656
rect 149145 334598 241836 334600
rect 149145 334595 149211 334598
rect 241830 334596 241836 334598
rect 241900 334596 241906 334660
rect 59118 334052 59124 334116
rect 59188 334114 59194 334116
rect 60641 334114 60707 334117
rect 59188 334112 60707 334114
rect 59188 334056 60646 334112
rect 60702 334056 60707 334112
rect 59188 334054 60707 334056
rect 59188 334052 59194 334054
rect 60641 334051 60707 334054
rect 41229 333978 41295 333981
rect 70393 333978 70459 333981
rect 41229 333976 70459 333978
rect 41229 333920 41234 333976
rect 41290 333920 70398 333976
rect 70454 333920 70459 333976
rect 41229 333918 70459 333920
rect 41229 333915 41295 333918
rect 70393 333915 70459 333918
rect 70393 333298 70459 333301
rect 250294 333298 250300 333300
rect 70393 333296 250300 333298
rect 70393 333240 70398 333296
rect 70454 333240 250300 333296
rect 70393 333238 250300 333240
rect 70393 333235 70459 333238
rect 250294 333236 250300 333238
rect 250364 333236 250370 333300
rect -960 332196 480 332436
rect 68686 331740 68692 331804
rect 68756 331802 68762 331804
rect 248454 331802 248460 331804
rect 68756 331742 248460 331802
rect 68756 331740 68762 331742
rect 248454 331740 248460 331742
rect 248524 331740 248530 331804
rect 80973 330442 81039 330445
rect 245694 330442 245700 330444
rect 80973 330440 245700 330442
rect 80973 330384 80978 330440
rect 81034 330384 245700 330440
rect 80973 330382 245700 330384
rect 80973 330379 81039 330382
rect 245694 330380 245700 330382
rect 245764 330380 245770 330444
rect 121862 329700 121868 329764
rect 121932 329762 121938 329764
rect 122005 329762 122071 329765
rect 121932 329760 122071 329762
rect 121932 329704 122010 329760
rect 122066 329704 122071 329760
rect 121932 329702 122071 329704
rect 121932 329700 121938 329702
rect 122005 329699 122071 329702
rect 125593 328402 125659 328405
rect 125726 328402 125732 328404
rect 125593 328400 125732 328402
rect 125593 328344 125598 328400
rect 125654 328344 125732 328400
rect 125593 328342 125732 328344
rect 125593 328339 125659 328342
rect 125726 328340 125732 328342
rect 125796 328340 125802 328404
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect 67541 323642 67607 323645
rect 121678 323642 121684 323644
rect 67541 323640 121684 323642
rect 67541 323584 67546 323640
rect 67602 323584 121684 323640
rect 67541 323582 121684 323584
rect 67541 323579 67607 323582
rect 121678 323580 121684 323582
rect 121748 323580 121754 323644
rect -960 319290 480 319380
rect 3233 319290 3299 319293
rect -960 319288 3299 319290
rect -960 319232 3238 319288
rect 3294 319232 3299 319288
rect -960 319230 3299 319232
rect -960 319140 480 319230
rect 3233 319227 3299 319230
rect 67265 312626 67331 312629
rect 121862 312626 121868 312628
rect 67265 312624 121868 312626
rect 67265 312568 67270 312624
rect 67326 312568 121868 312624
rect 67265 312566 121868 312568
rect 67265 312563 67331 312566
rect 121862 312564 121868 312566
rect 121932 312564 121938 312628
rect 75913 312490 75979 312493
rect 240358 312490 240364 312492
rect 75913 312488 240364 312490
rect 75913 312432 75918 312488
rect 75974 312432 240364 312488
rect 75913 312430 240364 312432
rect 75913 312427 75979 312430
rect 240358 312428 240364 312430
rect 240428 312428 240434 312492
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect 69105 311130 69171 311133
rect 309174 311130 309180 311132
rect 69105 311128 309180 311130
rect 69105 311072 69110 311128
rect 69166 311072 309180 311128
rect 69105 311070 309180 311072
rect 69105 311067 69171 311070
rect 309174 311068 309180 311070
rect 309244 311068 309250 311132
rect 88977 309770 89043 309773
rect 247718 309770 247724 309772
rect 88977 309768 247724 309770
rect 88977 309712 88982 309768
rect 89038 309712 247724 309768
rect 88977 309710 247724 309712
rect 88977 309707 89043 309710
rect 247718 309708 247724 309710
rect 247788 309708 247794 309772
rect 64638 308348 64644 308412
rect 64708 308410 64714 308412
rect 242934 308410 242940 308412
rect 64708 308350 242940 308410
rect 64708 308348 64714 308350
rect 242934 308348 242940 308350
rect 243004 308348 243010 308412
rect 71078 307124 71084 307188
rect 71148 307186 71154 307188
rect 94221 307186 94287 307189
rect 71148 307184 94287 307186
rect 71148 307128 94226 307184
rect 94282 307128 94287 307184
rect 71148 307126 94287 307128
rect 71148 307124 71154 307126
rect 94221 307123 94287 307126
rect 70894 306988 70900 307052
rect 70964 307050 70970 307052
rect 293217 307050 293283 307053
rect 70964 307048 293283 307050
rect 70964 306992 293222 307048
rect 293278 306992 293283 307048
rect 70964 306990 293283 306992
rect 70964 306988 70970 306990
rect 293217 306987 293283 306990
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 79225 302290 79291 302293
rect 252686 302290 252692 302292
rect 79225 302288 252692 302290
rect 79225 302232 79230 302288
rect 79286 302232 252692 302288
rect 79225 302230 252692 302232
rect 79225 302227 79291 302230
rect 252686 302228 252692 302230
rect 252756 302228 252762 302292
rect 108389 301610 108455 301613
rect 108389 301608 132510 301610
rect 108389 301552 108394 301608
rect 108450 301552 132510 301608
rect 108389 301550 132510 301552
rect 108389 301547 108455 301550
rect 61469 301474 61535 301477
rect 124305 301474 124371 301477
rect 61469 301472 124371 301474
rect 61469 301416 61474 301472
rect 61530 301416 124310 301472
rect 124366 301416 124371 301472
rect 61469 301414 124371 301416
rect 132450 301474 132510 301550
rect 137134 301474 137140 301476
rect 132450 301414 137140 301474
rect 61469 301411 61535 301414
rect 124305 301411 124371 301414
rect 137134 301412 137140 301414
rect 137204 301474 137210 301476
rect 209129 301474 209195 301477
rect 137204 301472 209195 301474
rect 137204 301416 209134 301472
rect 209190 301416 209195 301472
rect 137204 301414 209195 301416
rect 137204 301412 137210 301414
rect 209129 301411 209195 301414
rect 56317 300114 56383 300117
rect 56317 300112 64890 300114
rect 56317 300056 56322 300112
rect 56378 300056 64890 300112
rect 56317 300054 64890 300056
rect 56317 300051 56383 300054
rect 64830 299570 64890 300054
rect 77293 299570 77359 299573
rect 178677 299570 178743 299573
rect 64830 299568 178743 299570
rect 64830 299512 77298 299568
rect 77354 299512 178682 299568
rect 178738 299512 178743 299568
rect 64830 299510 178743 299512
rect 77293 299507 77359 299510
rect 178677 299507 178743 299510
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 29637 298346 29703 298349
rect 118325 298346 118391 298349
rect 147949 298346 148015 298349
rect 29637 298344 148015 298346
rect 29637 298288 29642 298344
rect 29698 298288 118330 298344
rect 118386 298288 147954 298344
rect 148010 298288 148015 298344
rect 29637 298286 148015 298288
rect 29637 298283 29703 298286
rect 118325 298283 118391 298286
rect 147949 298283 148015 298286
rect 68921 298210 68987 298213
rect 282913 298210 282979 298213
rect 68921 298208 282979 298210
rect 68921 298152 68926 298208
rect 68982 298152 282918 298208
rect 282974 298152 282979 298208
rect 68921 298150 282979 298152
rect 68921 298147 68987 298150
rect 282913 298147 282979 298150
rect 80973 296986 81039 296989
rect 236494 296986 236500 296988
rect 80973 296984 236500 296986
rect 80973 296928 80978 296984
rect 81034 296928 236500 296984
rect 80973 296926 236500 296928
rect 80973 296923 81039 296926
rect 236494 296924 236500 296926
rect 236564 296924 236570 296988
rect 69841 296850 69907 296853
rect 241646 296850 241652 296852
rect 69841 296848 241652 296850
rect 69841 296792 69846 296848
rect 69902 296792 241652 296848
rect 69841 296790 241652 296792
rect 69841 296787 69907 296790
rect 241646 296788 241652 296790
rect 241716 296788 241722 296852
rect 65977 296034 66043 296037
rect 121821 296034 121887 296037
rect 65977 296032 121887 296034
rect 65977 295976 65982 296032
rect 66038 295976 121826 296032
rect 121882 295976 121887 296032
rect 65977 295974 121887 295976
rect 65977 295971 66043 295974
rect 121821 295971 121887 295974
rect 89989 295490 90055 295493
rect 126329 295490 126395 295493
rect 89989 295488 126395 295490
rect 89989 295432 89994 295488
rect 90050 295432 126334 295488
rect 126390 295432 126395 295488
rect 89989 295430 126395 295432
rect 89989 295427 90055 295430
rect 126329 295427 126395 295430
rect 114461 295354 114527 295357
rect 188429 295354 188495 295357
rect 114461 295352 188495 295354
rect 114461 295296 114466 295352
rect 114522 295296 188434 295352
rect 188490 295296 188495 295352
rect 114461 295294 188495 295296
rect 114461 295291 114527 295294
rect 188429 295291 188495 295294
rect 75821 294402 75887 294405
rect 213177 294402 213243 294405
rect 75821 294400 213243 294402
rect 75821 294344 75826 294400
rect 75882 294344 213182 294400
rect 213238 294344 213243 294400
rect 75821 294342 213243 294344
rect 75821 294339 75887 294342
rect 213177 294339 213243 294342
rect 77937 294266 78003 294269
rect 123334 294266 123340 294268
rect 77937 294264 123340 294266
rect 77937 294208 77942 294264
rect 77998 294208 123340 294264
rect 77937 294206 123340 294208
rect 77937 294203 78003 294206
rect 123334 294204 123340 294206
rect 123404 294204 123410 294268
rect 95785 294130 95851 294133
rect 177246 294130 177252 294132
rect 95785 294128 177252 294130
rect 95785 294072 95790 294128
rect 95846 294072 177252 294128
rect 95785 294070 177252 294072
rect 95785 294067 95851 294070
rect 177246 294068 177252 294070
rect 177316 294068 177322 294132
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 79409 293178 79475 293181
rect 131113 293178 131179 293181
rect 79409 293176 131179 293178
rect 79409 293120 79414 293176
rect 79470 293120 131118 293176
rect 131174 293120 131179 293176
rect 79409 293118 131179 293120
rect 79409 293115 79475 293118
rect 131113 293115 131179 293118
rect 111885 292770 111951 292773
rect 129733 292770 129799 292773
rect 111885 292768 129799 292770
rect 111885 292712 111890 292768
rect 111946 292712 129738 292768
rect 129794 292712 129799 292768
rect 111885 292710 129799 292712
rect 111885 292707 111951 292710
rect 129733 292707 129799 292710
rect 115289 292634 115355 292637
rect 115749 292634 115815 292637
rect 162209 292634 162275 292637
rect 115289 292632 162275 292634
rect 115289 292576 115294 292632
rect 115350 292576 115754 292632
rect 115810 292576 162214 292632
rect 162270 292576 162275 292632
rect 115289 292574 162275 292576
rect 115289 292571 115355 292574
rect 115749 292571 115815 292574
rect 162209 292571 162275 292574
rect 71037 292362 71103 292365
rect 70718 292360 71103 292362
rect 70718 292304 71042 292360
rect 71098 292304 71103 292360
rect 70718 292302 71103 292304
rect 70718 291788 70778 292302
rect 71037 292299 71103 292302
rect 119061 292092 119127 292093
rect 119061 292088 119108 292092
rect 119172 292090 119178 292092
rect 119061 292032 119066 292088
rect 119061 292028 119108 292032
rect 119172 292030 119218 292090
rect 119172 292028 119178 292030
rect 119061 292027 119127 292028
rect 117957 291954 118023 291957
rect 146937 291954 147003 291957
rect 117957 291952 147003 291954
rect 117957 291896 117962 291952
rect 118018 291896 146942 291952
rect 146998 291896 147003 291952
rect 117957 291894 147003 291896
rect 117957 291891 118023 291894
rect 146937 291891 147003 291894
rect 121545 291818 121611 291821
rect 119876 291816 121611 291818
rect 119876 291760 121550 291816
rect 121606 291760 121611 291816
rect 119876 291758 121611 291760
rect 121545 291755 121611 291758
rect 69982 291214 70226 291274
rect 67449 291138 67515 291141
rect 67633 291138 67699 291141
rect 69982 291138 70042 291214
rect 67449 291136 70042 291138
rect 67449 291080 67454 291136
rect 67510 291080 67638 291136
rect 67694 291080 70042 291136
rect 70166 291108 70226 291214
rect 121637 291138 121703 291141
rect 119876 291136 121703 291138
rect 67449 291078 70042 291080
rect 119876 291080 121642 291136
rect 121698 291080 121703 291136
rect 119876 291078 121703 291080
rect 67449 291075 67515 291078
rect 67633 291075 67699 291078
rect 121637 291075 121703 291078
rect 69841 290866 69907 290869
rect 69841 290864 70226 290866
rect 69841 290808 69846 290864
rect 69902 290808 70226 290864
rect 69841 290806 70226 290808
rect 69841 290803 69907 290806
rect 70166 290428 70226 290806
rect 121545 290458 121611 290461
rect 119876 290456 121611 290458
rect 119876 290400 121550 290456
rect 121606 290400 121611 290456
rect 119876 290398 121611 290400
rect 121545 290395 121611 290398
rect 121729 289778 121795 289781
rect 119876 289776 121795 289778
rect 66897 289234 66963 289237
rect 70166 289234 70226 289748
rect 119876 289720 121734 289776
rect 121790 289720 121795 289776
rect 119876 289718 121795 289720
rect 121729 289715 121795 289718
rect 66897 289232 70226 289234
rect 66897 289176 66902 289232
rect 66958 289176 70226 289232
rect 66897 289174 70226 289176
rect 66897 289171 66963 289174
rect 121637 289098 121703 289101
rect 119876 289096 121703 289098
rect 67633 288826 67699 288829
rect 70166 288826 70226 289068
rect 119876 289040 121642 289096
rect 121698 289040 121703 289096
rect 119876 289038 121703 289040
rect 121637 289035 121703 289038
rect 67633 288824 70226 288826
rect 67633 288768 67638 288824
rect 67694 288768 70226 288824
rect 67633 288766 70226 288768
rect 67633 288763 67699 288766
rect 69982 288494 70226 288554
rect 67725 288418 67791 288421
rect 69982 288418 70042 288494
rect 67725 288416 70042 288418
rect 67725 288360 67730 288416
rect 67786 288360 70042 288416
rect 70166 288388 70226 288494
rect 122281 288418 122347 288421
rect 119876 288416 122347 288418
rect 67725 288358 70042 288360
rect 119876 288360 122286 288416
rect 122342 288360 122347 288416
rect 119876 288358 122347 288360
rect 67725 288355 67791 288358
rect 122281 288355 122347 288358
rect 68185 288146 68251 288149
rect 68185 288144 70226 288146
rect 68185 288088 68190 288144
rect 68246 288088 70226 288144
rect 68185 288086 70226 288088
rect 68185 288083 68251 288086
rect 70166 287708 70226 288086
rect 121545 287738 121611 287741
rect 119876 287736 121611 287738
rect 119876 287680 121550 287736
rect 121606 287680 121611 287736
rect 119876 287678 121611 287680
rect 121545 287675 121611 287678
rect 69105 287058 69171 287061
rect 69982 287058 70226 287070
rect 121545 287058 121611 287061
rect 69105 287056 70226 287058
rect 69105 287000 69110 287056
rect 69166 287010 70226 287056
rect 119876 287056 121611 287058
rect 69166 287000 70042 287010
rect 69105 286998 70042 287000
rect 119876 287000 121550 287056
rect 121606 287000 121611 287056
rect 119876 286998 121611 287000
rect 69105 286995 69171 286998
rect 121545 286995 121611 286998
rect 70526 286724 70532 286788
rect 70596 286724 70602 286788
rect 70534 286348 70594 286724
rect 119286 286452 119292 286516
rect 119356 286514 119362 286516
rect 285622 286514 285628 286516
rect 119356 286454 285628 286514
rect 119356 286452 119362 286454
rect 285622 286452 285628 286454
rect 285692 286452 285698 286516
rect 121637 286378 121703 286381
rect 119876 286376 121703 286378
rect 119876 286320 121642 286376
rect 121698 286320 121703 286376
rect 119876 286318 121703 286320
rect 121637 286315 121703 286318
rect 68921 286106 68987 286109
rect 68921 286104 70226 286106
rect 68921 286048 68926 286104
rect 68982 286048 70226 286104
rect 68921 286046 70226 286048
rect 68921 286043 68987 286046
rect 70166 285668 70226 286046
rect 121453 285698 121519 285701
rect 119876 285696 121519 285698
rect 119876 285640 121458 285696
rect 121514 285640 121519 285696
rect 119876 285638 121519 285640
rect 121453 285635 121519 285638
rect 67541 285426 67607 285429
rect 67541 285424 70226 285426
rect 67541 285368 67546 285424
rect 67602 285368 70226 285424
rect 67541 285366 70226 285368
rect 67541 285363 67607 285366
rect 70166 284988 70226 285366
rect 583520 285276 584960 285516
rect 121453 285018 121519 285021
rect 119876 285016 121519 285018
rect 119876 284960 121458 285016
rect 121514 284960 121519 285016
rect 119876 284958 121519 284960
rect 121453 284955 121519 284958
rect 67633 284474 67699 284477
rect 67633 284472 70226 284474
rect 67633 284416 67638 284472
rect 67694 284416 70226 284472
rect 67633 284414 70226 284416
rect 67633 284411 67699 284414
rect 70166 284308 70226 284414
rect 120901 284338 120967 284341
rect 119876 284336 120967 284338
rect 119876 284280 120906 284336
rect 120962 284280 120967 284336
rect 119876 284278 120967 284280
rect 120901 284275 120967 284278
rect 68829 283794 68895 283797
rect 68829 283792 70226 283794
rect 68829 283736 68834 283792
rect 68890 283736 70226 283792
rect 68829 283734 70226 283736
rect 68829 283731 68895 283734
rect 70166 283628 70226 283734
rect 67725 283386 67791 283389
rect 67725 283384 70226 283386
rect 67725 283328 67730 283384
rect 67786 283328 70226 283384
rect 67725 283326 70226 283328
rect 67725 283323 67791 283326
rect 70166 282948 70226 283326
rect 119846 283114 119906 283628
rect 119846 283054 122850 283114
rect 121453 282978 121519 282981
rect 119876 282976 121519 282978
rect 119876 282920 121458 282976
rect 121514 282920 121519 282976
rect 119876 282918 121519 282920
rect 121453 282915 121519 282918
rect 122790 282842 122850 283054
rect 132493 282842 132559 282845
rect 133781 282842 133847 282845
rect 122790 282840 133847 282842
rect 122790 282784 132498 282840
rect 132554 282784 133786 282840
rect 133842 282784 133847 282840
rect 122790 282782 133847 282784
rect 132493 282779 132559 282782
rect 133781 282779 133847 282782
rect 69197 282162 69263 282165
rect 69197 282160 70226 282162
rect 69197 282104 69202 282160
rect 69258 282104 70226 282160
rect 69197 282102 70226 282104
rect 69197 282099 69263 282102
rect 70166 281588 70226 282102
rect 119846 281890 119906 282268
rect 133781 282162 133847 282165
rect 304206 282162 304212 282164
rect 133781 282160 304212 282162
rect 133781 282104 133786 282160
rect 133842 282104 304212 282160
rect 133781 282102 304212 282104
rect 133781 282099 133847 282102
rect 304206 282100 304212 282102
rect 304276 282100 304282 282164
rect 227662 281890 227668 281892
rect 119846 281830 227668 281890
rect 227662 281828 227668 281830
rect 227732 281828 227738 281892
rect 121453 281618 121519 281621
rect 119876 281616 121519 281618
rect 119876 281560 121458 281616
rect 121514 281560 121519 281616
rect 119876 281558 121519 281560
rect 121453 281555 121519 281558
rect 67725 280530 67791 280533
rect 70166 280530 70226 280908
rect 67725 280528 70226 280530
rect 67725 280472 67730 280528
rect 67786 280472 70226 280528
rect 67725 280470 70226 280472
rect 119846 280530 119906 280908
rect 285806 280530 285812 280532
rect 119846 280470 285812 280530
rect 67725 280467 67791 280470
rect 285806 280468 285812 280470
rect 285876 280468 285882 280532
rect 67633 280394 67699 280397
rect 67633 280392 70226 280394
rect 67633 280336 67638 280392
rect 67694 280336 70226 280392
rect 67633 280334 70226 280336
rect 67633 280331 67699 280334
rect 70166 280228 70226 280334
rect 121453 280258 121519 280261
rect 119876 280256 121519 280258
rect -960 279972 480 280212
rect 119876 280200 121458 280256
rect 121514 280200 121519 280256
rect 119876 280198 121519 280200
rect 121453 280195 121519 280198
rect 121545 279578 121611 279581
rect 119876 279576 121611 279578
rect 67633 279170 67699 279173
rect 70166 279170 70226 279548
rect 119876 279520 121550 279576
rect 121606 279520 121611 279576
rect 119876 279518 121611 279520
rect 121545 279515 121611 279518
rect 67633 279168 70226 279170
rect 67633 279112 67638 279168
rect 67694 279112 70226 279168
rect 67633 279110 70226 279112
rect 67633 279107 67699 279110
rect 58566 278972 58572 279036
rect 58636 279034 58642 279036
rect 58636 278974 70226 279034
rect 58636 278972 58642 278974
rect 70166 278868 70226 278974
rect 121453 278898 121519 278901
rect 119876 278896 121519 278898
rect 119876 278840 121458 278896
rect 121514 278840 121519 278896
rect 119876 278838 121519 278840
rect 121453 278835 121519 278838
rect 121545 278218 121611 278221
rect 119876 278216 121611 278218
rect 67633 277810 67699 277813
rect 70166 277810 70226 278188
rect 119876 278160 121550 278216
rect 121606 278160 121611 278216
rect 119876 278158 121611 278160
rect 121545 278155 121611 278158
rect 67633 277808 70226 277810
rect 67633 277752 67638 277808
rect 67694 277752 70226 277808
rect 67633 277750 70226 277752
rect 67633 277747 67699 277750
rect 68277 277674 68343 277677
rect 68277 277672 70226 277674
rect 68277 277616 68282 277672
rect 68338 277616 70226 277672
rect 68277 277614 70226 277616
rect 68277 277611 68343 277614
rect 70166 277508 70226 277614
rect 121453 277538 121519 277541
rect 119876 277536 121519 277538
rect 119876 277480 121458 277536
rect 121514 277480 121519 277536
rect 119876 277478 121519 277480
rect 121453 277475 121519 277478
rect 121862 276858 121868 276860
rect 67725 276450 67791 276453
rect 70166 276450 70226 276828
rect 119876 276798 121868 276858
rect 121862 276796 121868 276798
rect 121932 276796 121938 276860
rect 67725 276448 70226 276450
rect 67725 276392 67730 276448
rect 67786 276392 70226 276448
rect 67725 276390 70226 276392
rect 67725 276387 67791 276390
rect 67633 276314 67699 276317
rect 67633 276312 70226 276314
rect 67633 276256 67638 276312
rect 67694 276256 70226 276312
rect 67633 276254 70226 276256
rect 67633 276251 67699 276254
rect 70166 276148 70226 276254
rect 120022 276252 120028 276316
rect 120092 276314 120098 276316
rect 121637 276314 121703 276317
rect 120092 276312 121703 276314
rect 120092 276256 121642 276312
rect 121698 276256 121703 276312
rect 120092 276254 121703 276256
rect 120092 276252 120098 276254
rect 121637 276251 121703 276254
rect 121453 276178 121519 276181
rect 119876 276176 121519 276178
rect 119876 276120 121458 276176
rect 121514 276120 121519 276176
rect 119876 276118 121519 276120
rect 121453 276115 121519 276118
rect 121913 276044 121979 276045
rect 121862 276042 121868 276044
rect 121822 275982 121868 276042
rect 121932 276040 121979 276044
rect 121974 275984 121979 276040
rect 121862 275980 121868 275982
rect 121932 275980 121979 275984
rect 121913 275979 121979 275980
rect 121545 275498 121611 275501
rect 119876 275496 121611 275498
rect 67725 275090 67791 275093
rect 70166 275090 70226 275468
rect 119876 275440 121550 275496
rect 121606 275440 121611 275496
rect 119876 275438 121611 275440
rect 121545 275435 121611 275438
rect 67725 275088 70226 275090
rect 67725 275032 67730 275088
rect 67786 275032 70226 275088
rect 67725 275030 70226 275032
rect 67725 275027 67791 275030
rect 67633 274954 67699 274957
rect 67633 274952 70226 274954
rect 67633 274896 67638 274952
rect 67694 274896 70226 274952
rect 67633 274894 70226 274896
rect 67633 274891 67699 274894
rect 70166 274788 70226 274894
rect 121453 274818 121519 274821
rect 119876 274816 121519 274818
rect 119876 274760 121458 274816
rect 121514 274760 121519 274816
rect 119876 274758 121519 274760
rect 121453 274755 121519 274758
rect 122097 274138 122163 274141
rect 119876 274136 122163 274138
rect 69054 273594 69060 273596
rect 64830 273534 69060 273594
rect 39849 273458 39915 273461
rect 64830 273458 64890 273534
rect 69054 273532 69060 273534
rect 69124 273594 69130 273596
rect 70166 273594 70226 274108
rect 119876 274080 122102 274136
rect 122158 274080 122163 274136
rect 119876 274078 122163 274080
rect 122097 274075 122163 274078
rect 69124 273534 70226 273594
rect 69124 273532 69130 273534
rect 121453 273458 121519 273461
rect 39849 273456 64890 273458
rect 39849 273400 39854 273456
rect 39910 273400 64890 273456
rect 119876 273456 121519 273458
rect 39849 273398 64890 273400
rect 39849 273395 39915 273398
rect 67633 273322 67699 273325
rect 67633 273320 69858 273322
rect 67633 273264 67638 273320
rect 67694 273264 69858 273320
rect 67633 273262 69858 273264
rect 67633 273259 67699 273262
rect 69798 273186 69858 273262
rect 70350 273186 70410 273428
rect 119876 273400 121458 273456
rect 121514 273400 121519 273456
rect 119876 273398 121519 273400
rect 121453 273395 121519 273398
rect 69798 273126 70410 273186
rect 121453 272778 121519 272781
rect 119876 272776 121519 272778
rect 67633 272370 67699 272373
rect 70166 272370 70226 272748
rect 119876 272720 121458 272776
rect 121514 272720 121519 272776
rect 119876 272718 121519 272720
rect 121453 272715 121519 272718
rect 121913 272506 121979 272509
rect 298686 272506 298692 272508
rect 121913 272504 298692 272506
rect 121913 272448 121918 272504
rect 121974 272448 298692 272504
rect 121913 272446 298692 272448
rect 121913 272443 121979 272446
rect 298686 272444 298692 272446
rect 298756 272444 298762 272508
rect 67633 272368 70226 272370
rect 67633 272312 67638 272368
rect 67694 272312 70226 272368
rect 67633 272310 70226 272312
rect 67633 272307 67699 272310
rect 68093 272234 68159 272237
rect 580257 272234 580323 272237
rect 583520 272234 584960 272324
rect 68093 272232 70226 272234
rect 68093 272176 68098 272232
rect 68154 272176 70226 272232
rect 68093 272174 70226 272176
rect 68093 272171 68159 272174
rect 70166 272068 70226 272174
rect 580257 272232 584960 272234
rect 580257 272176 580262 272232
rect 580318 272176 584960 272232
rect 580257 272174 584960 272176
rect 580257 272171 580323 272174
rect 121453 272098 121519 272101
rect 119876 272096 121519 272098
rect 119876 272040 121458 272096
rect 121514 272040 121519 272096
rect 583520 272084 584960 272174
rect 119876 272038 121519 272040
rect 121453 272035 121519 272038
rect 67725 271554 67791 271557
rect 67725 271552 70226 271554
rect 67725 271496 67730 271552
rect 67786 271496 70226 271552
rect 67725 271494 70226 271496
rect 67725 271491 67791 271494
rect 70166 271388 70226 271494
rect 121453 271418 121519 271421
rect 119876 271416 121519 271418
rect 119876 271360 121458 271416
rect 121514 271360 121519 271416
rect 119876 271358 121519 271360
rect 121453 271355 121519 271358
rect 67633 271146 67699 271149
rect 67633 271144 70226 271146
rect 67633 271088 67638 271144
rect 67694 271088 70226 271144
rect 67633 271086 70226 271088
rect 67633 271083 67699 271086
rect 70166 270708 70226 271086
rect 121453 270058 121519 270061
rect 119876 270056 121519 270058
rect 67725 269650 67791 269653
rect 70166 269650 70226 270028
rect 119876 270000 121458 270056
rect 121514 270000 121519 270056
rect 119876 269998 121519 270000
rect 121453 269995 121519 269998
rect 67725 269648 70226 269650
rect 67725 269592 67730 269648
rect 67786 269592 70226 269648
rect 67725 269590 70226 269592
rect 67725 269587 67791 269590
rect 67633 269514 67699 269517
rect 67633 269512 70226 269514
rect 67633 269456 67638 269512
rect 67694 269456 70226 269512
rect 67633 269454 70226 269456
rect 67633 269451 67699 269454
rect 70166 269348 70226 269454
rect 121545 269378 121611 269381
rect 119876 269376 121611 269378
rect 119876 269320 121550 269376
rect 121606 269320 121611 269376
rect 119876 269318 121611 269320
rect 121545 269315 121611 269318
rect 67449 268834 67515 268837
rect 67449 268832 70226 268834
rect 67449 268776 67454 268832
rect 67510 268776 70226 268832
rect 67449 268774 70226 268776
rect 67449 268771 67515 268774
rect 70166 268668 70226 268774
rect 121453 268698 121519 268701
rect 119876 268696 121519 268698
rect 119876 268640 121458 268696
rect 121514 268640 121519 268696
rect 119876 268638 121519 268640
rect 121453 268635 121519 268638
rect 67725 268426 67791 268429
rect 67725 268424 70226 268426
rect 67725 268368 67730 268424
rect 67786 268368 70226 268424
rect 67725 268366 70226 268368
rect 67725 268363 67791 268366
rect 70166 267988 70226 268366
rect 121545 268018 121611 268021
rect 119876 268016 121611 268018
rect 119876 267960 121550 268016
rect 121606 267960 121611 268016
rect 119876 267958 121611 267960
rect 121545 267955 121611 267958
rect 121637 267338 121703 267341
rect 119876 267336 121703 267338
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 67725 266930 67791 266933
rect 70166 266930 70226 267308
rect 119876 267280 121642 267336
rect 121698 267280 121703 267336
rect 119876 267278 121703 267280
rect 121637 267275 121703 267278
rect 67725 266928 70226 266930
rect 67725 266872 67730 266928
rect 67786 266872 70226 266928
rect 67725 266870 70226 266872
rect 67725 266867 67791 266870
rect 67633 266794 67699 266797
rect 67633 266792 70226 266794
rect 67633 266736 67638 266792
rect 67694 266736 70226 266792
rect 67633 266734 70226 266736
rect 67633 266731 67699 266734
rect 70166 266628 70226 266734
rect 121545 266658 121611 266661
rect 119876 266656 121611 266658
rect 119876 266600 121550 266656
rect 121606 266600 121611 266656
rect 119876 266598 121611 266600
rect 121545 266595 121611 266598
rect 121637 265978 121703 265981
rect 119876 265976 121703 265978
rect 61694 265644 61700 265708
rect 61764 265706 61770 265708
rect 62021 265706 62087 265709
rect 61764 265704 62087 265706
rect 61764 265648 62026 265704
rect 62082 265648 62087 265704
rect 61764 265646 62087 265648
rect 61764 265644 61770 265646
rect 62021 265643 62087 265646
rect 67725 265570 67791 265573
rect 70166 265570 70226 265948
rect 119876 265920 121642 265976
rect 121698 265920 121703 265976
rect 119876 265918 121703 265920
rect 121637 265915 121703 265918
rect 67725 265568 70226 265570
rect 67725 265512 67730 265568
rect 67786 265512 70226 265568
rect 67725 265510 70226 265512
rect 67725 265507 67791 265510
rect 67633 265434 67699 265437
rect 67633 265432 70226 265434
rect 67633 265376 67638 265432
rect 67694 265376 70226 265432
rect 67633 265374 70226 265376
rect 67633 265371 67699 265374
rect 70166 265268 70226 265374
rect 121545 265298 121611 265301
rect 119876 265296 121611 265298
rect 119876 265240 121550 265296
rect 121606 265240 121611 265296
rect 119876 265238 121611 265240
rect 121545 265235 121611 265238
rect 67633 264890 67699 264893
rect 67633 264888 70226 264890
rect 67633 264832 67638 264888
rect 67694 264832 70226 264888
rect 67633 264830 70226 264832
rect 67633 264827 67699 264830
rect 70166 264588 70226 264830
rect 124305 264618 124371 264621
rect 119876 264616 124371 264618
rect 119876 264560 124310 264616
rect 124366 264560 124371 264616
rect 119876 264558 124371 264560
rect 124305 264555 124371 264558
rect 121637 263938 121703 263941
rect 119876 263936 121703 263938
rect 68921 263666 68987 263669
rect 70166 263666 70226 263908
rect 119876 263880 121642 263936
rect 121698 263880 121703 263936
rect 119876 263878 121703 263880
rect 121637 263875 121703 263878
rect 68921 263664 70226 263666
rect 68921 263608 68926 263664
rect 68982 263608 70226 263664
rect 68921 263606 70226 263608
rect 68921 263603 68987 263606
rect 121545 263258 121611 263261
rect 119876 263256 121611 263258
rect 67725 262850 67791 262853
rect 70166 262850 70226 263228
rect 119876 263200 121550 263256
rect 121606 263200 121611 263256
rect 119876 263198 121611 263200
rect 121545 263195 121611 263198
rect 67725 262848 70226 262850
rect 67725 262792 67730 262848
rect 67786 262792 70226 262848
rect 67725 262790 70226 262792
rect 124305 262850 124371 262853
rect 302734 262850 302740 262852
rect 124305 262848 302740 262850
rect 124305 262792 124310 262848
rect 124366 262792 302740 262848
rect 124305 262790 302740 262792
rect 67725 262787 67791 262790
rect 124305 262787 124371 262790
rect 302734 262788 302740 262790
rect 302804 262788 302810 262852
rect 121545 262578 121611 262581
rect 119876 262576 121611 262578
rect 67633 262306 67699 262309
rect 70166 262306 70226 262548
rect 119876 262520 121550 262576
rect 121606 262520 121611 262576
rect 119876 262518 121611 262520
rect 121545 262515 121611 262518
rect 67633 262304 70226 262306
rect 67633 262248 67638 262304
rect 67694 262248 70226 262304
rect 67633 262246 70226 262248
rect 67633 262243 67699 262246
rect 121637 261898 121703 261901
rect 119876 261896 121703 261898
rect 67725 261490 67791 261493
rect 70166 261490 70226 261868
rect 119876 261840 121642 261896
rect 121698 261840 121703 261896
rect 119876 261838 121703 261840
rect 121637 261835 121703 261838
rect 67725 261488 70226 261490
rect 67725 261432 67730 261488
rect 67786 261432 70226 261488
rect 67725 261430 70226 261432
rect 67725 261427 67791 261430
rect 121545 261218 121611 261221
rect 119876 261216 121611 261218
rect 66110 260884 66116 260948
rect 66180 260946 66186 260948
rect 70166 260946 70226 261188
rect 119876 261160 121550 261216
rect 121606 261160 121611 261216
rect 119876 261158 121611 261160
rect 121545 261155 121611 261158
rect 66180 260886 70226 260946
rect 66180 260884 66186 260886
rect 67633 260810 67699 260813
rect 67633 260808 70226 260810
rect 67633 260752 67638 260808
rect 67694 260752 70226 260808
rect 67633 260750 70226 260752
rect 67633 260747 67699 260750
rect 70166 260508 70226 260750
rect 121545 260538 121611 260541
rect 119876 260536 121611 260538
rect 119876 260480 121550 260536
rect 121606 260480 121611 260536
rect 119876 260478 121611 260480
rect 121545 260475 121611 260478
rect 121545 259858 121611 259861
rect 119876 259856 121611 259858
rect 67633 259586 67699 259589
rect 70350 259586 70410 259828
rect 119876 259800 121550 259856
rect 121606 259800 121611 259856
rect 119876 259798 121611 259800
rect 121545 259795 121611 259798
rect 67633 259584 70410 259586
rect 67633 259528 67638 259584
rect 67694 259528 70410 259584
rect 67633 259526 70410 259528
rect 67633 259523 67699 259526
rect 121729 259178 121795 259181
rect 119876 259176 121795 259178
rect 67725 258634 67791 258637
rect 70166 258634 70226 259148
rect 119876 259120 121734 259176
rect 121790 259120 121795 259176
rect 119876 259118 121795 259120
rect 121729 259115 121795 259118
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 123334 258708 123340 258772
rect 123404 258770 123410 258772
rect 430614 258770 430620 258772
rect 123404 258710 430620 258770
rect 123404 258708 123410 258710
rect 430614 258708 430620 258710
rect 430684 258708 430690 258772
rect 583520 258756 584960 258846
rect 67725 258632 70226 258634
rect 67725 258576 67730 258632
rect 67786 258576 70226 258632
rect 67725 258574 70226 258576
rect 67725 258571 67791 258574
rect 121545 258498 121611 258501
rect 119876 258496 121611 258498
rect 67633 258226 67699 258229
rect 70166 258226 70226 258468
rect 119876 258440 121550 258496
rect 121606 258440 121611 258496
rect 119876 258438 121611 258440
rect 121545 258435 121611 258438
rect 67633 258224 70226 258226
rect 67633 258168 67638 258224
rect 67694 258168 70226 258224
rect 67633 258166 70226 258168
rect 67633 258163 67699 258166
rect 121453 257818 121519 257821
rect 119876 257816 121519 257818
rect 67725 257274 67791 257277
rect 70166 257274 70226 257788
rect 119876 257760 121458 257816
rect 121514 257760 121519 257816
rect 119876 257758 121519 257760
rect 121453 257755 121519 257758
rect 67725 257272 70226 257274
rect 67725 257216 67730 257272
rect 67786 257216 70226 257272
rect 67725 257214 70226 257216
rect 67725 257211 67791 257214
rect 121269 257138 121335 257141
rect 119876 257136 121335 257138
rect 67633 256866 67699 256869
rect 70166 256866 70226 257108
rect 119876 257080 121274 257136
rect 121330 257080 121335 257136
rect 119876 257078 121335 257080
rect 121269 257075 121335 257078
rect 67633 256864 70226 256866
rect 67633 256808 67638 256864
rect 67694 256808 70226 256864
rect 67633 256806 70226 256808
rect 67633 256803 67699 256806
rect 121453 256458 121519 256461
rect 119876 256456 121519 256458
rect 67633 255914 67699 255917
rect 70166 255914 70226 256428
rect 119876 256400 121458 256456
rect 121514 256400 121519 256456
rect 119876 256398 121519 256400
rect 121453 256395 121519 256398
rect 67633 255912 70226 255914
rect 67633 255856 67638 255912
rect 67694 255856 70226 255912
rect 67633 255854 70226 255856
rect 67633 255851 67699 255854
rect 122741 255778 122807 255781
rect 119876 255776 122807 255778
rect 67725 255370 67791 255373
rect 70166 255370 70226 255748
rect 119876 255720 122746 255776
rect 122802 255720 122807 255776
rect 119876 255718 122807 255720
rect 122741 255715 122807 255718
rect 67725 255368 70226 255370
rect 67725 255312 67730 255368
rect 67786 255312 70226 255368
rect 67725 255310 70226 255312
rect 67725 255307 67791 255310
rect 67633 255234 67699 255237
rect 67633 255232 70226 255234
rect 67633 255176 67638 255232
rect 67694 255176 70226 255232
rect 67633 255174 70226 255176
rect 67633 255171 67699 255174
rect 70166 255068 70226 255174
rect 121637 255098 121703 255101
rect 119876 255096 121703 255098
rect 119876 255040 121642 255096
rect 121698 255040 121703 255096
rect 119876 255038 121703 255040
rect 121637 255035 121703 255038
rect 67633 254554 67699 254557
rect 67633 254552 70226 254554
rect 67633 254496 67638 254552
rect 67694 254496 70226 254552
rect 67633 254494 70226 254496
rect 67633 254491 67699 254494
rect 70166 254388 70226 254494
rect 121453 254418 121519 254421
rect 119876 254416 121519 254418
rect 119876 254360 121458 254416
rect 121514 254360 121519 254416
rect 119876 254358 121519 254360
rect 121453 254355 121519 254358
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 121637 253738 121703 253741
rect 119876 253736 121703 253738
rect 69013 253194 69079 253197
rect 70166 253194 70226 253708
rect 119876 253680 121642 253736
rect 121698 253680 121703 253736
rect 119876 253678 121703 253680
rect 121637 253675 121703 253678
rect 69013 253192 70226 253194
rect 69013 253136 69018 253192
rect 69074 253136 70226 253192
rect 69013 253134 70226 253136
rect 69013 253131 69079 253134
rect 121453 253058 121519 253061
rect 119876 253056 121519 253058
rect 68093 252650 68159 252653
rect 70166 252650 70226 253028
rect 119876 253000 121458 253056
rect 121514 253000 121519 253056
rect 119876 252998 121519 253000
rect 121453 252995 121519 252998
rect 68093 252648 70226 252650
rect 68093 252592 68098 252648
rect 68154 252592 70226 252648
rect 68093 252590 70226 252592
rect 68093 252587 68159 252590
rect 121729 252378 121795 252381
rect 119876 252376 121795 252378
rect 67633 251834 67699 251837
rect 70166 251834 70226 252348
rect 119876 252320 121734 252376
rect 121790 252320 121795 252376
rect 119876 252318 121795 252320
rect 121729 252315 121795 252318
rect 67633 251832 70226 251834
rect 67633 251776 67638 251832
rect 67694 251776 70226 251832
rect 67633 251774 70226 251776
rect 67633 251771 67699 251774
rect 121453 251698 121519 251701
rect 119876 251696 121519 251698
rect 69105 251290 69171 251293
rect 70166 251290 70226 251668
rect 119876 251640 121458 251696
rect 121514 251640 121519 251696
rect 119876 251638 121519 251640
rect 121453 251635 121519 251638
rect 69105 251288 70226 251290
rect 69105 251232 69110 251288
rect 69166 251232 70226 251288
rect 69105 251230 70226 251232
rect 69105 251227 69171 251230
rect 120073 251018 120139 251021
rect 119876 251016 120139 251018
rect 67725 250474 67791 250477
rect 70166 250474 70226 250988
rect 119876 250960 120078 251016
rect 120134 250960 120139 251016
rect 119876 250958 120139 250960
rect 120073 250955 120139 250958
rect 67725 250472 70226 250474
rect 67725 250416 67730 250472
rect 67786 250416 70226 250472
rect 67725 250414 70226 250416
rect 67725 250411 67791 250414
rect 121453 250338 121519 250341
rect 119876 250336 121519 250338
rect 67633 249930 67699 249933
rect 70166 249930 70226 250308
rect 119876 250280 121458 250336
rect 121514 250280 121519 250336
rect 119876 250278 121519 250280
rect 121453 250275 121519 250278
rect 67633 249928 70226 249930
rect 67633 249872 67638 249928
rect 67694 249872 70226 249928
rect 67633 249870 70226 249872
rect 67633 249867 67699 249870
rect 121637 249658 121703 249661
rect 119876 249656 121703 249658
rect 67725 249114 67791 249117
rect 70166 249114 70226 249628
rect 119876 249600 121642 249656
rect 121698 249600 121703 249656
rect 119876 249598 121703 249600
rect 121637 249595 121703 249598
rect 67725 249112 70226 249114
rect 67725 249056 67730 249112
rect 67786 249056 70226 249112
rect 67725 249054 70226 249056
rect 67725 249051 67791 249054
rect 121453 248978 121519 248981
rect 119876 248976 121519 248978
rect 67633 248570 67699 248573
rect 70166 248570 70226 248948
rect 119876 248920 121458 248976
rect 121514 248920 121519 248976
rect 119876 248918 121519 248920
rect 121453 248915 121519 248918
rect 67633 248568 70226 248570
rect 67633 248512 67638 248568
rect 67694 248512 70226 248568
rect 67633 248510 70226 248512
rect 67633 248507 67699 248510
rect 121453 248298 121519 248301
rect 119876 248296 121519 248298
rect 67725 247754 67791 247757
rect 70166 247754 70226 248268
rect 119876 248240 121458 248296
rect 121514 248240 121519 248296
rect 119876 248238 121519 248240
rect 121453 248235 121519 248238
rect 67725 247752 70226 247754
rect 67725 247696 67730 247752
rect 67786 247696 70226 247752
rect 67725 247694 70226 247696
rect 67725 247691 67791 247694
rect 121361 247618 121427 247621
rect 119876 247616 121427 247618
rect 67633 247210 67699 247213
rect 70166 247210 70226 247588
rect 119876 247560 121366 247616
rect 121422 247560 121427 247616
rect 119876 247558 121427 247560
rect 121361 247555 121427 247558
rect 67633 247208 70226 247210
rect 67633 247152 67638 247208
rect 67694 247152 70226 247208
rect 67633 247150 70226 247152
rect 67633 247147 67699 247150
rect 57838 247014 67650 247074
rect 50705 246938 50771 246941
rect 57094 246938 57100 246940
rect 50705 246936 57100 246938
rect 50705 246880 50710 246936
rect 50766 246880 57100 246936
rect 50705 246878 57100 246880
rect 50705 246875 50771 246878
rect 57094 246876 57100 246878
rect 57164 246938 57170 246940
rect 57838 246938 57898 247014
rect 57164 246878 57898 246938
rect 67590 246938 67650 247014
rect 69982 247014 70226 247074
rect 69982 246938 70042 247014
rect 67590 246878 70042 246938
rect 70166 246908 70226 247014
rect 121545 246938 121611 246941
rect 119876 246936 121611 246938
rect 119876 246880 121550 246936
rect 121606 246880 121611 246936
rect 119876 246878 121611 246880
rect 57164 246876 57170 246878
rect 121545 246875 121611 246878
rect 121453 246258 121519 246261
rect 119876 246256 121519 246258
rect 67357 245714 67423 245717
rect 70166 245714 70226 246228
rect 119876 246200 121458 246256
rect 121514 246200 121519 246256
rect 119876 246198 121519 246200
rect 121453 246195 121519 246198
rect 67357 245712 70226 245714
rect 67357 245656 67362 245712
rect 67418 245656 70226 245712
rect 67357 245654 70226 245656
rect 67357 245651 67423 245654
rect 121545 245578 121611 245581
rect 119876 245576 121611 245578
rect 69197 245034 69263 245037
rect 70166 245034 70226 245548
rect 119876 245520 121550 245576
rect 121606 245520 121611 245576
rect 119876 245518 121611 245520
rect 121545 245515 121611 245518
rect 579981 245578 580047 245581
rect 583520 245578 584960 245668
rect 579981 245576 584960 245578
rect 579981 245520 579986 245576
rect 580042 245520 584960 245576
rect 579981 245518 584960 245520
rect 579981 245515 580047 245518
rect 583520 245428 584960 245518
rect 69197 245032 70226 245034
rect 69197 244976 69202 245032
rect 69258 244976 70226 245032
rect 69197 244974 70226 244976
rect 69197 244971 69263 244974
rect 121453 244898 121519 244901
rect 119876 244896 121519 244898
rect 67633 244626 67699 244629
rect 70166 244626 70226 244868
rect 119876 244840 121458 244896
rect 121514 244840 121519 244896
rect 119876 244838 121519 244840
rect 121453 244835 121519 244838
rect 67633 244624 70226 244626
rect 67633 244568 67638 244624
rect 67694 244568 70226 244624
rect 67633 244566 70226 244568
rect 67633 244563 67699 244566
rect 121545 244218 121611 244221
rect 119876 244216 121611 244218
rect 67725 243674 67791 243677
rect 70166 243674 70226 244188
rect 119876 244160 121550 244216
rect 121606 244160 121611 244216
rect 119876 244158 121611 244160
rect 121545 244155 121611 244158
rect 67725 243672 70226 243674
rect 67725 243616 67730 243672
rect 67786 243616 70226 243672
rect 67725 243614 70226 243616
rect 67725 243611 67791 243614
rect 121678 243538 121684 243540
rect 67633 243266 67699 243269
rect 70166 243266 70226 243508
rect 119876 243478 121684 243538
rect 121678 243476 121684 243478
rect 121748 243538 121754 243540
rect 122097 243538 122163 243541
rect 121748 243536 122163 243538
rect 121748 243480 122102 243536
rect 122158 243480 122163 243536
rect 121748 243478 122163 243480
rect 121748 243476 121754 243478
rect 122097 243475 122163 243478
rect 67633 243264 70226 243266
rect 67633 243208 67638 243264
rect 67694 243208 70226 243264
rect 67633 243206 70226 243208
rect 67633 243203 67699 243206
rect 121453 242858 121519 242861
rect 119876 242856 121519 242858
rect 69841 242314 69907 242317
rect 70166 242314 70226 242828
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 121453 242795 121519 242798
rect 69841 242312 70226 242314
rect 69841 242256 69846 242312
rect 69902 242256 70226 242312
rect 69841 242254 70226 242256
rect 69841 242251 69907 242254
rect 121545 242178 121611 242181
rect 119876 242176 121611 242178
rect 68185 241634 68251 241637
rect 70166 241634 70226 242148
rect 119876 242120 121550 242176
rect 121606 242120 121611 242176
rect 119876 242118 121611 242120
rect 121545 242115 121611 242118
rect 68185 241632 70226 241634
rect 68185 241576 68190 241632
rect 68246 241576 70226 241632
rect 68185 241574 70226 241576
rect 68185 241571 68251 241574
rect 121637 241498 121703 241501
rect 119876 241496 121703 241498
rect -960 241090 480 241180
rect 3141 241090 3207 241093
rect -960 241088 3207 241090
rect -960 241032 3146 241088
rect 3202 241032 3207 241088
rect -960 241030 3207 241032
rect -960 240940 480 241030
rect 3141 241027 3207 241030
rect 67633 240954 67699 240957
rect 70166 240954 70226 241468
rect 119876 241440 121642 241496
rect 121698 241440 121703 241496
rect 119876 241438 121703 241440
rect 121637 241435 121703 241438
rect 67633 240952 70226 240954
rect 67633 240896 67638 240952
rect 67694 240896 70226 240952
rect 67633 240894 70226 240896
rect 67633 240891 67699 240894
rect 121453 240818 121519 240821
rect 119876 240816 121519 240818
rect 70534 240276 70594 240788
rect 119876 240760 121458 240816
rect 121514 240760 121519 240816
rect 119876 240758 121519 240760
rect 121453 240755 121519 240758
rect 122741 240818 122807 240821
rect 427854 240818 427860 240820
rect 122741 240816 427860 240818
rect 122741 240760 122746 240816
rect 122802 240760 427860 240816
rect 122741 240758 427860 240760
rect 122741 240755 122807 240758
rect 427854 240756 427860 240758
rect 427924 240756 427930 240820
rect 70526 240212 70532 240276
rect 70596 240212 70602 240276
rect 122097 240138 122163 240141
rect 119876 240136 122163 240138
rect 119876 240080 122102 240136
rect 122158 240080 122163 240136
rect 119876 240078 122163 240080
rect 122097 240075 122163 240078
rect 68829 239458 68895 239461
rect 170254 239458 170260 239460
rect 68829 239456 170260 239458
rect 68829 239400 68834 239456
rect 68890 239400 170260 239456
rect 68829 239398 170260 239400
rect 68829 239395 68895 239398
rect 170254 239396 170260 239398
rect 170324 239396 170330 239460
rect 50838 238580 50844 238644
rect 50908 238642 50914 238644
rect 98361 238642 98427 238645
rect 50908 238640 98427 238642
rect 50908 238584 98366 238640
rect 98422 238584 98427 238640
rect 50908 238582 98427 238584
rect 50908 238580 50914 238582
rect 98361 238579 98427 238582
rect 86125 237962 86191 237965
rect 169017 237962 169083 237965
rect 86125 237960 169083 237962
rect 86125 237904 86130 237960
rect 86186 237904 169022 237960
rect 169078 237904 169083 237960
rect 86125 237902 169083 237904
rect 86125 237899 86191 237902
rect 169017 237899 169083 237902
rect 59118 237220 59124 237284
rect 59188 237282 59194 237284
rect 76557 237282 76623 237285
rect 59188 237280 76623 237282
rect 59188 237224 76562 237280
rect 76618 237224 76623 237280
rect 59188 237222 76623 237224
rect 59188 237220 59194 237222
rect 76557 237219 76623 237222
rect 113817 237282 113883 237285
rect 129774 237282 129780 237284
rect 113817 237280 129780 237282
rect 113817 237224 113822 237280
rect 113878 237224 129780 237280
rect 113817 237222 129780 237224
rect 113817 237219 113883 237222
rect 129774 237220 129780 237222
rect 129844 237220 129850 237284
rect 113817 236058 113883 236061
rect 114461 236058 114527 236061
rect 113817 236056 114527 236058
rect 113817 236000 113822 236056
rect 113878 236000 114466 236056
rect 114522 236000 114527 236056
rect 113817 235998 114527 236000
rect 113817 235995 113883 235998
rect 114461 235995 114527 235998
rect 44030 235860 44036 235924
rect 44100 235922 44106 235924
rect 107377 235922 107443 235925
rect 44100 235920 107443 235922
rect 44100 235864 107382 235920
rect 107438 235864 107443 235920
rect 44100 235862 107443 235864
rect 44100 235860 44106 235862
rect 107377 235859 107443 235862
rect 55070 235724 55076 235788
rect 55140 235786 55146 235788
rect 95785 235786 95851 235789
rect 98637 235786 98703 235789
rect 55140 235784 98703 235786
rect 55140 235728 95790 235784
rect 95846 235728 98642 235784
rect 98698 235728 98703 235784
rect 55140 235726 98703 235728
rect 55140 235724 55146 235726
rect 95785 235723 95851 235726
rect 98637 235723 98703 235726
rect 67633 234562 67699 234565
rect 124254 234562 124260 234564
rect 67633 234560 124260 234562
rect 67633 234504 67638 234560
rect 67694 234504 124260 234560
rect 67633 234502 124260 234504
rect 67633 234499 67699 234502
rect 124254 234500 124260 234502
rect 124324 234562 124330 234564
rect 376753 234562 376819 234565
rect 377397 234562 377463 234565
rect 124324 234560 377463 234562
rect 124324 234504 376758 234560
rect 376814 234504 377402 234560
rect 377458 234504 377463 234560
rect 124324 234502 377463 234504
rect 124324 234500 124330 234502
rect 376753 234499 376819 234502
rect 377397 234499 377463 234502
rect 91277 234426 91343 234429
rect 140865 234426 140931 234429
rect 91277 234424 142170 234426
rect 91277 234368 91282 234424
rect 91338 234368 140870 234424
rect 140926 234368 142170 234424
rect 91277 234366 142170 234368
rect 91277 234363 91343 234366
rect 140865 234363 140931 234366
rect 142110 233882 142170 234366
rect 291878 233882 291884 233884
rect 142110 233822 291884 233882
rect 291878 233820 291884 233822
rect 291948 233820 291954 233884
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 69054 231100 69060 231164
rect 69124 231162 69130 231164
rect 430757 231162 430823 231165
rect 69124 231160 430823 231162
rect 69124 231104 430762 231160
rect 430818 231104 430823 231160
rect 69124 231102 430823 231104
rect 69124 231100 69130 231102
rect 430757 231099 430823 231102
rect -960 227884 480 228124
rect 61694 226884 61700 226948
rect 61764 226946 61770 226948
rect 359457 226946 359523 226949
rect 61764 226944 359523 226946
rect 61764 226888 359462 226944
rect 359518 226888 359523 226944
rect 61764 226886 359523 226888
rect 61764 226884 61770 226886
rect 359457 226883 359523 226886
rect 103605 222866 103671 222869
rect 287094 222866 287100 222868
rect 103605 222864 287100 222866
rect 103605 222808 103610 222864
rect 103666 222808 287100 222864
rect 103605 222806 287100 222808
rect 103605 222803 103671 222806
rect 287094 222804 287100 222806
rect 287164 222804 287170 222868
rect 76557 220146 76623 220149
rect 294454 220146 294460 220148
rect 76557 220144 294460 220146
rect 76557 220088 76562 220144
rect 76618 220088 294460 220144
rect 76557 220086 294460 220088
rect 76557 220083 76623 220086
rect 294454 220084 294460 220086
rect 294524 220084 294530 220148
rect 114645 219330 114711 219333
rect 143625 219330 143691 219333
rect 114645 219328 143691 219330
rect 114645 219272 114650 219328
rect 114706 219272 143630 219328
rect 143686 219272 143691 219328
rect 114645 219270 143691 219272
rect 114645 219267 114711 219270
rect 143625 219267 143691 219270
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 143625 218650 143691 218653
rect 293166 218650 293172 218652
rect 143625 218648 293172 218650
rect 143625 218592 143630 218648
rect 143686 218592 293172 218648
rect 143625 218590 293172 218592
rect 143625 218587 143691 218590
rect 293166 218588 293172 218590
rect 293236 218588 293242 218652
rect 70393 216066 70459 216069
rect 233182 216066 233188 216068
rect 70393 216064 233188 216066
rect 70393 216008 70398 216064
rect 70454 216008 233188 216064
rect 70393 216006 233188 216008
rect 70393 216003 70459 216006
rect 233182 216004 233188 216006
rect 233252 216004 233258 216068
rect 87045 215930 87111 215933
rect 287278 215930 287284 215932
rect 87045 215928 287284 215930
rect 87045 215872 87050 215928
rect 87106 215872 287284 215928
rect 87045 215870 287284 215872
rect 87045 215867 87111 215870
rect 287278 215868 287284 215870
rect 287348 215868 287354 215932
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 106273 212530 106339 212533
rect 139393 212530 139459 212533
rect 106273 212528 139459 212530
rect 106273 212472 106278 212528
rect 106334 212472 139398 212528
rect 139454 212472 139459 212528
rect 106273 212470 139459 212472
rect 106273 212467 106339 212470
rect 139393 212467 139459 212470
rect 139393 211850 139459 211853
rect 295926 211850 295932 211852
rect 139393 211848 295932 211850
rect 139393 211792 139398 211848
rect 139454 211792 295932 211848
rect 139393 211790 295932 211792
rect 139393 211787 139459 211790
rect 295926 211788 295932 211790
rect 295996 211788 296002 211852
rect 77385 208994 77451 208997
rect 288382 208994 288388 208996
rect 77385 208992 288388 208994
rect 77385 208936 77390 208992
rect 77446 208936 288388 208992
rect 77385 208934 288388 208936
rect 77385 208931 77451 208934
rect 288382 208932 288388 208934
rect 288452 208932 288458 208996
rect 119337 206274 119403 206277
rect 429142 206274 429148 206276
rect 119337 206272 429148 206274
rect 119337 206216 119342 206272
rect 119398 206216 429148 206272
rect 119337 206214 429148 206216
rect 119337 206211 119403 206214
rect 429142 206212 429148 206214
rect 429212 206212 429218 206276
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 57094 202132 57100 202196
rect 57164 202194 57170 202196
rect 336273 202194 336339 202197
rect 57164 202192 336339 202194
rect 57164 202136 336278 202192
rect 336334 202136 336339 202192
rect 57164 202134 336339 202136
rect 57164 202132 57170 202134
rect 336273 202131 336339 202134
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 68921 199338 68987 199341
rect 280286 199338 280292 199340
rect 68921 199336 280292 199338
rect 68921 199280 68926 199336
rect 68982 199280 280292 199336
rect 68921 199278 280292 199280
rect 68921 199275 68987 199278
rect 280286 199276 280292 199278
rect 280356 199276 280362 199340
rect 133137 198114 133203 198117
rect 238518 198114 238524 198116
rect 133137 198112 238524 198114
rect 133137 198056 133142 198112
rect 133198 198056 238524 198112
rect 133137 198054 238524 198056
rect 133137 198051 133203 198054
rect 238518 198052 238524 198054
rect 238588 198052 238594 198116
rect 155309 197978 155375 197981
rect 290590 197978 290596 197980
rect 155309 197976 290596 197978
rect 155309 197920 155314 197976
rect 155370 197920 290596 197976
rect 155309 197918 290596 197920
rect 155309 197915 155375 197918
rect 290590 197916 290596 197918
rect 290660 197916 290666 197980
rect 66110 196556 66116 196620
rect 66180 196618 66186 196620
rect 281625 196618 281691 196621
rect 66180 196616 281691 196618
rect 66180 196560 281630 196616
rect 281686 196560 281691 196616
rect 66180 196558 281691 196560
rect 66180 196556 66186 196558
rect 281625 196555 281691 196558
rect 56501 195258 56567 195261
rect 237414 195258 237420 195260
rect 56501 195256 237420 195258
rect 56501 195200 56506 195256
rect 56562 195200 237420 195256
rect 56501 195198 237420 195200
rect 56501 195195 56567 195198
rect 237414 195196 237420 195198
rect 237484 195196 237490 195260
rect 84285 192538 84351 192541
rect 284334 192538 284340 192540
rect 84285 192536 284340 192538
rect 84285 192480 84290 192536
rect 84346 192480 284340 192536
rect 84285 192478 284340 192480
rect 84285 192475 84351 192478
rect 284334 192476 284340 192478
rect 284404 192476 284410 192540
rect 580901 192538 580967 192541
rect 583520 192538 584960 192628
rect 580901 192536 584960 192538
rect 580901 192480 580906 192536
rect 580962 192480 584960 192536
rect 580901 192478 584960 192480
rect 580901 192475 580967 192478
rect 583520 192388 584960 192478
rect 53465 191042 53531 191045
rect 394693 191042 394759 191045
rect 53465 191040 394759 191042
rect 53465 190984 53470 191040
rect 53526 190984 394698 191040
rect 394754 190984 394759 191040
rect 53465 190982 394759 190984
rect 53465 190979 53531 190982
rect 394693 190979 394759 190982
rect 224309 189682 224375 189685
rect 298134 189682 298140 189684
rect 224309 189680 298140 189682
rect 224309 189624 224314 189680
rect 224370 189624 298140 189680
rect 224309 189622 298140 189624
rect 224309 189619 224375 189622
rect 298134 189620 298140 189622
rect 298204 189620 298210 189684
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 147581 188322 147647 188325
rect 344277 188322 344343 188325
rect 147581 188320 344343 188322
rect 147581 188264 147586 188320
rect 147642 188264 344282 188320
rect 344338 188264 344343 188320
rect 147581 188262 344343 188264
rect 147581 188259 147647 188262
rect 344277 188259 344343 188262
rect 349102 188260 349108 188324
rect 349172 188322 349178 188324
rect 580257 188322 580323 188325
rect 349172 188320 580323 188322
rect 349172 188264 580262 188320
rect 580318 188264 580323 188320
rect 349172 188262 580323 188264
rect 349172 188260 349178 188262
rect 580257 188259 580323 188262
rect 211797 186962 211863 186965
rect 244222 186962 244228 186964
rect 211797 186960 244228 186962
rect 211797 186904 211802 186960
rect 211858 186904 244228 186960
rect 211797 186902 244228 186904
rect 211797 186899 211863 186902
rect 244222 186900 244228 186902
rect 244292 186900 244298 186964
rect 74533 185602 74599 185605
rect 233366 185602 233372 185604
rect 74533 185600 233372 185602
rect 74533 185544 74538 185600
rect 74594 185544 233372 185600
rect 74533 185542 233372 185544
rect 74533 185539 74599 185542
rect 233366 185540 233372 185542
rect 233436 185540 233442 185604
rect 78673 182882 78739 182885
rect 245878 182882 245884 182884
rect 78673 182880 245884 182882
rect 78673 182824 78678 182880
rect 78734 182824 245884 182880
rect 78673 182822 245884 182824
rect 78673 182819 78739 182822
rect 245878 182820 245884 182822
rect 245948 182820 245954 182884
rect 41321 181386 41387 181389
rect 199469 181386 199535 181389
rect 41321 181384 199535 181386
rect 41321 181328 41326 181384
rect 41382 181328 199474 181384
rect 199530 181328 199535 181384
rect 41321 181326 199535 181328
rect 41321 181323 41387 181326
rect 199469 181323 199535 181326
rect 70894 180100 70900 180164
rect 70964 180162 70970 180164
rect 203609 180162 203675 180165
rect 70964 180160 203675 180162
rect 70964 180104 203614 180160
rect 203670 180104 203675 180160
rect 70964 180102 203675 180104
rect 70964 180100 70970 180102
rect 203609 180099 203675 180102
rect 63309 180026 63375 180029
rect 231894 180026 231900 180028
rect 63309 180024 231900 180026
rect 63309 179968 63314 180024
rect 63370 179968 231900 180024
rect 63309 179966 231900 179968
rect 63309 179963 63375 179966
rect 231894 179964 231900 179966
rect 231964 179964 231970 180028
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 166257 178666 166323 178669
rect 180057 178666 180123 178669
rect 166257 178664 180123 178666
rect 166257 178608 166262 178664
rect 166318 178608 180062 178664
rect 180118 178608 180123 178664
rect 166257 178606 180123 178608
rect 166257 178603 166323 178606
rect 180057 178603 180123 178606
rect 218697 178666 218763 178669
rect 237598 178666 237604 178668
rect 218697 178664 237604 178666
rect 218697 178608 218702 178664
rect 218758 178608 237604 178664
rect 218697 178606 237604 178608
rect 218697 178603 218763 178606
rect 237598 178604 237604 178606
rect 237668 178604 237674 178668
rect 269941 178666 270007 178669
rect 278998 178666 279004 178668
rect 269941 178664 279004 178666
rect 269941 178608 269946 178664
rect 270002 178608 279004 178664
rect 269941 178606 279004 178608
rect 269941 178603 270007 178606
rect 278998 178604 279004 178606
rect 279068 178604 279074 178668
rect 221549 177850 221615 177853
rect 228950 177850 228956 177852
rect 221549 177848 228956 177850
rect 221549 177792 221554 177848
rect 221610 177792 228956 177848
rect 221549 177790 228956 177792
rect 221549 177787 221615 177790
rect 228950 177788 228956 177790
rect 229020 177788 229026 177852
rect 104566 177652 104572 177716
rect 104636 177714 104642 177716
rect 104801 177714 104867 177717
rect 104636 177712 104867 177714
rect 104636 177656 104806 177712
rect 104862 177656 104867 177712
rect 104636 177654 104867 177656
rect 104636 177652 104642 177654
rect 104801 177651 104867 177654
rect 105670 177652 105676 177716
rect 105740 177714 105746 177716
rect 106181 177714 106247 177717
rect 105740 177712 106247 177714
rect 105740 177656 106186 177712
rect 106242 177656 106247 177712
rect 105740 177654 106247 177656
rect 105740 177652 105746 177654
rect 106181 177651 106247 177654
rect 108062 177652 108068 177716
rect 108132 177714 108138 177716
rect 108941 177714 109007 177717
rect 116945 177716 117011 177717
rect 119521 177716 119587 177717
rect 116894 177714 116900 177716
rect 108132 177712 109007 177714
rect 108132 177656 108946 177712
rect 109002 177656 109007 177712
rect 108132 177654 109007 177656
rect 116854 177654 116900 177714
rect 116964 177712 117011 177716
rect 119470 177714 119476 177716
rect 117006 177656 117011 177712
rect 108132 177652 108138 177654
rect 108941 177651 109007 177654
rect 116894 177652 116900 177654
rect 116964 177652 117011 177656
rect 119430 177654 119476 177714
rect 119540 177712 119587 177716
rect 119582 177656 119587 177712
rect 119470 177652 119476 177654
rect 119540 177652 119587 177656
rect 121862 177652 121868 177716
rect 121932 177714 121938 177716
rect 122005 177714 122071 177717
rect 121932 177712 122071 177714
rect 121932 177656 122010 177712
rect 122066 177656 122071 177712
rect 121932 177654 122071 177656
rect 121932 177652 121938 177654
rect 116945 177651 117011 177652
rect 119521 177651 119587 177652
rect 122005 177651 122071 177654
rect 129406 177652 129412 177716
rect 129476 177714 129482 177716
rect 129641 177714 129707 177717
rect 129476 177712 129707 177714
rect 129476 177656 129646 177712
rect 129702 177656 129707 177712
rect 129476 177654 129707 177656
rect 129476 177652 129482 177654
rect 129641 177651 129707 177654
rect 130694 177652 130700 177716
rect 130764 177714 130770 177716
rect 131021 177714 131087 177717
rect 132401 177716 132467 177717
rect 132350 177714 132356 177716
rect 130764 177712 131087 177714
rect 130764 177656 131026 177712
rect 131082 177656 131087 177712
rect 130764 177654 131087 177656
rect 132310 177654 132356 177714
rect 132420 177712 132467 177716
rect 132462 177656 132467 177712
rect 130764 177652 130770 177654
rect 131021 177651 131087 177654
rect 132350 177652 132356 177654
rect 132420 177652 132467 177656
rect 132401 177651 132467 177652
rect 226977 177442 227043 177445
rect 234654 177442 234660 177444
rect 226977 177440 234660 177442
rect 226977 177384 226982 177440
rect 227038 177384 234660 177440
rect 226977 177382 234660 177384
rect 226977 177379 227043 177382
rect 234654 177380 234660 177382
rect 234724 177380 234730 177444
rect 276657 177442 276723 177445
rect 288566 177442 288572 177444
rect 276657 177440 288572 177442
rect 276657 177384 276662 177440
rect 276718 177384 288572 177440
rect 276657 177382 288572 177384
rect 276657 177379 276723 177382
rect 288566 177380 288572 177382
rect 288636 177380 288642 177444
rect 213269 177306 213335 177309
rect 240542 177306 240548 177308
rect 213269 177304 240548 177306
rect 213269 177248 213274 177304
rect 213330 177248 240548 177304
rect 213269 177246 240548 177248
rect 213269 177243 213335 177246
rect 240542 177244 240548 177246
rect 240612 177244 240618 177308
rect 260097 177306 260163 177309
rect 291694 177306 291700 177308
rect 260097 177304 291700 177306
rect 260097 177248 260102 177304
rect 260158 177248 291700 177304
rect 260097 177246 291700 177248
rect 260097 177243 260163 177246
rect 291694 177244 291700 177246
rect 291764 177244 291770 177308
rect 115841 177172 115907 177173
rect 115790 177170 115796 177172
rect 115750 177110 115796 177170
rect 115860 177168 115907 177172
rect 115902 177112 115907 177168
rect 115790 177108 115796 177110
rect 115860 177108 115907 177112
rect 120758 177108 120764 177172
rect 120828 177170 120834 177172
rect 120993 177170 121059 177173
rect 133137 177172 133203 177173
rect 133086 177170 133092 177172
rect 120828 177168 121059 177170
rect 120828 177112 120998 177168
rect 121054 177112 121059 177168
rect 120828 177110 121059 177112
rect 133046 177110 133092 177170
rect 133156 177168 133203 177172
rect 133198 177112 133203 177168
rect 120828 177108 120834 177110
rect 115841 177107 115907 177108
rect 120993 177107 121059 177110
rect 133086 177108 133092 177110
rect 133156 177108 133203 177112
rect 133137 177107 133203 177108
rect 97022 176972 97028 177036
rect 97092 177034 97098 177036
rect 97349 177034 97415 177037
rect 97092 177032 97415 177034
rect 97092 176976 97354 177032
rect 97410 176976 97415 177032
rect 97092 176974 97415 176976
rect 97092 176972 97098 176974
rect 97349 176971 97415 176974
rect 100702 176972 100708 177036
rect 100772 177034 100778 177036
rect 168230 177034 168236 177036
rect 100772 176974 168236 177034
rect 100772 176972 100778 176974
rect 168230 176972 168236 176974
rect 168300 176972 168306 177036
rect 106958 176836 106964 176900
rect 107028 176898 107034 176900
rect 107028 176838 110890 176898
rect 107028 176836 107034 176838
rect 100661 176762 100727 176765
rect 102041 176764 102107 176765
rect 101990 176762 101996 176764
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 101950 176702 101996 176762
rect 102060 176760 102107 176764
rect 103421 176762 103487 176765
rect 102102 176704 102107 176760
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 101990 176700 101996 176702
rect 102060 176700 102107 176704
rect 102041 176699 102107 176700
rect 103286 176760 103487 176762
rect 103286 176704 103426 176760
rect 103482 176704 103487 176760
rect 103286 176702 103487 176704
rect 103286 176492 103346 176702
rect 103421 176699 103487 176702
rect 109534 176700 109540 176764
rect 109604 176762 109610 176764
rect 109769 176762 109835 176765
rect 110689 176764 110755 176765
rect 110638 176762 110644 176764
rect 109604 176760 109835 176762
rect 109604 176704 109774 176760
rect 109830 176704 109835 176760
rect 109604 176702 109835 176704
rect 110598 176702 110644 176762
rect 110708 176760 110755 176764
rect 110750 176704 110755 176760
rect 109604 176700 109610 176702
rect 109769 176699 109835 176702
rect 110638 176700 110644 176702
rect 110708 176700 110755 176704
rect 110830 176762 110890 176838
rect 112110 176836 112116 176900
rect 112180 176898 112186 176900
rect 112253 176898 112319 176901
rect 166206 176898 166212 176900
rect 112180 176896 112319 176898
rect 112180 176840 112258 176896
rect 112314 176840 112319 176896
rect 112180 176838 112319 176840
rect 112180 176836 112186 176838
rect 112253 176835 112319 176838
rect 113130 176838 166212 176898
rect 113130 176762 113190 176838
rect 166206 176836 166212 176838
rect 166276 176836 166282 176900
rect 114369 176764 114435 176765
rect 118417 176764 118483 176765
rect 124489 176764 124555 176765
rect 125777 176764 125843 176765
rect 127065 176764 127131 176765
rect 134425 176764 134491 176765
rect 148225 176764 148291 176765
rect 114318 176762 114324 176764
rect 110830 176702 113190 176762
rect 114278 176702 114324 176762
rect 114388 176760 114435 176764
rect 118366 176762 118372 176764
rect 114430 176704 114435 176760
rect 114318 176700 114324 176702
rect 114388 176700 114435 176704
rect 118326 176702 118372 176762
rect 118436 176760 118483 176764
rect 124438 176762 124444 176764
rect 118478 176704 118483 176760
rect 118366 176700 118372 176702
rect 118436 176700 118483 176704
rect 124398 176702 124444 176762
rect 124508 176760 124555 176764
rect 125726 176762 125732 176764
rect 124550 176704 124555 176760
rect 124438 176700 124444 176702
rect 124508 176700 124555 176704
rect 125686 176702 125732 176762
rect 125796 176760 125843 176764
rect 127014 176762 127020 176764
rect 125838 176704 125843 176760
rect 125726 176700 125732 176702
rect 125796 176700 125843 176704
rect 126974 176702 127020 176762
rect 127084 176760 127131 176764
rect 134374 176762 134380 176764
rect 127126 176704 127131 176760
rect 127014 176700 127020 176702
rect 127084 176700 127131 176704
rect 134334 176702 134380 176762
rect 134444 176760 134491 176764
rect 148174 176762 148180 176764
rect 134486 176704 134491 176760
rect 134374 176700 134380 176702
rect 134444 176700 134491 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 110689 176699 110755 176700
rect 114369 176699 114435 176700
rect 118417 176699 118483 176700
rect 124489 176699 124555 176700
rect 125777 176699 125843 176700
rect 127065 176699 127131 176700
rect 134425 176699 134491 176700
rect 148225 176699 148291 176700
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 227069 176354 227135 176357
rect 229093 176354 229159 176357
rect 227069 176352 229159 176354
rect 227069 176296 227074 176352
rect 227130 176296 229098 176352
rect 229154 176296 229159 176352
rect 227069 176294 229159 176296
rect 227069 176291 227135 176294
rect 229093 176291 229159 176294
rect 425697 176082 425763 176085
rect 435030 176082 435036 176084
rect 425697 176080 435036 176082
rect -960 175796 480 176036
rect 425697 176024 425702 176080
rect 425758 176024 435036 176080
rect 425697 176022 435036 176024
rect 425697 176019 425763 176022
rect 435030 176020 435036 176022
rect 435100 176020 435106 176084
rect 109401 175946 109467 175949
rect 440417 175946 440483 175949
rect 109401 175944 440483 175946
rect 109401 175888 109406 175944
rect 109462 175888 440422 175944
rect 440478 175888 440483 175944
rect 109401 175886 440483 175888
rect 109401 175883 109467 175886
rect 440417 175883 440483 175886
rect 213913 175810 213979 175813
rect 227713 175810 227779 175813
rect 278313 175810 278379 175813
rect 279325 175810 279391 175813
rect 213913 175808 217242 175810
rect 213913 175752 213918 175808
rect 213974 175752 217242 175808
rect 213913 175750 217242 175752
rect 213913 175747 213979 175750
rect 217182 175644 217242 175750
rect 227713 175808 228282 175810
rect 227713 175752 227718 175808
rect 227774 175752 228282 175808
rect 227713 175750 228282 175752
rect 227713 175747 227779 175750
rect 228222 175644 228282 175750
rect 278313 175808 279391 175810
rect 278313 175752 278318 175808
rect 278374 175752 279330 175808
rect 279386 175752 279391 175808
rect 278313 175750 279391 175752
rect 278313 175747 278379 175750
rect 279325 175747 279391 175750
rect 279509 175810 279575 175813
rect 279509 175808 279618 175810
rect 279509 175752 279514 175808
rect 279570 175752 279618 175808
rect 279509 175747 279618 175752
rect 135713 175540 135779 175541
rect 135662 175538 135668 175540
rect 135622 175478 135668 175538
rect 135732 175536 135779 175540
rect 135774 175480 135779 175536
rect 135662 175476 135668 175478
rect 135732 175476 135779 175480
rect 135713 175475 135779 175476
rect 98361 175404 98427 175405
rect 128169 175404 128235 175405
rect 158897 175404 158963 175405
rect 98310 175402 98316 175404
rect 98270 175342 98316 175402
rect 98380 175400 98427 175404
rect 128118 175402 128124 175404
rect 98422 175344 98427 175400
rect 98310 175340 98316 175342
rect 98380 175340 98427 175344
rect 128078 175342 128124 175402
rect 128188 175400 128235 175404
rect 158846 175402 158852 175404
rect 128230 175344 128235 175400
rect 128118 175340 128124 175342
rect 128188 175340 128235 175344
rect 158806 175342 158852 175402
rect 158916 175400 158963 175404
rect 158958 175344 158963 175400
rect 158846 175340 158852 175342
rect 158916 175340 158963 175344
rect 98361 175339 98427 175340
rect 128169 175339 128235 175340
rect 158897 175339 158963 175340
rect 264421 175402 264487 175405
rect 268150 175402 268210 175644
rect 279558 175508 279618 175747
rect 264421 175400 268210 175402
rect 264421 175344 264426 175400
rect 264482 175344 268210 175400
rect 264421 175342 268210 175344
rect 264421 175339 264487 175342
rect 229134 175266 229140 175268
rect 228968 175206 229140 175266
rect 229134 175204 229140 175206
rect 229204 175204 229210 175268
rect 279417 175266 279483 175269
rect 279374 175264 279483 175266
rect 213913 175130 213979 175133
rect 213913 175128 217242 175130
rect 213913 175072 213918 175128
rect 213974 175072 217242 175128
rect 213913 175070 217242 175072
rect 213913 175067 213979 175070
rect 113173 174996 113239 174997
rect 123109 174996 123175 174997
rect 113136 174932 113142 174996
rect 113206 174994 113239 174996
rect 123064 174994 123070 174996
rect 113206 174992 113298 174994
rect 113234 174936 113298 174992
rect 113206 174934 113298 174936
rect 123018 174934 123070 174994
rect 123134 174992 123175 174996
rect 123170 174936 123175 174992
rect 217182 174964 217242 175070
rect 265893 174994 265959 174997
rect 268150 174994 268210 175236
rect 265893 174992 268210 174994
rect 113206 174932 113239 174934
rect 123064 174932 123070 174934
rect 123134 174932 123175 174936
rect 113173 174931 113239 174932
rect 123109 174931 123175 174932
rect 265893 174936 265898 174992
rect 265954 174936 268210 174992
rect 265893 174934 268210 174936
rect 279374 175208 279422 175264
rect 279478 175208 279483 175264
rect 279374 175203 279483 175208
rect 427813 175266 427879 175269
rect 427813 175264 427922 175266
rect 427813 175208 427818 175264
rect 427874 175208 427922 175264
rect 427813 175203 427922 175208
rect 265893 174931 265959 174934
rect 214005 174722 214071 174725
rect 229134 174722 229140 174724
rect 214005 174720 217242 174722
rect 214005 174664 214010 174720
rect 214066 174664 217242 174720
rect 214005 174662 217242 174664
rect 228968 174662 229140 174722
rect 214005 174659 214071 174662
rect 217182 174284 217242 174662
rect 229134 174660 229140 174662
rect 229204 174660 229210 174724
rect 265985 174586 266051 174589
rect 268150 174586 268210 174828
rect 279374 174692 279434 175203
rect 427862 174964 427922 175203
rect 347497 174722 347563 174725
rect 347497 174720 350060 174722
rect 347497 174664 347502 174720
rect 347558 174664 350060 174720
rect 347497 174662 350060 174664
rect 347497 174659 347563 174662
rect 265985 174584 268210 174586
rect 265985 174528 265990 174584
rect 266046 174528 268210 174584
rect 265985 174526 268210 174528
rect 265985 174523 266051 174526
rect 279325 174450 279391 174453
rect 279325 174448 279434 174450
rect 229093 174314 229159 174317
rect 228968 174312 229159 174314
rect 228968 174256 229098 174312
rect 229154 174256 229159 174312
rect 228968 174254 229159 174256
rect 229093 174251 229159 174254
rect 265341 174178 265407 174181
rect 268150 174178 268210 174420
rect 279325 174392 279330 174448
rect 279386 174392 279434 174448
rect 279325 174387 279434 174392
rect 265341 174176 268210 174178
rect 265341 174120 265346 174176
rect 265402 174120 268210 174176
rect 265341 174118 268210 174120
rect 265341 174115 265407 174118
rect 265801 174042 265867 174045
rect 265801 174040 267842 174042
rect 265801 173984 265806 174040
rect 265862 173984 267842 174040
rect 279374 174012 279434 174387
rect 265801 173982 267842 173984
rect 265801 173979 265867 173982
rect 213913 173770 213979 173773
rect 229553 173770 229619 173773
rect 213913 173768 217242 173770
rect 213913 173712 213918 173768
rect 213974 173712 217242 173768
rect 213913 173710 217242 173712
rect 228968 173768 229619 173770
rect 228968 173712 229558 173768
rect 229614 173712 229619 173768
rect 228968 173710 229619 173712
rect 267782 173770 267842 173982
rect 268334 173770 268394 174012
rect 267782 173710 268394 173770
rect 213913 173707 213979 173710
rect 217182 173604 217242 173710
rect 229553 173707 229619 173710
rect 279366 173708 279372 173772
rect 279436 173708 279442 173772
rect 214005 173362 214071 173365
rect 231393 173362 231459 173365
rect 214005 173360 217242 173362
rect 214005 173304 214010 173360
rect 214066 173304 217242 173360
rect 214005 173302 217242 173304
rect 228968 173360 231459 173362
rect 228968 173304 231398 173360
rect 231454 173304 231459 173360
rect 228968 173302 231459 173304
rect 214005 173299 214071 173302
rect 217182 172924 217242 173302
rect 231393 173299 231459 173302
rect 265249 173226 265315 173229
rect 268150 173226 268210 173604
rect 265249 173224 268210 173226
rect 265249 173168 265254 173224
rect 265310 173168 268210 173224
rect 279374 173196 279434 173708
rect 428230 173362 428290 173876
rect 429193 173362 429259 173365
rect 428230 173360 429259 173362
rect 428230 173304 429198 173360
rect 429254 173304 429259 173360
rect 428230 173302 429259 173304
rect 429193 173299 429259 173302
rect 430573 173226 430639 173229
rect 428230 173224 430639 173226
rect 265249 173166 268210 173168
rect 428230 173168 430578 173224
rect 430634 173168 430639 173224
rect 428230 173166 430639 173168
rect 265249 173163 265315 173166
rect 347497 173090 347563 173093
rect 347497 173088 350060 173090
rect 229461 172818 229527 172821
rect 228968 172816 229527 172818
rect 228968 172760 229466 172816
rect 229522 172760 229527 172816
rect 228968 172758 229527 172760
rect 229461 172755 229527 172758
rect 265341 172818 265407 172821
rect 268150 172818 268210 173060
rect 347497 173032 347502 173088
rect 347558 173032 350060 173088
rect 347497 173030 350060 173032
rect 347497 173027 347563 173030
rect 265341 172816 268210 172818
rect 265341 172760 265346 172816
rect 265402 172760 268210 172816
rect 428230 172788 428290 173166
rect 430573 173163 430639 173166
rect 265341 172758 268210 172760
rect 265341 172755 265407 172758
rect 265801 172546 265867 172549
rect 265801 172544 267842 172546
rect 265801 172488 265806 172544
rect 265862 172488 267842 172544
rect 265801 172486 267842 172488
rect 265801 172483 265867 172486
rect 213913 172410 213979 172413
rect 231761 172410 231827 172413
rect 213913 172408 217242 172410
rect 213913 172352 213918 172408
rect 213974 172352 217242 172408
rect 213913 172350 217242 172352
rect 228968 172408 231827 172410
rect 228968 172352 231766 172408
rect 231822 172352 231827 172408
rect 228968 172350 231827 172352
rect 267782 172410 267842 172486
rect 268334 172410 268394 172652
rect 281533 172410 281599 172413
rect 267782 172350 268394 172410
rect 279956 172408 281599 172410
rect 279956 172352 281538 172408
rect 281594 172352 281599 172408
rect 279956 172350 281599 172352
rect 213913 172347 213979 172350
rect 217182 172244 217242 172350
rect 231761 172347 231827 172350
rect 281533 172347 281599 172350
rect 429377 172274 429443 172277
rect 428230 172272 429443 172274
rect 214097 172002 214163 172005
rect 265065 172002 265131 172005
rect 268150 172002 268210 172244
rect 214097 172000 217242 172002
rect 214097 171944 214102 172000
rect 214158 171944 217242 172000
rect 214097 171942 217242 171944
rect 214097 171939 214163 171942
rect 167085 171594 167151 171597
rect 164694 171592 167151 171594
rect 164694 171536 167090 171592
rect 167146 171536 167151 171592
rect 217182 171564 217242 171942
rect 265065 172000 268210 172002
rect 265065 171944 265070 172000
rect 265126 171944 268210 172000
rect 265065 171942 268210 171944
rect 428230 172216 429382 172272
rect 429438 172216 429443 172272
rect 428230 172214 429443 172216
rect 265065 171939 265131 171942
rect 229369 171866 229435 171869
rect 228968 171864 229435 171866
rect 228968 171808 229374 171864
rect 229430 171808 229435 171864
rect 228968 171806 229435 171808
rect 229369 171803 229435 171806
rect 265157 171594 265223 171597
rect 268150 171594 268210 171836
rect 428230 171700 428290 172214
rect 429377 172211 429443 172214
rect 265157 171592 268210 171594
rect 164694 171534 167151 171536
rect 167085 171531 167151 171534
rect 265157 171536 265162 171592
rect 265218 171536 268210 171592
rect 265157 171534 268210 171536
rect 265157 171531 265223 171534
rect 231669 171458 231735 171461
rect 228968 171456 231735 171458
rect 228968 171400 231674 171456
rect 231730 171400 231735 171456
rect 228968 171398 231735 171400
rect 231669 171395 231735 171398
rect 265341 171186 265407 171189
rect 268150 171186 268210 171428
rect 216998 171126 217242 171186
rect 216998 171050 217058 171126
rect 215250 170990 217058 171050
rect 217182 171020 217242 171126
rect 265341 171184 268210 171186
rect 265341 171128 265346 171184
rect 265402 171128 268210 171184
rect 265341 171126 268210 171128
rect 279926 171186 279986 171700
rect 347497 171322 347563 171325
rect 347497 171320 350060 171322
rect 347497 171264 347502 171320
rect 347558 171264 350060 171320
rect 347497 171262 350060 171264
rect 347497 171259 347563 171262
rect 288566 171186 288572 171188
rect 279926 171126 288572 171186
rect 265341 171123 265407 171126
rect 288566 171124 288572 171126
rect 288636 171124 288642 171188
rect 429377 171186 429443 171189
rect 434846 171186 434852 171188
rect 429377 171184 434852 171186
rect 429377 171128 429382 171184
rect 429438 171128 434852 171184
rect 429377 171126 434852 171128
rect 429377 171123 429443 171126
rect 434846 171124 434852 171126
rect 434916 171124 434922 171188
rect 214005 170914 214071 170917
rect 215250 170914 215310 170990
rect 231669 170914 231735 170917
rect 214005 170912 215310 170914
rect 214005 170856 214010 170912
rect 214066 170856 215310 170912
rect 214005 170854 215310 170856
rect 228968 170912 231735 170914
rect 228968 170856 231674 170912
rect 231730 170856 231735 170912
rect 228968 170854 231735 170856
rect 214005 170851 214071 170854
rect 231669 170851 231735 170854
rect 213913 170778 213979 170781
rect 213913 170776 217242 170778
rect 213913 170720 213918 170776
rect 213974 170720 217242 170776
rect 213913 170718 217242 170720
rect 213913 170715 213979 170718
rect 217182 170340 217242 170718
rect 265433 170642 265499 170645
rect 268150 170642 268210 171020
rect 282821 170914 282887 170917
rect 279956 170912 282887 170914
rect 279956 170856 282826 170912
rect 282882 170856 282887 170912
rect 279956 170854 282887 170856
rect 282821 170851 282887 170854
rect 265433 170640 268210 170642
rect 265433 170584 265438 170640
rect 265494 170584 268210 170640
rect 265433 170582 268210 170584
rect 265433 170579 265499 170582
rect 231761 170506 231827 170509
rect 228968 170504 231827 170506
rect 228968 170448 231766 170504
rect 231822 170448 231827 170504
rect 228968 170446 231827 170448
rect 231761 170443 231827 170446
rect 265249 170234 265315 170237
rect 268150 170234 268210 170476
rect 265249 170232 268210 170234
rect 265249 170176 265254 170232
rect 265310 170176 268210 170232
rect 265249 170174 268210 170176
rect 265249 170171 265315 170174
rect 282729 170098 282795 170101
rect 279956 170096 282795 170098
rect 231761 169962 231827 169965
rect 228968 169960 231827 169962
rect 228968 169904 231766 169960
rect 231822 169904 231827 169960
rect 228968 169902 231827 169904
rect 231761 169899 231827 169902
rect 265617 169826 265683 169829
rect 268150 169826 268210 170068
rect 279956 170040 282734 170096
rect 282790 170040 282795 170096
rect 279956 170038 282795 170040
rect 282729 170035 282795 170038
rect 428230 169962 428290 170476
rect 430665 169962 430731 169965
rect 432045 169962 432111 169965
rect 428230 169960 432111 169962
rect 428230 169904 430670 169960
rect 430726 169904 432050 169960
rect 432106 169904 432111 169960
rect 428230 169902 432111 169904
rect 430665 169899 430731 169902
rect 432045 169899 432111 169902
rect 216998 169766 217242 169826
rect 213913 169690 213979 169693
rect 216998 169690 217058 169766
rect 213913 169688 217058 169690
rect 213913 169632 213918 169688
rect 213974 169632 217058 169688
rect 217182 169660 217242 169766
rect 265617 169824 268210 169826
rect 265617 169768 265622 169824
rect 265678 169768 268210 169824
rect 265617 169766 268210 169768
rect 265617 169763 265683 169766
rect 347037 169690 347103 169693
rect 347037 169688 350060 169690
rect 213913 169630 217058 169632
rect 213913 169627 213979 169630
rect 231761 169554 231827 169557
rect 228968 169552 231827 169554
rect 228968 169496 231766 169552
rect 231822 169496 231827 169552
rect 228968 169494 231827 169496
rect 231761 169491 231827 169494
rect 214005 169418 214071 169421
rect 265893 169418 265959 169421
rect 268150 169418 268210 169660
rect 347037 169632 347042 169688
rect 347098 169632 350060 169688
rect 347037 169630 350060 169632
rect 347037 169627 347103 169630
rect 281901 169418 281967 169421
rect 214005 169416 217242 169418
rect 214005 169360 214010 169416
rect 214066 169360 217242 169416
rect 214005 169358 217242 169360
rect 214005 169355 214071 169358
rect 217182 168980 217242 169358
rect 265893 169416 268210 169418
rect 265893 169360 265898 169416
rect 265954 169360 268210 169416
rect 265893 169358 268210 169360
rect 279956 169416 281967 169418
rect 279956 169360 281906 169416
rect 281962 169360 281967 169416
rect 279956 169358 281967 169360
rect 265893 169355 265959 169358
rect 281901 169355 281967 169358
rect 231669 169010 231735 169013
rect 228968 169008 231735 169010
rect 228968 168952 231674 169008
rect 231730 168952 231735 169008
rect 228968 168950 231735 168952
rect 231669 168947 231735 168950
rect 265433 169010 265499 169013
rect 268150 169010 268210 169252
rect 265433 169008 268210 169010
rect 265433 168952 265438 169008
rect 265494 168952 268210 169008
rect 265433 168950 268210 168952
rect 265433 168947 265499 168950
rect 428230 168874 428290 169388
rect 429285 168874 429351 168877
rect 430798 168874 430804 168876
rect 428230 168872 430804 168874
rect 231393 168602 231459 168605
rect 228968 168600 231459 168602
rect 228968 168544 231398 168600
rect 231454 168544 231459 168600
rect 228968 168542 231459 168544
rect 231393 168539 231459 168542
rect 265341 168602 265407 168605
rect 268150 168602 268210 168844
rect 428230 168816 429290 168872
rect 429346 168816 430804 168872
rect 428230 168814 430804 168816
rect 429285 168811 429351 168814
rect 430798 168812 430804 168814
rect 430868 168812 430874 168876
rect 281625 168602 281691 168605
rect 265341 168600 268210 168602
rect 265341 168544 265346 168600
rect 265402 168544 268210 168600
rect 265341 168542 268210 168544
rect 279956 168600 281691 168602
rect 279956 168544 281630 168600
rect 281686 168544 281691 168600
rect 279956 168542 281691 168544
rect 265341 168539 265407 168542
rect 281625 168539 281691 168542
rect 265801 168466 265867 168469
rect 216998 168406 217242 168466
rect 213913 168330 213979 168333
rect 216998 168330 217058 168406
rect 213913 168328 217058 168330
rect 213913 168272 213918 168328
rect 213974 168272 217058 168328
rect 217182 168300 217242 168406
rect 265801 168464 267842 168466
rect 265801 168408 265806 168464
rect 265862 168408 267842 168464
rect 265801 168406 267842 168408
rect 265801 168403 265867 168406
rect 238753 168332 238819 168333
rect 213913 168270 217058 168272
rect 213913 168267 213979 168270
rect 238702 168268 238708 168332
rect 238772 168330 238819 168332
rect 238772 168328 238864 168330
rect 238814 168272 238864 168328
rect 238772 168270 238864 168272
rect 238772 168268 238819 168270
rect 238753 168267 238819 168268
rect 267782 168194 267842 168406
rect 268334 168194 268394 168436
rect 267782 168134 268394 168194
rect 214005 168058 214071 168061
rect 231761 168058 231827 168061
rect 214005 168056 217242 168058
rect 214005 168000 214010 168056
rect 214066 168000 217242 168056
rect 214005 167998 217242 168000
rect 228968 168056 231827 168058
rect 228968 168000 231766 168056
rect 231822 168000 231827 168056
rect 228968 167998 231827 168000
rect 214005 167995 214071 167998
rect 217182 167620 217242 167998
rect 231761 167995 231827 167998
rect 347497 167922 347563 167925
rect 347497 167920 350060 167922
rect 240542 167650 240548 167652
rect 228968 167590 240548 167650
rect 240542 167588 240548 167590
rect 240612 167588 240618 167652
rect 265249 167650 265315 167653
rect 268150 167650 268210 167892
rect 347497 167864 347502 167920
rect 347558 167864 350060 167920
rect 347497 167862 350060 167864
rect 347497 167859 347563 167862
rect 281901 167786 281967 167789
rect 279956 167784 281967 167786
rect 279956 167728 281906 167784
rect 281962 167728 281967 167784
rect 279956 167726 281967 167728
rect 428230 167786 428290 168300
rect 429285 167786 429351 167789
rect 428230 167784 429351 167786
rect 428230 167728 429290 167784
rect 429346 167728 429351 167784
rect 428230 167726 429351 167728
rect 281901 167723 281967 167726
rect 429285 167723 429351 167726
rect 265249 167648 268210 167650
rect 265249 167592 265254 167648
rect 265310 167592 268210 167648
rect 265249 167590 268210 167592
rect 265249 167587 265315 167590
rect 265525 167242 265591 167245
rect 268150 167242 268210 167484
rect 265525 167240 268210 167242
rect 265525 167184 265530 167240
rect 265586 167184 268210 167240
rect 265525 167182 268210 167184
rect 265525 167179 265591 167182
rect 231209 167106 231275 167109
rect 228968 167104 231275 167106
rect 228968 167048 231214 167104
rect 231270 167048 231275 167104
rect 228968 167046 231275 167048
rect 231209 167043 231275 167046
rect 265157 167106 265223 167109
rect 282361 167106 282427 167109
rect 265157 167104 268026 167106
rect 265157 167048 265162 167104
rect 265218 167048 268026 167104
rect 279956 167104 282427 167106
rect 265157 167046 268026 167048
rect 265157 167043 265223 167046
rect 267966 167010 268026 167046
rect 268150 167010 268210 167076
rect 279956 167048 282366 167104
rect 282422 167048 282427 167104
rect 279956 167046 282427 167048
rect 282361 167043 282427 167046
rect 214097 166970 214163 166973
rect 216998 166970 217242 167010
rect 214097 166968 217242 166970
rect 214097 166912 214102 166968
rect 214158 166950 217242 166968
rect 267966 166950 268210 167010
rect 427862 166973 427922 167212
rect 427862 166968 427971 166973
rect 214158 166912 217058 166950
rect 217182 166940 217242 166950
rect 214097 166910 217058 166912
rect 427862 166912 427910 166968
rect 427966 166912 427971 166968
rect 427862 166910 427971 166912
rect 214097 166907 214163 166910
rect 427905 166907 427971 166910
rect 214649 166698 214715 166701
rect 231761 166698 231827 166701
rect 214649 166696 217242 166698
rect 214649 166640 214654 166696
rect 214710 166640 217242 166696
rect 214649 166638 217242 166640
rect 228968 166696 231827 166698
rect 228968 166640 231766 166696
rect 231822 166640 231827 166696
rect 228968 166638 231827 166640
rect 214649 166635 214715 166638
rect 217182 166396 217242 166638
rect 231761 166635 231827 166638
rect 265617 166426 265683 166429
rect 268150 166426 268210 166668
rect 265617 166424 268210 166426
rect 265617 166368 265622 166424
rect 265678 166368 268210 166424
rect 265617 166366 268210 166368
rect 265617 166363 265683 166366
rect 282085 166290 282151 166293
rect 279956 166288 282151 166290
rect 213913 166154 213979 166157
rect 231485 166154 231551 166157
rect 213913 166152 217242 166154
rect 213913 166096 213918 166152
rect 213974 166096 217242 166152
rect 213913 166094 217242 166096
rect 228968 166152 231551 166154
rect 228968 166096 231490 166152
rect 231546 166096 231551 166152
rect 228968 166094 231551 166096
rect 213913 166091 213979 166094
rect 217182 165716 217242 166094
rect 231485 166091 231551 166094
rect 265893 166018 265959 166021
rect 268150 166018 268210 166260
rect 279956 166232 282090 166288
rect 282146 166232 282151 166288
rect 279956 166230 282151 166232
rect 282085 166227 282151 166230
rect 346853 166290 346919 166293
rect 346853 166288 350060 166290
rect 346853 166232 346858 166288
rect 346914 166232 350060 166288
rect 346853 166230 350060 166232
rect 346853 166227 346919 166230
rect 429101 166154 429167 166157
rect 265893 166016 268210 166018
rect 265893 165960 265898 166016
rect 265954 165960 268210 166016
rect 265893 165958 268210 165960
rect 428230 166152 429167 166154
rect 428230 166096 429106 166152
rect 429162 166096 429167 166152
rect 428230 166094 429167 166096
rect 265893 165955 265959 165958
rect 231577 165746 231643 165749
rect 228968 165744 231643 165746
rect 228968 165688 231582 165744
rect 231638 165688 231643 165744
rect 228968 165686 231643 165688
rect 231577 165683 231643 165686
rect 265801 165746 265867 165749
rect 265801 165744 267842 165746
rect 265801 165688 265806 165744
rect 265862 165688 267842 165744
rect 265801 165686 267842 165688
rect 265801 165683 265867 165686
rect 267782 165610 267842 165686
rect 268334 165610 268394 165852
rect 427997 165746 428063 165749
rect 428230 165746 428290 166094
rect 429101 166091 429167 166094
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 427997 165744 428290 165746
rect 427997 165688 428002 165744
rect 428058 165688 428290 165744
rect 583520 165732 584960 165822
rect 427997 165686 428290 165688
rect 427997 165683 428063 165686
rect 267782 165550 268394 165610
rect 282361 165474 282427 165477
rect 279956 165472 282427 165474
rect 279956 165416 282366 165472
rect 282422 165416 282427 165472
rect 279956 165414 282427 165416
rect 282361 165411 282427 165414
rect 213913 165338 213979 165341
rect 213913 165336 217242 165338
rect 213913 165280 213918 165336
rect 213974 165280 217242 165336
rect 213913 165278 217242 165280
rect 213913 165275 213979 165278
rect 217182 165036 217242 165278
rect 231025 165202 231091 165205
rect 228968 165200 231091 165202
rect 228968 165144 231030 165200
rect 231086 165144 231091 165200
rect 228968 165142 231091 165144
rect 231025 165139 231091 165142
rect 264237 165066 264303 165069
rect 268150 165066 268210 165308
rect 430665 165066 430731 165069
rect 435030 165066 435036 165068
rect 264237 165064 268210 165066
rect 264237 165008 264242 165064
rect 264298 165008 268210 165064
rect 264237 165006 268210 165008
rect 428230 165064 435036 165066
rect 428230 165008 430670 165064
rect 430726 165008 435036 165064
rect 428230 165006 435036 165008
rect 264237 165003 264303 165006
rect 263041 164930 263107 164933
rect 263041 164928 268026 164930
rect 263041 164872 263046 164928
rect 263102 164896 268026 164928
rect 428230 164900 428290 165006
rect 430665 165003 430731 165006
rect 435030 165004 435036 165006
rect 435100 165004 435106 165068
rect 268150 164896 268210 164900
rect 263102 164872 268210 164896
rect 263041 164870 268210 164872
rect 263041 164867 263107 164870
rect 267966 164836 268210 164870
rect 214005 164794 214071 164797
rect 237414 164794 237420 164796
rect 214005 164792 217242 164794
rect 214005 164736 214010 164792
rect 214066 164736 217242 164792
rect 214005 164734 217242 164736
rect 228968 164734 237420 164794
rect 214005 164731 214071 164734
rect 217182 164356 217242 164734
rect 237414 164732 237420 164734
rect 237484 164732 237490 164796
rect 282085 164794 282151 164797
rect 279956 164792 282151 164794
rect 279956 164736 282090 164792
rect 282146 164736 282151 164792
rect 279956 164734 282151 164736
rect 282085 164731 282151 164734
rect 258030 164598 268210 164658
rect 239254 164460 239260 164524
rect 239324 164522 239330 164524
rect 258030 164522 258090 164598
rect 239324 164462 258090 164522
rect 268150 164492 268210 164598
rect 347497 164522 347563 164525
rect 347497 164520 350060 164522
rect 347497 164464 347502 164520
rect 347558 164464 350060 164520
rect 347497 164462 350060 164464
rect 239324 164460 239330 164462
rect 347497 164459 347563 164462
rect 231117 164386 231183 164389
rect 228968 164384 231183 164386
rect 228968 164328 231122 164384
rect 231178 164328 231183 164384
rect 228968 164326 231183 164328
rect 231117 164323 231183 164326
rect 213913 164114 213979 164117
rect 213913 164112 217242 164114
rect 213913 164056 213918 164112
rect 213974 164056 217242 164112
rect 213913 164054 217242 164056
rect 213913 164051 213979 164054
rect 217182 163676 217242 164054
rect 231761 163842 231827 163845
rect 228968 163840 231827 163842
rect 228968 163784 231766 163840
rect 231822 163784 231827 163840
rect 228968 163782 231827 163784
rect 231761 163779 231827 163782
rect 265985 163842 266051 163845
rect 268150 163842 268210 164084
rect 282821 163978 282887 163981
rect 430573 163978 430639 163981
rect 279956 163976 282887 163978
rect 279956 163920 282826 163976
rect 282882 163920 282887 163976
rect 279956 163918 282887 163920
rect 282821 163915 282887 163918
rect 428230 163976 430639 163978
rect 428230 163920 430578 163976
rect 430634 163920 430639 163976
rect 428230 163918 430639 163920
rect 265985 163840 268210 163842
rect 265985 163784 265990 163840
rect 266046 163784 268210 163840
rect 428230 163812 428290 163918
rect 430573 163915 430639 163918
rect 265985 163782 268210 163784
rect 265985 163779 266051 163782
rect 214005 163434 214071 163437
rect 231669 163434 231735 163437
rect 214005 163432 217242 163434
rect 214005 163376 214010 163432
rect 214066 163376 217242 163432
rect 214005 163374 217242 163376
rect 228968 163432 231735 163434
rect 228968 163376 231674 163432
rect 231730 163376 231735 163432
rect 228968 163374 231735 163376
rect 214005 163371 214071 163374
rect 217182 162996 217242 163374
rect 231669 163371 231735 163374
rect 265617 163434 265683 163437
rect 268150 163434 268210 163676
rect 265617 163432 268210 163434
rect 265617 163376 265622 163432
rect 265678 163376 268210 163432
rect 265617 163374 268210 163376
rect 265617 163371 265683 163374
rect 265525 163026 265591 163029
rect 268150 163026 268210 163268
rect 282177 163162 282243 163165
rect 279956 163160 282243 163162
rect 279956 163104 282182 163160
rect 282238 163104 282243 163160
rect 279956 163102 282243 163104
rect 282177 163099 282243 163102
rect 265525 163024 268210 163026
rect -960 162890 480 162980
rect 265525 162968 265530 163024
rect 265586 162968 268210 163024
rect 265525 162966 268210 162968
rect 265525 162963 265591 162966
rect 3417 162890 3483 162893
rect 231485 162890 231551 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect 228968 162888 231551 162890
rect 228968 162832 231490 162888
rect 231546 162832 231551 162888
rect 228968 162830 231551 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 231485 162827 231551 162830
rect 265433 162890 265499 162893
rect 346669 162890 346735 162893
rect 265433 162888 267842 162890
rect 265433 162832 265438 162888
rect 265494 162832 267842 162888
rect 346669 162888 350060 162890
rect 265433 162830 267842 162832
rect 265433 162827 265499 162830
rect 214557 162754 214623 162757
rect 214557 162752 217242 162754
rect 214557 162696 214562 162752
rect 214618 162696 217242 162752
rect 214557 162694 217242 162696
rect 214557 162691 214623 162694
rect 217182 162316 217242 162694
rect 267782 162618 267842 162830
rect 268334 162618 268394 162860
rect 346669 162832 346674 162888
rect 346730 162832 350060 162888
rect 346669 162830 350060 162832
rect 346669 162827 346735 162830
rect 267782 162558 268394 162618
rect 231945 162482 232011 162485
rect 282085 162482 282151 162485
rect 228968 162480 232011 162482
rect 228968 162424 231950 162480
rect 232006 162424 232011 162480
rect 228968 162422 232011 162424
rect 279956 162480 282151 162482
rect 279956 162424 282090 162480
rect 282146 162424 282151 162480
rect 279956 162422 282151 162424
rect 428046 162482 428106 162724
rect 430573 162482 430639 162485
rect 428046 162480 430639 162482
rect 428046 162424 430578 162480
rect 430634 162424 430639 162480
rect 428046 162422 430639 162424
rect 231945 162419 232011 162422
rect 282085 162419 282151 162422
rect 430573 162419 430639 162422
rect 213913 162074 213979 162077
rect 265709 162074 265775 162077
rect 268150 162074 268210 162316
rect 213913 162072 217242 162074
rect 213913 162016 213918 162072
rect 213974 162016 217242 162072
rect 213913 162014 217242 162016
rect 213913 162011 213979 162014
rect 217182 161772 217242 162014
rect 265709 162072 268210 162074
rect 265709 162016 265714 162072
rect 265770 162016 268210 162072
rect 265709 162014 268210 162016
rect 265709 162011 265775 162014
rect 231761 161938 231827 161941
rect 430573 161938 430639 161941
rect 228968 161936 231827 161938
rect 228968 161880 231766 161936
rect 231822 161880 231827 161936
rect 428230 161936 430639 161938
rect 228968 161878 231827 161880
rect 231761 161875 231827 161878
rect 265801 161666 265867 161669
rect 268518 161668 268578 161908
rect 428230 161880 430578 161936
rect 430634 161880 430639 161936
rect 428230 161878 430639 161880
rect 265801 161664 268210 161666
rect 265801 161608 265806 161664
rect 265862 161608 268210 161664
rect 265801 161606 268210 161608
rect 265801 161603 265867 161606
rect 229185 161530 229251 161533
rect 228968 161528 229251 161530
rect 228968 161472 229190 161528
rect 229246 161472 229251 161528
rect 268150 161500 268210 161606
rect 268510 161604 268516 161668
rect 268580 161604 268586 161668
rect 282821 161666 282887 161669
rect 279956 161664 282887 161666
rect 279956 161608 282826 161664
rect 282882 161608 282887 161664
rect 279956 161606 282887 161608
rect 282821 161603 282887 161606
rect 428230 161500 428290 161878
rect 430573 161875 430639 161878
rect 228968 161470 229251 161472
rect 229185 161467 229251 161470
rect 214741 161258 214807 161261
rect 264513 161258 264579 161261
rect 268510 161258 268516 161260
rect 214741 161256 217242 161258
rect 214741 161200 214746 161256
rect 214802 161200 217242 161256
rect 214741 161198 217242 161200
rect 214741 161195 214807 161198
rect 217182 161092 217242 161198
rect 264513 161256 268516 161258
rect 264513 161200 264518 161256
rect 264574 161200 268516 161256
rect 264513 161198 268516 161200
rect 264513 161195 264579 161198
rect 268510 161196 268516 161198
rect 268580 161196 268586 161260
rect 347497 161122 347563 161125
rect 347497 161120 350060 161122
rect 231301 160986 231367 160989
rect 228968 160984 231367 160986
rect 228968 160928 231306 160984
rect 231362 160928 231367 160984
rect 228968 160926 231367 160928
rect 231301 160923 231367 160926
rect 265341 160850 265407 160853
rect 268150 160850 268210 161092
rect 347497 161064 347502 161120
rect 347558 161064 350060 161120
rect 347497 161062 350060 161064
rect 347497 161059 347563 161062
rect 430573 160986 430639 160989
rect 428230 160984 430639 160986
rect 428230 160928 430578 160984
rect 430634 160928 430639 160984
rect 428230 160926 430639 160928
rect 282821 160850 282887 160853
rect 265341 160848 268210 160850
rect 265341 160792 265346 160848
rect 265402 160792 268210 160848
rect 265341 160790 268210 160792
rect 279956 160848 282887 160850
rect 279956 160792 282826 160848
rect 282882 160792 282887 160848
rect 279956 160790 282887 160792
rect 265341 160787 265407 160790
rect 282821 160787 282887 160790
rect 231761 160578 231827 160581
rect 228968 160576 231827 160578
rect 228968 160520 231766 160576
rect 231822 160520 231827 160576
rect 228968 160518 231827 160520
rect 231761 160515 231827 160518
rect 265617 160442 265683 160445
rect 268150 160442 268210 160684
rect 265617 160440 268210 160442
rect 166206 160108 166212 160172
rect 166276 160170 166282 160172
rect 217182 160170 217242 160412
rect 265617 160384 265622 160440
rect 265678 160384 268210 160440
rect 428230 160412 428290 160926
rect 430573 160923 430639 160926
rect 265617 160382 268210 160384
rect 265617 160379 265683 160382
rect 166276 160110 217242 160170
rect 265801 160170 265867 160173
rect 265801 160168 267842 160170
rect 265801 160112 265806 160168
rect 265862 160112 267842 160168
rect 265801 160110 267842 160112
rect 166276 160108 166282 160110
rect 265801 160107 265867 160110
rect 213913 160034 213979 160037
rect 231577 160034 231643 160037
rect 213913 160032 217242 160034
rect 213913 159976 213918 160032
rect 213974 159976 217242 160032
rect 213913 159974 217242 159976
rect 228968 160032 231643 160034
rect 228968 159976 231582 160032
rect 231638 159976 231643 160032
rect 228968 159974 231643 159976
rect 267782 160034 267842 160110
rect 268334 160034 268394 160276
rect 282729 160170 282795 160173
rect 279956 160168 282795 160170
rect 279956 160112 282734 160168
rect 282790 160112 282795 160168
rect 279956 160110 282795 160112
rect 282729 160107 282795 160110
rect 267782 159974 268394 160034
rect 213913 159971 213979 159974
rect 217182 159732 217242 159974
rect 231577 159971 231643 159974
rect 430573 159762 430639 159765
rect 428230 159760 430639 159762
rect 231025 159626 231091 159629
rect 228968 159624 231091 159626
rect 228968 159568 231030 159624
rect 231086 159568 231091 159624
rect 228968 159566 231091 159568
rect 231025 159563 231091 159566
rect 214005 159490 214071 159493
rect 265893 159490 265959 159493
rect 268150 159490 268210 159732
rect 428230 159704 430578 159760
rect 430634 159704 430639 159760
rect 428230 159702 430639 159704
rect 214005 159488 217242 159490
rect 214005 159432 214010 159488
rect 214066 159432 217242 159488
rect 214005 159430 217242 159432
rect 214005 159427 214071 159430
rect 217182 159052 217242 159430
rect 265893 159488 268210 159490
rect 265893 159432 265898 159488
rect 265954 159432 268210 159488
rect 265893 159430 268210 159432
rect 347497 159490 347563 159493
rect 347497 159488 350060 159490
rect 347497 159432 347502 159488
rect 347558 159432 350060 159488
rect 347497 159430 350060 159432
rect 265893 159427 265959 159430
rect 347497 159427 347563 159430
rect 282085 159354 282151 159357
rect 279956 159352 282151 159354
rect 231761 159082 231827 159085
rect 228968 159080 231827 159082
rect 228968 159024 231766 159080
rect 231822 159024 231827 159080
rect 228968 159022 231827 159024
rect 231761 159019 231827 159022
rect 265801 159082 265867 159085
rect 268150 159082 268210 159324
rect 279956 159296 282090 159352
rect 282146 159296 282151 159352
rect 428230 159324 428290 159702
rect 430573 159699 430639 159702
rect 279956 159294 282151 159296
rect 282085 159291 282151 159294
rect 265801 159080 268210 159082
rect 265801 159024 265806 159080
rect 265862 159024 268210 159080
rect 265801 159022 268210 159024
rect 265801 159019 265867 159022
rect 265709 158810 265775 158813
rect 265709 158808 267842 158810
rect 265709 158752 265714 158808
rect 265770 158752 267842 158808
rect 265709 158750 267842 158752
rect 265709 158747 265775 158750
rect 213913 158674 213979 158677
rect 230473 158674 230539 158677
rect 213913 158672 217242 158674
rect 213913 158616 213918 158672
rect 213974 158616 217242 158672
rect 213913 158614 217242 158616
rect 228968 158672 230539 158674
rect 228968 158616 230478 158672
rect 230534 158616 230539 158672
rect 228968 158614 230539 158616
rect 267782 158674 267842 158750
rect 268334 158674 268394 158916
rect 267782 158614 268394 158674
rect 213913 158611 213979 158614
rect 217182 158372 217242 158614
rect 230473 158611 230539 158614
rect 282821 158538 282887 158541
rect 430573 158538 430639 158541
rect 279956 158536 282887 158538
rect 265709 158266 265775 158269
rect 268150 158266 268210 158508
rect 279956 158480 282826 158536
rect 282882 158480 282887 158536
rect 279956 158478 282887 158480
rect 282821 158475 282887 158478
rect 428230 158536 430639 158538
rect 428230 158480 430578 158536
rect 430634 158480 430639 158536
rect 428230 158478 430639 158480
rect 265709 158264 268210 158266
rect 265709 158208 265714 158264
rect 265770 158208 268210 158264
rect 428230 158236 428290 158478
rect 430573 158475 430639 158478
rect 265709 158206 268210 158208
rect 265709 158203 265775 158206
rect 213361 158130 213427 158133
rect 231209 158130 231275 158133
rect 213361 158128 217242 158130
rect 213361 158072 213366 158128
rect 213422 158072 217242 158128
rect 213361 158070 217242 158072
rect 228968 158128 231275 158130
rect 228968 158072 231214 158128
rect 231270 158072 231275 158128
rect 228968 158070 231275 158072
rect 213361 158067 213427 158070
rect 168230 157932 168236 157996
rect 168300 157994 168306 157996
rect 214005 157994 214071 157997
rect 168300 157992 214071 157994
rect 168300 157936 214010 157992
rect 214066 157936 214071 157992
rect 168300 157934 214071 157936
rect 168300 157932 168306 157934
rect 214005 157931 214071 157934
rect 217182 157692 217242 158070
rect 231209 158067 231275 158070
rect 265617 157858 265683 157861
rect 268150 157858 268210 158100
rect 282729 157858 282795 157861
rect 265617 157856 268210 157858
rect 265617 157800 265622 157856
rect 265678 157800 268210 157856
rect 265617 157798 268210 157800
rect 279956 157856 282795 157858
rect 279956 157800 282734 157856
rect 282790 157800 282795 157856
rect 279956 157798 282795 157800
rect 265617 157795 265683 157798
rect 282729 157795 282795 157798
rect 347497 157858 347563 157861
rect 347497 157856 350060 157858
rect 347497 157800 347502 157856
rect 347558 157800 350060 157856
rect 347497 157798 350060 157800
rect 347497 157795 347563 157798
rect 231761 157722 231827 157725
rect 228968 157720 231827 157722
rect 228968 157664 231766 157720
rect 231822 157664 231827 157720
rect 228968 157662 231827 157664
rect 231761 157659 231827 157662
rect 230105 157450 230171 157453
rect 237598 157450 237604 157452
rect 230105 157448 237604 157450
rect 230105 157392 230110 157448
rect 230166 157392 237604 157448
rect 230105 157390 237604 157392
rect 230105 157387 230171 157390
rect 237598 157388 237604 157390
rect 237668 157388 237674 157452
rect 265157 157450 265223 157453
rect 268334 157450 268394 157692
rect 265157 157448 268394 157450
rect 265157 157392 265162 157448
rect 265218 157392 268394 157448
rect 265157 157390 268394 157392
rect 265157 157387 265223 157390
rect 214005 157314 214071 157317
rect 214005 157312 217242 157314
rect 214005 157256 214010 157312
rect 214066 157256 217242 157312
rect 214005 157254 217242 157256
rect 214005 157251 214071 157254
rect 217182 157148 217242 157254
rect 231761 157178 231827 157181
rect 430573 157178 430639 157181
rect 228968 157176 231827 157178
rect 228968 157120 231766 157176
rect 231822 157120 231827 157176
rect 428230 157176 430639 157178
rect 228968 157118 231827 157120
rect 231761 157115 231827 157118
rect 213913 156906 213979 156909
rect 265525 156906 265591 156909
rect 268150 156906 268210 157148
rect 428230 157120 430578 157176
rect 430634 157120 430639 157176
rect 428230 157118 430639 157120
rect 282085 157042 282151 157045
rect 279956 157040 282151 157042
rect 279956 156984 282090 157040
rect 282146 156984 282151 157040
rect 428230 157012 428290 157118
rect 430573 157115 430639 157118
rect 279956 156982 282151 156984
rect 282085 156979 282151 156982
rect 213913 156904 217242 156906
rect 213913 156848 213918 156904
rect 213974 156848 217242 156904
rect 213913 156846 217242 156848
rect 213913 156843 213979 156846
rect 217182 156468 217242 156846
rect 265525 156904 268210 156906
rect 265525 156848 265530 156904
rect 265586 156848 268210 156904
rect 265525 156846 268210 156848
rect 265525 156843 265591 156846
rect 231117 156770 231183 156773
rect 228968 156768 231183 156770
rect 228968 156712 231122 156768
rect 231178 156712 231183 156768
rect 228968 156710 231183 156712
rect 231117 156707 231183 156710
rect 265893 156498 265959 156501
rect 268150 156498 268210 156740
rect 265893 156496 268210 156498
rect 265893 156440 265898 156496
rect 265954 156440 268210 156496
rect 265893 156438 268210 156440
rect 265893 156435 265959 156438
rect 280337 156362 280403 156365
rect 279956 156360 280403 156362
rect 230933 156226 230999 156229
rect 228968 156224 230999 156226
rect 228968 156168 230938 156224
rect 230994 156168 230999 156224
rect 228968 156166 230999 156168
rect 230933 156163 230999 156166
rect 265985 156090 266051 156093
rect 268150 156090 268210 156332
rect 279956 156304 280342 156360
rect 280398 156304 280403 156360
rect 279956 156302 280403 156304
rect 280337 156299 280403 156302
rect 265985 156088 268210 156090
rect 265985 156032 265990 156088
rect 266046 156032 268210 156088
rect 265985 156030 268210 156032
rect 347037 156090 347103 156093
rect 347037 156088 350060 156090
rect 347037 156032 347042 156088
rect 347098 156032 350060 156088
rect 347037 156030 350060 156032
rect 265985 156027 266051 156030
rect 347037 156027 347103 156030
rect 213913 155954 213979 155957
rect 213913 155952 217242 155954
rect 213913 155896 213918 155952
rect 213974 155896 217242 155952
rect 213913 155894 217242 155896
rect 213913 155891 213979 155894
rect 217182 155788 217242 155894
rect 232037 155818 232103 155821
rect 228968 155816 232103 155818
rect 228968 155760 232042 155816
rect 232098 155760 232103 155816
rect 228968 155758 232103 155760
rect 232037 155755 232103 155758
rect 265525 155682 265591 155685
rect 268150 155682 268210 155924
rect 265525 155680 268210 155682
rect 265525 155624 265530 155680
rect 265586 155624 268210 155680
rect 265525 155622 268210 155624
rect 428046 155682 428106 155924
rect 430573 155682 430639 155685
rect 428046 155680 430639 155682
rect 428046 155624 430578 155680
rect 430634 155624 430639 155680
rect 428046 155622 430639 155624
rect 265525 155619 265591 155622
rect 430573 155619 430639 155622
rect 214005 155546 214071 155549
rect 282085 155546 282151 155549
rect 214005 155544 217242 155546
rect 214005 155488 214010 155544
rect 214066 155488 217242 155544
rect 279956 155544 282151 155546
rect 214005 155486 217242 155488
rect 214005 155483 214071 155486
rect 217182 155108 217242 155486
rect 231761 155274 231827 155277
rect 228968 155272 231827 155274
rect 228968 155216 231766 155272
rect 231822 155216 231827 155272
rect 228968 155214 231827 155216
rect 231761 155211 231827 155214
rect 265801 155274 265867 155277
rect 268150 155274 268210 155516
rect 279956 155488 282090 155544
rect 282146 155488 282151 155544
rect 279956 155486 282151 155488
rect 282085 155483 282151 155486
rect 430849 155410 430915 155413
rect 265801 155272 268210 155274
rect 265801 155216 265806 155272
rect 265862 155216 268210 155272
rect 265801 155214 268210 155216
rect 428230 155408 430915 155410
rect 428230 155352 430854 155408
rect 430910 155352 430915 155408
rect 428230 155350 430915 155352
rect 265801 155211 265867 155214
rect 231485 154866 231551 154869
rect 228968 154864 231551 154866
rect 228968 154808 231490 154864
rect 231546 154808 231551 154864
rect 228968 154806 231551 154808
rect 231485 154803 231551 154806
rect 265985 154730 266051 154733
rect 268518 154730 268578 155108
rect 428230 154836 428290 155350
rect 430849 155347 430915 155350
rect 282361 154730 282427 154733
rect 265985 154728 268578 154730
rect 265985 154672 265990 154728
rect 266046 154672 268578 154728
rect 265985 154670 268578 154672
rect 279956 154728 282427 154730
rect 279956 154672 282366 154728
rect 282422 154672 282427 154728
rect 279956 154670 282427 154672
rect 265985 154667 266051 154670
rect 282361 154667 282427 154670
rect 231158 154532 231164 154596
rect 231228 154594 231234 154596
rect 237373 154594 237439 154597
rect 231228 154592 237439 154594
rect 231228 154536 237378 154592
rect 237434 154536 237439 154592
rect 231228 154534 237439 154536
rect 231228 154532 231234 154534
rect 237373 154531 237439 154534
rect 265709 154594 265775 154597
rect 265709 154592 267842 154594
rect 265709 154536 265714 154592
rect 265770 154536 267842 154592
rect 265709 154534 267842 154536
rect 265709 154531 265775 154534
rect 214005 153914 214071 153917
rect 217182 153914 217242 154428
rect 231761 154322 231827 154325
rect 228968 154320 231827 154322
rect 228968 154264 231766 154320
rect 231822 154264 231827 154320
rect 228968 154262 231827 154264
rect 267782 154322 267842 154534
rect 268334 154322 268394 154564
rect 346669 154458 346735 154461
rect 346669 154456 350060 154458
rect 346669 154400 346674 154456
rect 346730 154400 350060 154456
rect 346669 154398 350060 154400
rect 346669 154395 346735 154398
rect 267782 154262 268394 154322
rect 231761 154259 231827 154262
rect 430573 154186 430639 154189
rect 428230 154184 430639 154186
rect 231669 153914 231735 153917
rect 214005 153912 217242 153914
rect 214005 153856 214010 153912
rect 214066 153856 217242 153912
rect 214005 153854 217242 153856
rect 228968 153912 231735 153914
rect 228968 153856 231674 153912
rect 231730 153856 231735 153912
rect 228968 153854 231735 153856
rect 214005 153851 214071 153854
rect 231669 153851 231735 153854
rect 265893 153914 265959 153917
rect 268150 153914 268210 154156
rect 428230 154128 430578 154184
rect 430634 154128 430639 154184
rect 428230 154126 430639 154128
rect 281901 154050 281967 154053
rect 279956 154048 281967 154050
rect 279956 153992 281906 154048
rect 281962 153992 281967 154048
rect 279956 153990 281967 153992
rect 281901 153987 281967 153990
rect 265893 153912 268210 153914
rect 265893 153856 265898 153912
rect 265954 153856 268210 153912
rect 265893 153854 268210 153856
rect 265893 153851 265959 153854
rect 428230 153748 428290 154126
rect 430573 154123 430639 154126
rect 213913 153506 213979 153509
rect 217182 153506 217242 153748
rect 213913 153504 217242 153506
rect 213913 153448 213918 153504
rect 213974 153448 217242 153504
rect 213913 153446 217242 153448
rect 265801 153506 265867 153509
rect 268150 153506 268210 153748
rect 265801 153504 268210 153506
rect 265801 153448 265806 153504
rect 265862 153448 268210 153504
rect 265801 153446 268210 153448
rect 213913 153443 213979 153446
rect 265801 153443 265867 153446
rect 233182 153370 233188 153372
rect 228968 153310 233188 153370
rect 233182 153308 233188 153310
rect 233252 153308 233258 153372
rect 265801 153234 265867 153237
rect 265801 153232 267842 153234
rect 265801 153176 265806 153232
rect 265862 153176 267842 153232
rect 265801 153174 267842 153176
rect 265801 153171 265867 153174
rect 267782 153098 267842 153174
rect 268334 153098 268394 153340
rect 282453 153234 282519 153237
rect 279956 153232 282519 153234
rect 279956 153176 282458 153232
rect 282514 153176 282519 153232
rect 279956 153174 282519 153176
rect 282453 153171 282519 153174
rect 213913 152690 213979 152693
rect 217182 152690 217242 153068
rect 267782 153038 268394 153098
rect 231761 152962 231827 152965
rect 228968 152960 231827 152962
rect 228968 152904 231766 152960
rect 231822 152904 231827 152960
rect 228968 152902 231827 152904
rect 231761 152899 231827 152902
rect 213913 152688 217242 152690
rect 213913 152632 213918 152688
rect 213974 152632 217242 152688
rect 213913 152630 217242 152632
rect 266077 152690 266143 152693
rect 268150 152690 268210 152932
rect 430573 152826 430639 152829
rect 428230 152824 430639 152826
rect 428230 152768 430578 152824
rect 430634 152768 430639 152824
rect 428230 152766 430639 152768
rect 266077 152688 268210 152690
rect 266077 152632 266082 152688
rect 266138 152632 268210 152688
rect 266077 152630 268210 152632
rect 346577 152690 346643 152693
rect 346577 152688 350060 152690
rect 346577 152632 346582 152688
rect 346638 152632 350060 152688
rect 346577 152630 350060 152632
rect 213913 152627 213979 152630
rect 266077 152627 266143 152630
rect 346577 152627 346643 152630
rect 241646 152554 241652 152556
rect 214005 152282 214071 152285
rect 217182 152282 217242 152524
rect 228968 152494 241652 152554
rect 241646 152492 241652 152494
rect 241716 152492 241722 152556
rect 428230 152524 428290 152766
rect 430573 152763 430639 152766
rect 582373 152690 582439 152693
rect 583520 152690 584960 152780
rect 582373 152688 584960 152690
rect 582373 152632 582378 152688
rect 582434 152632 584960 152688
rect 582373 152630 584960 152632
rect 582373 152627 582439 152630
rect 583520 152540 584960 152630
rect 237966 152356 237972 152420
rect 238036 152418 238042 152420
rect 265801 152418 265867 152421
rect 238036 152416 265867 152418
rect 238036 152360 265806 152416
rect 265862 152360 265867 152416
rect 238036 152358 265867 152360
rect 238036 152356 238042 152358
rect 265801 152355 265867 152358
rect 214005 152280 217242 152282
rect 214005 152224 214010 152280
rect 214066 152224 217242 152280
rect 214005 152222 217242 152224
rect 214005 152219 214071 152222
rect 265985 152146 266051 152149
rect 268150 152146 268210 152524
rect 281533 152418 281599 152421
rect 279956 152416 281599 152418
rect 279956 152360 281538 152416
rect 281594 152360 281599 152416
rect 279956 152358 281599 152360
rect 281533 152355 281599 152358
rect 265985 152144 268210 152146
rect 265985 152088 265990 152144
rect 266046 152088 268210 152144
rect 265985 152086 268210 152088
rect 265985 152083 266051 152086
rect 213913 152010 213979 152013
rect 231577 152010 231643 152013
rect 213913 152008 217242 152010
rect 213913 151952 213918 152008
rect 213974 151952 217242 152008
rect 213913 151950 217242 151952
rect 228968 152008 231643 152010
rect 228968 151952 231582 152008
rect 231638 151952 231643 152008
rect 228968 151950 231643 151952
rect 213913 151947 213979 151950
rect 217182 151844 217242 151950
rect 231577 151947 231643 151950
rect 265801 151874 265867 151877
rect 265801 151872 267842 151874
rect 265801 151816 265806 151872
rect 265862 151816 267842 151872
rect 265801 151814 267842 151816
rect 265801 151811 265867 151814
rect 267782 151738 267842 151814
rect 268334 151738 268394 151980
rect 281901 151738 281967 151741
rect 267782 151678 268394 151738
rect 279956 151736 281967 151738
rect 279956 151680 281906 151736
rect 281962 151680 281967 151736
rect 279956 151678 281967 151680
rect 281901 151675 281967 151678
rect 231761 151602 231827 151605
rect 430573 151602 430639 151605
rect 228968 151600 231827 151602
rect 228968 151544 231766 151600
rect 231822 151544 231827 151600
rect 428230 151600 430639 151602
rect 228968 151542 231827 151544
rect 231761 151539 231827 151542
rect 265893 151330 265959 151333
rect 268150 151330 268210 151572
rect 428230 151544 430578 151600
rect 430634 151544 430639 151600
rect 428230 151542 430639 151544
rect 428230 151436 428290 151542
rect 430573 151539 430639 151542
rect 265893 151328 268210 151330
rect 265893 151272 265898 151328
rect 265954 151272 268210 151328
rect 265893 151270 268210 151272
rect 265893 151267 265959 151270
rect 214649 150786 214715 150789
rect 217182 150786 217242 151164
rect 231669 151058 231735 151061
rect 228968 151056 231735 151058
rect 228968 151000 231674 151056
rect 231730 151000 231735 151056
rect 228968 150998 231735 151000
rect 231669 150995 231735 150998
rect 265801 150922 265867 150925
rect 268150 150922 268210 151164
rect 346669 151058 346735 151061
rect 346669 151056 350060 151058
rect 346669 151000 346674 151056
rect 346730 151000 350060 151056
rect 346669 150998 350060 151000
rect 346669 150995 346735 150998
rect 282269 150922 282335 150925
rect 265801 150920 268210 150922
rect 265801 150864 265806 150920
rect 265862 150864 268210 150920
rect 265801 150862 268210 150864
rect 279956 150920 282335 150922
rect 279956 150864 282274 150920
rect 282330 150864 282335 150920
rect 279956 150862 282335 150864
rect 265801 150859 265867 150862
rect 282269 150859 282335 150862
rect 214649 150784 217242 150786
rect 214649 150728 214654 150784
rect 214710 150728 217242 150784
rect 214649 150726 217242 150728
rect 214649 150723 214715 150726
rect 214005 150650 214071 150653
rect 230473 150650 230539 150653
rect 214005 150648 217242 150650
rect 214005 150592 214010 150648
rect 214066 150592 217242 150648
rect 214005 150590 217242 150592
rect 228968 150648 230539 150650
rect 228968 150592 230478 150648
rect 230534 150592 230539 150648
rect 228968 150590 230539 150592
rect 214005 150587 214071 150590
rect 217182 150484 217242 150590
rect 230473 150587 230539 150590
rect 265750 150452 265756 150516
rect 265820 150514 265826 150516
rect 268150 150514 268210 150756
rect 265820 150454 268210 150514
rect 265820 150452 265826 150454
rect 213913 150106 213979 150109
rect 234654 150106 234660 150108
rect 213913 150104 217242 150106
rect 213913 150048 213918 150104
rect 213974 150048 217242 150104
rect 213913 150046 217242 150048
rect 228968 150046 234660 150106
rect 213913 150043 213979 150046
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect 217182 149804 217242 150046
rect 234654 150044 234660 150046
rect 234724 150044 234730 150108
rect 265893 150106 265959 150109
rect 268150 150106 268210 150348
rect 282821 150106 282887 150109
rect 265893 150104 268210 150106
rect 265893 150048 265898 150104
rect 265954 150048 268210 150104
rect 265893 150046 268210 150048
rect 279956 150104 282887 150106
rect 279956 150048 282826 150104
rect 282882 150048 282887 150104
rect 279956 150046 282887 150048
rect 428046 150106 428106 150348
rect 430573 150106 430639 150109
rect 428046 150104 430639 150106
rect 428046 150048 430578 150104
rect 430634 150048 430639 150104
rect 428046 150046 430639 150048
rect 265893 150043 265959 150046
rect 282821 150043 282887 150046
rect 430573 150043 430639 150046
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 231761 149698 231827 149701
rect 228968 149696 231827 149698
rect 228968 149640 231766 149696
rect 231822 149640 231827 149696
rect 228968 149638 231827 149640
rect 231761 149635 231827 149638
rect 265249 149698 265315 149701
rect 268150 149698 268210 149940
rect 430849 149834 430915 149837
rect 265249 149696 268210 149698
rect 265249 149640 265254 149696
rect 265310 149640 268210 149696
rect 265249 149638 268210 149640
rect 428230 149832 430915 149834
rect 428230 149776 430854 149832
rect 430910 149776 430915 149832
rect 428230 149774 430915 149776
rect 265249 149635 265315 149638
rect 214557 149562 214623 149565
rect 214557 149560 217242 149562
rect 214557 149504 214562 149560
rect 214618 149504 217242 149560
rect 214557 149502 217242 149504
rect 214557 149499 214623 149502
rect 217182 149124 217242 149502
rect 231669 149154 231735 149157
rect 228968 149152 231735 149154
rect 228968 149096 231674 149152
rect 231730 149096 231735 149152
rect 228968 149094 231735 149096
rect 231669 149091 231735 149094
rect 265801 149154 265867 149157
rect 268150 149154 268210 149532
rect 282729 149426 282795 149429
rect 279956 149424 282795 149426
rect 279956 149368 282734 149424
rect 282790 149368 282795 149424
rect 279956 149366 282795 149368
rect 282729 149363 282795 149366
rect 347497 149290 347563 149293
rect 347497 149288 350060 149290
rect 347497 149232 347502 149288
rect 347558 149232 350060 149288
rect 428230 149260 428290 149774
rect 430849 149771 430915 149774
rect 347497 149230 350060 149232
rect 347497 149227 347563 149230
rect 265801 149152 268210 149154
rect 265801 149096 265806 149152
rect 265862 149096 268210 149152
rect 265801 149094 268210 149096
rect 265801 149091 265867 149094
rect 213913 148746 213979 148749
rect 233366 148746 233372 148748
rect 213913 148744 217242 148746
rect 213913 148688 213918 148744
rect 213974 148688 217242 148744
rect 213913 148686 217242 148688
rect 228968 148686 233372 148746
rect 213913 148683 213979 148686
rect 217182 148444 217242 148686
rect 233366 148684 233372 148686
rect 233436 148684 233442 148748
rect 265709 148746 265775 148749
rect 268150 148746 268210 148988
rect 265709 148744 268210 148746
rect 265709 148688 265714 148744
rect 265770 148688 268210 148744
rect 265709 148686 268210 148688
rect 265709 148683 265775 148686
rect 282821 148610 282887 148613
rect 430573 148610 430639 148613
rect 279956 148608 282887 148610
rect 265433 148338 265499 148341
rect 268150 148338 268210 148580
rect 279956 148552 282826 148608
rect 282882 148552 282887 148608
rect 279956 148550 282887 148552
rect 282821 148547 282887 148550
rect 428230 148608 430639 148610
rect 428230 148552 430578 148608
rect 430634 148552 430639 148608
rect 428230 148550 430639 148552
rect 265433 148336 268210 148338
rect 265433 148280 265438 148336
rect 265494 148280 268210 148336
rect 265433 148278 268210 148280
rect 265433 148275 265499 148278
rect 231301 148202 231367 148205
rect 228968 148200 231367 148202
rect 228968 148144 231306 148200
rect 231362 148144 231367 148200
rect 428230 148172 428290 148550
rect 430573 148547 430639 148550
rect 228968 148142 231367 148144
rect 231301 148139 231367 148142
rect 213913 148066 213979 148069
rect 213913 148064 217242 148066
rect 213913 148008 213918 148064
rect 213974 148008 217242 148064
rect 213913 148006 217242 148008
rect 213913 148003 213979 148006
rect 217182 147900 217242 148006
rect 265065 147930 265131 147933
rect 268518 147932 268578 148172
rect 265065 147928 268210 147930
rect 265065 147872 265070 147928
rect 265126 147872 268210 147928
rect 265065 147870 268210 147872
rect 265065 147867 265131 147870
rect 230749 147794 230815 147797
rect 228968 147792 230815 147794
rect 228968 147736 230754 147792
rect 230810 147736 230815 147792
rect 268150 147764 268210 147870
rect 268510 147868 268516 147932
rect 268580 147868 268586 147932
rect 280245 147794 280311 147797
rect 279956 147792 280311 147794
rect 228968 147734 230815 147736
rect 279956 147736 280250 147792
rect 280306 147736 280311 147792
rect 279956 147734 280311 147736
rect 230749 147731 230815 147734
rect 280245 147731 280311 147734
rect 346669 147658 346735 147661
rect 346669 147656 350060 147658
rect 346669 147600 346674 147656
rect 346730 147600 350060 147656
rect 346669 147598 350060 147600
rect 346669 147595 346735 147598
rect 432137 147522 432203 147525
rect 428230 147520 432203 147522
rect 428230 147464 432142 147520
rect 432198 147464 432203 147520
rect 428230 147462 432203 147464
rect 244222 147250 244228 147252
rect 213913 146706 213979 146709
rect 217182 146706 217242 147220
rect 228968 147190 244228 147250
rect 244222 147188 244228 147190
rect 244292 147188 244298 147252
rect 265709 147114 265775 147117
rect 268150 147114 268210 147356
rect 282821 147114 282887 147117
rect 265709 147112 268210 147114
rect 265709 147056 265714 147112
rect 265770 147056 268210 147112
rect 265709 147054 268210 147056
rect 279956 147112 282887 147114
rect 279956 147056 282826 147112
rect 282882 147056 282887 147112
rect 279956 147054 282887 147056
rect 265709 147051 265775 147054
rect 282821 147051 282887 147054
rect 233734 146916 233740 146980
rect 233804 146978 233810 146980
rect 265065 146978 265131 146981
rect 233804 146976 265131 146978
rect 233804 146920 265070 146976
rect 265126 146920 265131 146976
rect 428230 146948 428290 147462
rect 432137 147459 432203 147462
rect 233804 146918 265131 146920
rect 233804 146916 233810 146918
rect 265065 146915 265131 146918
rect 229277 146842 229343 146845
rect 228968 146840 229343 146842
rect 228968 146784 229282 146840
rect 229338 146784 229343 146840
rect 228968 146782 229343 146784
rect 229277 146779 229343 146782
rect 213913 146704 217242 146706
rect 213913 146648 213918 146704
rect 213974 146648 217242 146704
rect 213913 146646 217242 146648
rect 266169 146706 266235 146709
rect 268150 146706 268210 146948
rect 266169 146704 268210 146706
rect 266169 146648 266174 146704
rect 266230 146648 268210 146704
rect 266169 146646 268210 146648
rect 213913 146643 213979 146646
rect 266169 146643 266235 146646
rect 265433 146570 265499 146573
rect 265433 146568 268210 146570
rect 214097 146434 214163 146437
rect 214097 146432 216874 146434
rect 214097 146376 214102 146432
rect 214158 146376 216874 146432
rect 214097 146374 216874 146376
rect 214097 146371 214163 146374
rect 216814 146298 216874 146374
rect 217366 146298 217426 146540
rect 265433 146512 265438 146568
rect 265494 146512 268210 146568
rect 265433 146510 268210 146512
rect 265433 146507 265499 146510
rect 260373 146434 260439 146437
rect 265750 146434 265756 146436
rect 260373 146432 265756 146434
rect 260373 146376 260378 146432
rect 260434 146376 265756 146432
rect 260373 146374 265756 146376
rect 260373 146371 260439 146374
rect 265750 146372 265756 146374
rect 265820 146372 265826 146436
rect 268150 146404 268210 146510
rect 231761 146298 231827 146301
rect 282821 146298 282887 146301
rect 216814 146238 217426 146298
rect 228968 146296 231827 146298
rect 228968 146240 231766 146296
rect 231822 146240 231827 146296
rect 228968 146238 231827 146240
rect 279956 146296 282887 146298
rect 279956 146240 282826 146296
rect 282882 146240 282887 146296
rect 279956 146238 282887 146240
rect 231761 146235 231827 146238
rect 282821 146235 282887 146238
rect 261845 146162 261911 146165
rect 268510 146162 268516 146164
rect 261845 146160 268516 146162
rect 261845 146104 261850 146160
rect 261906 146104 268516 146160
rect 261845 146102 268516 146104
rect 261845 146099 261911 146102
rect 268510 146100 268516 146102
rect 268580 146100 268586 146164
rect 430573 146026 430639 146029
rect 428230 146024 430639 146026
rect 230841 145890 230907 145893
rect 228968 145888 230907 145890
rect 214005 145346 214071 145349
rect 217182 145346 217242 145860
rect 228968 145832 230846 145888
rect 230902 145832 230907 145888
rect 228968 145830 230907 145832
rect 230841 145827 230907 145830
rect 265893 145754 265959 145757
rect 268150 145754 268210 145996
rect 428230 145968 430578 146024
rect 430634 145968 430639 146024
rect 428230 145966 430639 145968
rect 346301 145890 346367 145893
rect 346485 145890 346551 145893
rect 346301 145888 350060 145890
rect 346301 145832 346306 145888
rect 346362 145832 346490 145888
rect 346546 145832 350060 145888
rect 428230 145860 428290 145966
rect 430573 145963 430639 145966
rect 346301 145830 350060 145832
rect 346301 145827 346367 145830
rect 346485 145827 346551 145830
rect 265893 145752 268210 145754
rect 265893 145696 265898 145752
rect 265954 145696 268210 145752
rect 265893 145694 268210 145696
rect 265893 145691 265959 145694
rect 231393 145346 231459 145349
rect 214005 145344 217242 145346
rect 214005 145288 214010 145344
rect 214066 145288 217242 145344
rect 214005 145286 217242 145288
rect 228968 145344 231459 145346
rect 228968 145288 231398 145344
rect 231454 145288 231459 145344
rect 228968 145286 231459 145288
rect 214005 145283 214071 145286
rect 231393 145283 231459 145286
rect 264329 145346 264395 145349
rect 268150 145346 268210 145588
rect 282729 145482 282795 145485
rect 279956 145480 282795 145482
rect 279956 145424 282734 145480
rect 282790 145424 282795 145480
rect 279956 145422 282795 145424
rect 282729 145419 282795 145422
rect 264329 145344 268210 145346
rect 264329 145288 264334 145344
rect 264390 145288 268210 145344
rect 264329 145286 268210 145288
rect 264329 145283 264395 145286
rect 213913 144938 213979 144941
rect 217366 144938 217426 145180
rect 245878 144938 245884 144940
rect 213913 144936 217426 144938
rect 213913 144880 213918 144936
rect 213974 144880 217426 144936
rect 213913 144878 217426 144880
rect 228968 144878 245884 144938
rect 213913 144875 213979 144878
rect 245878 144876 245884 144878
rect 245948 144876 245954 144940
rect 265801 144938 265867 144941
rect 268334 144938 268394 145180
rect 265801 144936 268394 144938
rect 265801 144880 265806 144936
rect 265862 144880 268394 144936
rect 265801 144878 268394 144880
rect 265801 144875 265867 144878
rect 282821 144802 282887 144805
rect 279956 144800 282887 144802
rect 265525 144530 265591 144533
rect 268150 144530 268210 144772
rect 279956 144744 282826 144800
rect 282882 144744 282887 144800
rect 279956 144742 282887 144744
rect 282821 144739 282887 144742
rect 265525 144528 268210 144530
rect 213913 143986 213979 143989
rect 217182 143986 217242 144500
rect 265525 144472 265530 144528
rect 265586 144472 268210 144528
rect 265525 144470 268210 144472
rect 428046 144530 428106 144772
rect 430573 144530 430639 144533
rect 428046 144528 430639 144530
rect 428046 144472 430578 144528
rect 430634 144472 430639 144528
rect 428046 144470 430639 144472
rect 265525 144467 265591 144470
rect 430573 144467 430639 144470
rect 231761 144394 231827 144397
rect 228968 144392 231827 144394
rect 228968 144336 231766 144392
rect 231822 144336 231827 144392
rect 228968 144334 231827 144336
rect 231761 144331 231827 144334
rect 231761 143986 231827 143989
rect 213913 143984 217242 143986
rect 213913 143928 213918 143984
rect 213974 143928 217242 143984
rect 213913 143926 217242 143928
rect 228968 143984 231827 143986
rect 228968 143928 231766 143984
rect 231822 143928 231827 143984
rect 228968 143926 231827 143928
rect 213913 143923 213979 143926
rect 231761 143923 231827 143926
rect 265709 143986 265775 143989
rect 268150 143986 268210 144364
rect 346669 144258 346735 144261
rect 346669 144256 350060 144258
rect 346669 144200 346674 144256
rect 346730 144200 350060 144256
rect 346669 144198 350060 144200
rect 346669 144195 346735 144198
rect 430849 144122 430915 144125
rect 428230 144120 430915 144122
rect 428230 144064 430854 144120
rect 430910 144064 430915 144120
rect 428230 144062 430915 144064
rect 282729 143986 282795 143989
rect 265709 143984 268210 143986
rect 265709 143928 265714 143984
rect 265770 143928 268210 143984
rect 265709 143926 268210 143928
rect 279956 143984 282795 143986
rect 279956 143928 282734 143984
rect 282790 143928 282795 143984
rect 279956 143926 282795 143928
rect 265709 143923 265775 143926
rect 282729 143923 282795 143926
rect 214005 143578 214071 143581
rect 217366 143578 217426 143820
rect 214005 143576 217426 143578
rect 214005 143520 214010 143576
rect 214066 143520 217426 143576
rect 214005 143518 217426 143520
rect 265801 143578 265867 143581
rect 268334 143578 268394 143820
rect 428230 143684 428290 144062
rect 430849 144059 430915 144062
rect 265801 143576 268394 143578
rect 265801 143520 265806 143576
rect 265862 143520 268394 143576
rect 265801 143518 268394 143520
rect 214005 143515 214071 143518
rect 265801 143515 265867 143518
rect 229921 143442 229987 143445
rect 228968 143440 229987 143442
rect 228968 143384 229926 143440
rect 229982 143384 229987 143440
rect 228968 143382 229987 143384
rect 229921 143379 229987 143382
rect 213269 142762 213335 142765
rect 217182 142762 217242 143276
rect 266077 143170 266143 143173
rect 268150 143170 268210 143412
rect 282085 143170 282151 143173
rect 266077 143168 268210 143170
rect 266077 143112 266082 143168
rect 266138 143112 268210 143168
rect 266077 143110 268210 143112
rect 279956 143168 282151 143170
rect 279956 143112 282090 143168
rect 282146 143112 282151 143168
rect 279956 143110 282151 143112
rect 266077 143107 266143 143110
rect 282085 143107 282151 143110
rect 231761 143034 231827 143037
rect 228968 143032 231827 143034
rect 228968 142976 231766 143032
rect 231822 142976 231827 143032
rect 228968 142974 231827 142976
rect 231761 142971 231827 142974
rect 213269 142760 217242 142762
rect 213269 142704 213274 142760
rect 213330 142704 217242 142760
rect 213269 142702 217242 142704
rect 213269 142699 213335 142702
rect 230974 142700 230980 142764
rect 231044 142762 231050 142764
rect 253105 142762 253171 142765
rect 231044 142760 253171 142762
rect 231044 142704 253110 142760
rect 253166 142704 253171 142760
rect 231044 142702 253171 142704
rect 231044 142700 231050 142702
rect 253105 142699 253171 142702
rect 265525 142762 265591 142765
rect 268150 142762 268210 143004
rect 265525 142760 268210 142762
rect 265525 142704 265530 142760
rect 265586 142704 268210 142760
rect 265525 142702 268210 142704
rect 265525 142699 265591 142702
rect 346577 142626 346643 142629
rect 346577 142624 350060 142626
rect 213913 142218 213979 142221
rect 217182 142218 217242 142596
rect 229737 142490 229803 142493
rect 228968 142488 229803 142490
rect 228968 142432 229742 142488
rect 229798 142432 229803 142488
rect 228968 142430 229803 142432
rect 229737 142427 229803 142430
rect 265617 142354 265683 142357
rect 268150 142354 268210 142596
rect 346577 142568 346582 142624
rect 346638 142568 350060 142624
rect 346577 142566 350060 142568
rect 346577 142563 346643 142566
rect 282821 142490 282887 142493
rect 279956 142488 282887 142490
rect 279956 142432 282826 142488
rect 282882 142432 282887 142488
rect 279956 142430 282887 142432
rect 282821 142427 282887 142430
rect 265617 142352 268210 142354
rect 265617 142296 265622 142352
rect 265678 142296 268210 142352
rect 265617 142294 268210 142296
rect 265617 142291 265683 142294
rect 213913 142216 217242 142218
rect 213913 142160 213918 142216
rect 213974 142160 217242 142216
rect 213913 142158 217242 142160
rect 265709 142218 265775 142221
rect 428046 142218 428106 142460
rect 430573 142218 430639 142221
rect 265709 142216 267842 142218
rect 265709 142160 265714 142216
rect 265770 142160 267842 142216
rect 428046 142216 430639 142218
rect 265709 142158 267842 142160
rect 213913 142155 213979 142158
rect 265709 142155 265775 142158
rect 236494 142082 236500 142084
rect 228968 142022 236500 142082
rect 236494 142020 236500 142022
rect 236564 142020 236570 142084
rect 267782 141946 267842 142158
rect 268334 141946 268394 142188
rect 428046 142160 430578 142216
rect 430634 142160 430639 142216
rect 428046 142158 430639 142160
rect 430573 142155 430639 142158
rect 214005 141402 214071 141405
rect 217182 141402 217242 141916
rect 267782 141886 268394 141946
rect 268510 141884 268516 141948
rect 268580 141884 268586 141948
rect 268518 141780 268578 141884
rect 231761 141674 231827 141677
rect 282821 141674 282887 141677
rect 228968 141672 231827 141674
rect 228968 141616 231766 141672
rect 231822 141616 231827 141672
rect 228968 141614 231827 141616
rect 279956 141672 282887 141674
rect 279956 141616 282826 141672
rect 282882 141616 282887 141672
rect 279956 141614 282887 141616
rect 231761 141611 231827 141614
rect 282821 141611 282887 141614
rect 264421 141538 264487 141541
rect 264421 141536 268578 141538
rect 264421 141480 264426 141536
rect 264482 141480 268578 141536
rect 264421 141478 268578 141480
rect 264421 141475 264487 141478
rect 214005 141400 217242 141402
rect 214005 141344 214010 141400
rect 214066 141344 217242 141400
rect 214005 141342 217242 141344
rect 214005 141339 214071 141342
rect 268518 141236 268578 141478
rect 213913 140994 213979 140997
rect 217182 140994 217242 141236
rect 231485 141130 231551 141133
rect 228968 141128 231551 141130
rect 228968 141072 231490 141128
rect 231546 141072 231551 141128
rect 228968 141070 231551 141072
rect 231485 141067 231551 141070
rect 213913 140992 217242 140994
rect 213913 140936 213918 140992
rect 213974 140936 217242 140992
rect 213913 140934 217242 140936
rect 265801 140994 265867 140997
rect 265801 140992 268210 140994
rect 265801 140936 265806 140992
rect 265862 140936 268210 140992
rect 265801 140934 268210 140936
rect 213913 140931 213979 140934
rect 265801 140931 265867 140934
rect 268150 140828 268210 140934
rect 282729 140858 282795 140861
rect 279956 140856 282795 140858
rect 279956 140800 282734 140856
rect 282790 140800 282795 140856
rect 279956 140798 282795 140800
rect 282729 140795 282795 140798
rect 346485 140858 346551 140861
rect 428230 140858 428290 141372
rect 429377 140858 429443 140861
rect 346485 140856 350060 140858
rect 346485 140800 346490 140856
rect 346546 140800 350060 140856
rect 346485 140798 350060 140800
rect 428230 140856 429443 140858
rect 428230 140800 429382 140856
rect 429438 140800 429443 140856
rect 428230 140798 429443 140800
rect 346485 140795 346551 140798
rect 429377 140795 429443 140798
rect 230657 140722 230723 140725
rect 228968 140720 230723 140722
rect 228968 140664 230662 140720
rect 230718 140664 230723 140720
rect 228968 140662 230723 140664
rect 230657 140659 230723 140662
rect 264605 140586 264671 140589
rect 268510 140586 268516 140588
rect 264605 140584 268516 140586
rect 213913 140042 213979 140045
rect 217182 140042 217242 140556
rect 264605 140528 264610 140584
rect 264666 140528 268516 140584
rect 264605 140526 268516 140528
rect 264605 140523 264671 140526
rect 268510 140524 268516 140526
rect 268580 140524 268586 140588
rect 430573 140586 430639 140589
rect 428230 140584 430639 140586
rect 428230 140528 430578 140584
rect 430634 140528 430639 140584
rect 428230 140526 430639 140528
rect 252686 140178 252692 140180
rect 228968 140118 252692 140178
rect 252686 140116 252692 140118
rect 252756 140116 252762 140180
rect 265893 140178 265959 140181
rect 268150 140178 268210 140420
rect 428230 140284 428290 140526
rect 430573 140523 430639 140526
rect 282821 140178 282887 140181
rect 265893 140176 268210 140178
rect 265893 140120 265898 140176
rect 265954 140120 268210 140176
rect 265893 140118 268210 140120
rect 279956 140176 282887 140178
rect 279956 140120 282826 140176
rect 282882 140120 282887 140176
rect 279956 140118 282887 140120
rect 265893 140115 265959 140118
rect 282821 140115 282887 140118
rect 213913 140040 217242 140042
rect 213913 139984 213918 140040
rect 213974 139984 217242 140040
rect 213913 139982 217242 139984
rect 213913 139979 213979 139982
rect 168230 139436 168236 139500
rect 168300 139498 168306 139500
rect 217182 139498 217242 139876
rect 231301 139770 231367 139773
rect 228968 139768 231367 139770
rect 228968 139712 231306 139768
rect 231362 139712 231367 139768
rect 228968 139710 231367 139712
rect 231301 139707 231367 139710
rect 265249 139770 265315 139773
rect 268150 139770 268210 140012
rect 306230 139980 306236 140044
rect 306300 140042 306306 140044
rect 344921 140042 344987 140045
rect 306300 140040 344987 140042
rect 306300 139984 344926 140040
rect 344982 139984 344987 140040
rect 306300 139982 344987 139984
rect 306300 139980 306306 139982
rect 344921 139979 344987 139982
rect 265249 139768 268210 139770
rect 265249 139712 265254 139768
rect 265310 139712 268210 139768
rect 265249 139710 268210 139712
rect 265249 139707 265315 139710
rect 168300 139438 217242 139498
rect 168300 139436 168306 139438
rect 264094 139436 264100 139500
rect 264164 139498 264170 139500
rect 264164 139438 267842 139498
rect 264164 139436 264170 139438
rect 267782 139362 267842 139438
rect 268334 139362 268394 139604
rect 282821 139362 282887 139365
rect 267782 139302 268394 139362
rect 279956 139360 282887 139362
rect 279956 139304 282826 139360
rect 282882 139304 282887 139360
rect 279956 139302 282887 139304
rect 282821 139299 282887 139302
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 231301 139226 231367 139229
rect 228968 139224 231367 139226
rect 213913 138818 213979 138821
rect 217182 138818 217242 139196
rect 228968 139168 231306 139224
rect 231362 139168 231367 139224
rect 347129 139226 347195 139229
rect 347129 139224 350060 139226
rect 228968 139166 231367 139168
rect 231301 139163 231367 139166
rect 231761 138818 231827 138821
rect 213913 138816 217242 138818
rect 213913 138760 213918 138816
rect 213974 138760 217242 138816
rect 213913 138758 217242 138760
rect 228968 138816 231827 138818
rect 228968 138760 231766 138816
rect 231822 138760 231827 138816
rect 228968 138758 231827 138760
rect 213913 138755 213979 138758
rect 231761 138755 231827 138758
rect 265433 138818 265499 138821
rect 268150 138818 268210 139196
rect 347129 139168 347134 139224
rect 347190 139168 350060 139224
rect 583520 139212 584960 139302
rect 347129 139166 350060 139168
rect 347129 139163 347195 139166
rect 428046 138954 428106 139196
rect 429469 138954 429535 138957
rect 429745 138954 429811 138957
rect 428046 138952 429811 138954
rect 428046 138896 429474 138952
rect 429530 138896 429750 138952
rect 429806 138896 429811 138952
rect 428046 138894 429811 138896
rect 429469 138891 429535 138894
rect 429745 138891 429811 138894
rect 265433 138816 268210 138818
rect 265433 138760 265438 138816
rect 265494 138760 268210 138816
rect 265433 138758 268210 138760
rect 265433 138755 265499 138758
rect 213361 138138 213427 138141
rect 217182 138138 217242 138652
rect 265157 138410 265223 138413
rect 268150 138410 268210 138652
rect 282729 138546 282795 138549
rect 279956 138544 282795 138546
rect 279956 138488 282734 138544
rect 282790 138488 282795 138544
rect 279956 138486 282795 138488
rect 282729 138483 282795 138486
rect 265157 138408 268210 138410
rect 265157 138352 265162 138408
rect 265218 138352 268210 138408
rect 265157 138350 268210 138352
rect 265157 138347 265223 138350
rect 231485 138274 231551 138277
rect 228968 138272 231551 138274
rect 228968 138216 231490 138272
rect 231546 138216 231551 138272
rect 228968 138214 231551 138216
rect 231485 138211 231551 138214
rect 264421 138274 264487 138277
rect 264421 138272 268026 138274
rect 264421 138216 264426 138272
rect 264482 138216 268026 138272
rect 264421 138214 268026 138216
rect 264421 138211 264487 138214
rect 213361 138136 217242 138138
rect 213361 138080 213366 138136
rect 213422 138080 217242 138136
rect 267966 138172 268026 138214
rect 268334 138172 268394 138244
rect 267966 138112 268394 138172
rect 213361 138078 217242 138080
rect 213361 138075 213427 138078
rect 217182 137458 217242 137972
rect 267966 137942 268210 138002
rect 230105 137866 230171 137869
rect 228968 137864 230171 137866
rect 228968 137808 230110 137864
rect 230166 137808 230171 137864
rect 228968 137806 230171 137808
rect 230105 137803 230171 137806
rect 264421 137866 264487 137869
rect 267966 137866 268026 137942
rect 264421 137864 268026 137866
rect 264421 137808 264426 137864
rect 264482 137808 268026 137864
rect 268150 137836 268210 137942
rect 282821 137866 282887 137869
rect 279956 137864 282887 137866
rect 264421 137806 268026 137808
rect 279956 137808 282826 137864
rect 282882 137808 282887 137864
rect 279956 137806 282887 137808
rect 264421 137803 264487 137806
rect 282821 137803 282887 137806
rect 428230 137730 428290 137972
rect 430573 137730 430639 137733
rect 428230 137728 430639 137730
rect 428230 137672 430578 137728
rect 430634 137672 430639 137728
rect 428230 137670 430639 137672
rect 430573 137667 430639 137670
rect 267966 137534 268210 137594
rect 200070 137398 217242 137458
rect 262949 137458 263015 137461
rect 267966 137458 268026 137534
rect 262949 137456 268026 137458
rect 262949 137400 262954 137456
rect 263010 137400 268026 137456
rect 268150 137428 268210 137534
rect 346669 137458 346735 137461
rect 430849 137458 430915 137461
rect 346669 137456 350060 137458
rect 262949 137398 268026 137400
rect 346669 137400 346674 137456
rect 346730 137400 350060 137456
rect 346669 137398 350060 137400
rect 428230 137456 430915 137458
rect 428230 137400 430854 137456
rect 430910 137400 430915 137456
rect 428230 137398 430915 137400
rect -960 136778 480 136868
rect 168966 136852 168972 136916
rect 169036 136914 169042 136916
rect 200070 136914 200130 137398
rect 262949 137395 263015 137398
rect 346669 137395 346735 137398
rect 231393 137322 231459 137325
rect 228968 137320 231459 137322
rect 169036 136854 200130 136914
rect 169036 136852 169042 136854
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 214557 136778 214623 136781
rect 217182 136778 217242 137292
rect 228968 137264 231398 137320
rect 231454 137264 231459 137320
rect 228968 137262 231459 137264
rect 231393 137259 231459 137262
rect 267966 137126 268210 137186
rect 266077 137050 266143 137053
rect 267966 137050 268026 137126
rect 266077 137048 268026 137050
rect 266077 136992 266082 137048
rect 266138 136992 268026 137048
rect 268150 137020 268210 137126
rect 282269 137050 282335 137053
rect 279956 137048 282335 137050
rect 266077 136990 268026 136992
rect 279956 136992 282274 137048
rect 282330 136992 282335 137048
rect 279956 136990 282335 136992
rect 266077 136987 266143 136990
rect 282269 136987 282335 136990
rect 231761 136914 231827 136917
rect 228968 136912 231827 136914
rect 228968 136856 231766 136912
rect 231822 136856 231827 136912
rect 428230 136884 428290 137398
rect 430849 137395 430915 137398
rect 228968 136854 231827 136856
rect 231761 136851 231827 136854
rect 214557 136776 217242 136778
rect 214557 136720 214562 136776
rect 214618 136720 217242 136776
rect 214557 136718 217242 136720
rect 214557 136715 214623 136718
rect 260925 136642 260991 136645
rect 267966 136642 268210 136676
rect 260925 136640 268210 136642
rect 214005 136098 214071 136101
rect 217182 136098 217242 136612
rect 260925 136584 260930 136640
rect 260986 136616 268210 136640
rect 260986 136584 268026 136616
rect 268150 136612 268210 136616
rect 260925 136582 268026 136584
rect 260925 136579 260991 136582
rect 231894 136370 231900 136372
rect 228968 136310 231900 136370
rect 231894 136308 231900 136310
rect 231964 136308 231970 136372
rect 280153 136370 280219 136373
rect 430573 136370 430639 136373
rect 267966 136310 268210 136370
rect 279956 136368 280219 136370
rect 279956 136312 280158 136368
rect 280214 136312 280219 136368
rect 279956 136310 280219 136312
rect 261109 136234 261175 136237
rect 267966 136234 268026 136310
rect 261109 136232 268026 136234
rect 261109 136176 261114 136232
rect 261170 136176 268026 136232
rect 268150 136204 268210 136310
rect 280153 136307 280219 136310
rect 428230 136368 430639 136370
rect 428230 136312 430578 136368
rect 430634 136312 430639 136368
rect 428230 136310 430639 136312
rect 261109 136174 268026 136176
rect 261109 136171 261175 136174
rect 214005 136096 217242 136098
rect 214005 136040 214010 136096
rect 214066 136040 217242 136096
rect 214005 136038 217242 136040
rect 214005 136035 214071 136038
rect 231393 135962 231459 135965
rect 228968 135960 231459 135962
rect 214649 135554 214715 135557
rect 217182 135554 217242 135932
rect 228968 135904 231398 135960
rect 231454 135904 231459 135960
rect 228968 135902 231459 135904
rect 231393 135899 231459 135902
rect 264421 135962 264487 135965
rect 264421 135960 268578 135962
rect 264421 135904 264426 135960
rect 264482 135904 268578 135960
rect 264421 135902 268578 135904
rect 264421 135899 264487 135902
rect 268518 135660 268578 135902
rect 347497 135826 347563 135829
rect 347497 135824 350060 135826
rect 347497 135768 347502 135824
rect 347558 135768 350060 135824
rect 428230 135796 428290 136310
rect 430573 136307 430639 136310
rect 347497 135766 350060 135768
rect 347497 135763 347563 135766
rect 282361 135554 282427 135557
rect 214649 135552 217242 135554
rect 214649 135496 214654 135552
rect 214710 135496 217242 135552
rect 214649 135494 217242 135496
rect 279956 135552 282427 135554
rect 279956 135496 282366 135552
rect 282422 135496 282427 135552
rect 279956 135494 282427 135496
rect 214649 135491 214715 135494
rect 282361 135491 282427 135494
rect 213913 135418 213979 135421
rect 230749 135418 230815 135421
rect 213913 135416 217242 135418
rect 213913 135360 213918 135416
rect 213974 135360 217242 135416
rect 213913 135358 217242 135360
rect 228968 135416 230815 135418
rect 228968 135360 230754 135416
rect 230810 135360 230815 135416
rect 228968 135358 230815 135360
rect 213913 135355 213979 135358
rect 217182 135252 217242 135358
rect 230749 135355 230815 135358
rect 265801 135418 265867 135421
rect 265801 135416 268210 135418
rect 265801 135360 265806 135416
rect 265862 135360 268210 135416
rect 265801 135358 268210 135360
rect 265801 135355 265867 135358
rect 268150 135252 268210 135358
rect 231761 135010 231827 135013
rect 430573 135010 430639 135013
rect 228968 135008 231827 135010
rect 228968 134952 231766 135008
rect 231822 134952 231827 135008
rect 228968 134950 231827 134952
rect 231761 134947 231827 134950
rect 428230 135008 430639 135010
rect 428230 134952 430578 135008
rect 430634 134952 430639 135008
rect 428230 134950 430639 134952
rect 265801 134602 265867 134605
rect 268150 134602 268210 134844
rect 282821 134738 282887 134741
rect 279956 134736 282887 134738
rect 279956 134680 282826 134736
rect 282882 134680 282887 134736
rect 428230 134708 428290 134950
rect 430573 134947 430639 134950
rect 279956 134678 282887 134680
rect 282821 134675 282887 134678
rect 265801 134600 268210 134602
rect 166390 134132 166396 134196
rect 166460 134194 166466 134196
rect 217182 134194 217242 134572
rect 265801 134544 265806 134600
rect 265862 134544 268210 134600
rect 265801 134542 268210 134544
rect 265801 134539 265867 134542
rect 231669 134466 231735 134469
rect 228968 134464 231735 134466
rect 228968 134408 231674 134464
rect 231730 134408 231735 134464
rect 228968 134406 231735 134408
rect 231669 134403 231735 134406
rect 166460 134134 217242 134194
rect 265709 134194 265775 134197
rect 268150 134194 268210 134436
rect 305494 134404 305500 134468
rect 305564 134466 305570 134468
rect 338297 134466 338363 134469
rect 305564 134464 338363 134466
rect 305564 134408 338302 134464
rect 338358 134408 338363 134464
rect 305564 134406 338363 134408
rect 305564 134404 305570 134406
rect 338297 134403 338363 134406
rect 265709 134192 268210 134194
rect 265709 134136 265714 134192
rect 265770 134136 268210 134192
rect 265709 134134 268210 134136
rect 166460 134132 166466 134134
rect 265709 134131 265775 134134
rect 213913 134058 213979 134061
rect 230565 134058 230631 134061
rect 282729 134058 282795 134061
rect 213913 134056 217242 134058
rect 213913 134000 213918 134056
rect 213974 134000 217242 134056
rect 213913 133998 217242 134000
rect 228968 134056 230631 134058
rect 228968 134000 230570 134056
rect 230626 134000 230631 134056
rect 279956 134056 282795 134058
rect 228968 133998 230631 134000
rect 213913 133995 213979 133998
rect 217182 133892 217242 133998
rect 230565 133995 230631 133998
rect 265525 133922 265591 133925
rect 265525 133920 267842 133922
rect 265525 133864 265530 133920
rect 265586 133864 267842 133920
rect 265525 133862 267842 133864
rect 265525 133859 265591 133862
rect 267782 133786 267842 133862
rect 268334 133786 268394 134028
rect 279956 134000 282734 134056
rect 282790 134000 282795 134056
rect 279956 133998 282795 134000
rect 282729 133995 282795 133998
rect 338297 134058 338363 134061
rect 338297 134056 350060 134058
rect 338297 134000 338302 134056
rect 338358 134000 350060 134056
rect 338297 133998 350060 134000
rect 338297 133995 338363 133998
rect 428457 133786 428523 133789
rect 430573 133786 430639 133789
rect 267782 133726 268394 133786
rect 428230 133784 430639 133786
rect 428230 133728 428462 133784
rect 428518 133728 430578 133784
rect 430634 133728 430639 133784
rect 428230 133726 430639 133728
rect 231761 133514 231827 133517
rect 228968 133512 231827 133514
rect 228968 133456 231766 133512
rect 231822 133456 231827 133512
rect 228968 133454 231827 133456
rect 231761 133451 231827 133454
rect 214005 132834 214071 132837
rect 217182 132834 217242 133348
rect 265893 133242 265959 133245
rect 268150 133242 268210 133620
rect 428230 133484 428290 133726
rect 428457 133723 428523 133726
rect 430573 133723 430639 133726
rect 281993 133242 282059 133245
rect 265893 133240 268210 133242
rect 265893 133184 265898 133240
rect 265954 133184 268210 133240
rect 265893 133182 268210 133184
rect 279956 133240 282059 133242
rect 279956 133184 281998 133240
rect 282054 133184 282059 133240
rect 279956 133182 282059 133184
rect 265893 133179 265959 133182
rect 281993 133179 282059 133182
rect 231669 133106 231735 133109
rect 228968 133104 231735 133106
rect 228968 133048 231674 133104
rect 231730 133048 231735 133104
rect 228968 133046 231735 133048
rect 231669 133043 231735 133046
rect 214005 132832 217242 132834
rect 214005 132776 214010 132832
rect 214066 132776 217242 132832
rect 214005 132774 217242 132776
rect 265709 132834 265775 132837
rect 268150 132834 268210 133076
rect 265709 132832 268210 132834
rect 265709 132776 265714 132832
rect 265770 132776 268210 132832
rect 265709 132774 268210 132776
rect 214005 132771 214071 132774
rect 265709 132771 265775 132774
rect 213913 132562 213979 132565
rect 213913 132560 216874 132562
rect 213913 132504 213918 132560
rect 213974 132510 216874 132560
rect 217366 132510 217426 132668
rect 231577 132562 231643 132565
rect 213974 132504 217426 132510
rect 213913 132502 217426 132504
rect 228968 132560 231643 132562
rect 228968 132504 231582 132560
rect 231638 132504 231643 132560
rect 228968 132502 231643 132504
rect 213913 132499 213979 132502
rect 216814 132450 217426 132502
rect 231577 132499 231643 132502
rect 265801 132562 265867 132565
rect 265801 132560 267842 132562
rect 265801 132504 265806 132560
rect 265862 132504 267842 132560
rect 265801 132502 267842 132504
rect 265801 132499 265867 132502
rect 267782 132426 267842 132502
rect 268334 132426 268394 132668
rect 282269 132426 282335 132429
rect 267782 132366 268394 132426
rect 279956 132424 282335 132426
rect 279956 132368 282274 132424
rect 282330 132368 282335 132424
rect 279956 132366 282335 132368
rect 282269 132363 282335 132366
rect 347405 132426 347471 132429
rect 347405 132424 350060 132426
rect 347405 132368 347410 132424
rect 347466 132368 350060 132424
rect 347405 132366 350060 132368
rect 347405 132363 347471 132366
rect 230657 132154 230723 132157
rect 228968 132152 230723 132154
rect 228968 132096 230662 132152
rect 230718 132096 230723 132152
rect 228968 132094 230723 132096
rect 230657 132091 230723 132094
rect 265893 132018 265959 132021
rect 268150 132018 268210 132260
rect 428046 132154 428106 132396
rect 430573 132154 430639 132157
rect 428046 132152 430639 132154
rect 428046 132096 430578 132152
rect 430634 132096 430639 132152
rect 428046 132094 430639 132096
rect 430573 132091 430639 132094
rect 265893 132016 268210 132018
rect 213913 131474 213979 131477
rect 217182 131474 217242 131988
rect 265893 131960 265898 132016
rect 265954 131960 268210 132016
rect 265893 131958 268210 131960
rect 265893 131955 265959 131958
rect 430849 131882 430915 131885
rect 428230 131880 430915 131882
rect 231669 131610 231735 131613
rect 228968 131608 231735 131610
rect 228968 131552 231674 131608
rect 231730 131552 231735 131608
rect 228968 131550 231735 131552
rect 231669 131547 231735 131550
rect 265709 131610 265775 131613
rect 268150 131610 268210 131852
rect 428230 131824 430854 131880
rect 430910 131824 430915 131880
rect 428230 131822 430915 131824
rect 282821 131746 282887 131749
rect 279956 131744 282887 131746
rect 279956 131688 282826 131744
rect 282882 131688 282887 131744
rect 279956 131686 282887 131688
rect 282821 131683 282887 131686
rect 265709 131608 268210 131610
rect 265709 131552 265714 131608
rect 265770 131552 268210 131608
rect 265709 131550 268210 131552
rect 265709 131547 265775 131550
rect 213913 131472 217242 131474
rect 213913 131416 213918 131472
rect 213974 131416 217242 131472
rect 213913 131414 217242 131416
rect 213913 131411 213979 131414
rect 173014 131140 173020 131204
rect 173084 131202 173090 131204
rect 173084 131142 216874 131202
rect 173084 131140 173090 131142
rect 216814 131066 216874 131142
rect 217366 131066 217426 131308
rect 231761 131202 231827 131205
rect 228968 131200 231827 131202
rect 228968 131144 231766 131200
rect 231822 131144 231827 131200
rect 228968 131142 231827 131144
rect 231761 131139 231827 131142
rect 265433 131202 265499 131205
rect 268334 131202 268394 131444
rect 428230 131308 428290 131822
rect 430849 131819 430915 131822
rect 265433 131200 268394 131202
rect 265433 131144 265438 131200
rect 265494 131144 268394 131200
rect 265433 131142 268394 131144
rect 265433 131139 265499 131142
rect 216814 131006 217426 131066
rect 231761 130658 231827 130661
rect 268150 130658 268210 131036
rect 294454 131004 294460 131068
rect 294524 131066 294530 131068
rect 349153 131066 349219 131069
rect 294524 131064 349219 131066
rect 294524 131008 349158 131064
rect 349214 131008 349219 131064
rect 294524 131006 349219 131008
rect 294524 131004 294530 131006
rect 349153 131003 349219 131006
rect 281625 130930 281691 130933
rect 279956 130928 281691 130930
rect 279956 130872 281630 130928
rect 281686 130872 281691 130928
rect 279956 130870 281691 130872
rect 281625 130867 281691 130870
rect 430614 130794 430620 130796
rect 428230 130734 430620 130794
rect 228968 130656 231827 130658
rect 166206 130052 166212 130116
rect 166276 130114 166282 130116
rect 217182 130114 217242 130628
rect 228968 130600 231766 130656
rect 231822 130600 231827 130656
rect 228968 130598 231827 130600
rect 231761 130595 231827 130598
rect 258030 130598 268210 130658
rect 349153 130658 349219 130661
rect 349153 130656 350060 130658
rect 349153 130600 349158 130656
rect 349214 130600 350060 130656
rect 349153 130598 350060 130600
rect 231393 130250 231459 130253
rect 228968 130248 231459 130250
rect 228968 130192 231398 130248
rect 231454 130192 231459 130248
rect 228968 130190 231459 130192
rect 231393 130187 231459 130190
rect 257286 130188 257292 130252
rect 257356 130250 257362 130252
rect 258030 130250 258090 130598
rect 349153 130595 349219 130598
rect 257356 130190 258090 130250
rect 265249 130250 265315 130253
rect 268150 130250 268210 130492
rect 265249 130248 268210 130250
rect 265249 130192 265254 130248
rect 265310 130192 268210 130248
rect 428230 130220 428290 130734
rect 430614 130732 430620 130734
rect 430684 130732 430690 130796
rect 265249 130190 268210 130192
rect 257356 130188 257362 130190
rect 265249 130187 265315 130190
rect 281625 130114 281691 130117
rect 166276 130054 217242 130114
rect 279956 130112 281691 130114
rect 166276 130052 166282 130054
rect 169150 129916 169156 129980
rect 169220 129978 169226 129980
rect 169220 129918 216874 129978
rect 169220 129916 169226 129918
rect 216814 129706 216874 129918
rect 217366 129706 217426 129948
rect 231301 129842 231367 129845
rect 228968 129840 231367 129842
rect 228968 129784 231306 129840
rect 231362 129784 231367 129840
rect 228968 129782 231367 129784
rect 231301 129779 231367 129782
rect 262806 129780 262812 129844
rect 262876 129842 262882 129844
rect 268150 129842 268210 130084
rect 279956 130056 281630 130112
rect 281686 130056 281691 130112
rect 279956 130054 281691 130056
rect 281625 130051 281691 130054
rect 262876 129782 268210 129842
rect 262876 129780 262882 129782
rect 216814 129646 217426 129706
rect 268150 129434 268210 129676
rect 430573 129434 430639 129437
rect 258030 129374 268210 129434
rect 428230 129432 430639 129434
rect 66161 129298 66227 129301
rect 68142 129298 68816 129304
rect 231761 129298 231827 129301
rect 66161 129296 68816 129298
rect 66161 129240 66166 129296
rect 66222 129244 68816 129296
rect 228968 129296 231827 129298
rect 66222 129240 68202 129244
rect 66161 129238 68202 129240
rect 66161 129235 66227 129238
rect 214005 128890 214071 128893
rect 217182 128890 217242 129268
rect 228968 129240 231766 129296
rect 231822 129240 231827 129296
rect 228968 129238 231827 129240
rect 231761 129235 231827 129238
rect 244774 128964 244780 129028
rect 244844 129026 244850 129028
rect 258030 129026 258090 129374
rect 244844 128966 258090 129026
rect 244844 128964 244850 128966
rect 265750 128964 265756 129028
rect 265820 129026 265826 129028
rect 268150 129026 268210 129268
rect 265820 128966 268210 129026
rect 265820 128964 265826 128966
rect 231393 128890 231459 128893
rect 214005 128888 217242 128890
rect 214005 128832 214010 128888
rect 214066 128832 217242 128888
rect 214005 128830 217242 128832
rect 228968 128888 231459 128890
rect 228968 128832 231398 128888
rect 231454 128832 231459 128888
rect 228968 128830 231459 128832
rect 214005 128827 214071 128830
rect 231393 128827 231459 128830
rect 213913 128482 213979 128485
rect 217182 128482 217242 128724
rect 265709 128618 265775 128621
rect 268518 128620 268578 128860
rect 279926 128754 279986 129404
rect 428230 129376 430578 129432
rect 430634 129376 430639 129432
rect 428230 129374 430639 129376
rect 428230 128996 428290 129374
rect 430573 129371 430639 129374
rect 288382 128754 288388 128756
rect 279926 128694 288388 128754
rect 288382 128692 288388 128694
rect 288452 128692 288458 128756
rect 265709 128616 268210 128618
rect 265709 128560 265714 128616
rect 265770 128560 268210 128616
rect 265709 128558 268210 128560
rect 265709 128555 265775 128558
rect 213913 128480 217242 128482
rect 213913 128424 213918 128480
rect 213974 128424 217242 128480
rect 268150 128452 268210 128558
rect 268510 128556 268516 128620
rect 268580 128556 268586 128620
rect 282821 128618 282887 128621
rect 279956 128616 282887 128618
rect 279956 128560 282826 128616
rect 282882 128560 282887 128616
rect 279956 128558 282887 128560
rect 282821 128555 282887 128558
rect 350030 128485 350090 128996
rect 347681 128482 347747 128485
rect 349981 128482 350090 128485
rect 347681 128480 350090 128482
rect 213913 128422 217242 128424
rect 347681 128424 347686 128480
rect 347742 128424 349986 128480
rect 350042 128424 350090 128480
rect 347681 128422 350090 128424
rect 213913 128419 213979 128422
rect 347681 128419 347747 128422
rect 349981 128419 350047 128422
rect 231761 128346 231827 128349
rect 228968 128344 231827 128346
rect 228968 128288 231766 128344
rect 231822 128288 231827 128344
rect 228968 128286 231827 128288
rect 231761 128283 231827 128286
rect 427854 128284 427860 128348
rect 427924 128284 427930 128348
rect 264421 128210 264487 128213
rect 268510 128210 268516 128212
rect 264421 128208 268516 128210
rect 264421 128152 264426 128208
rect 264482 128152 268516 128208
rect 264421 128150 268516 128152
rect 264421 128147 264487 128150
rect 268510 128148 268516 128150
rect 268580 128148 268586 128212
rect 66069 128074 66135 128077
rect 68142 128074 68816 128080
rect 66069 128072 68816 128074
rect 66069 128016 66074 128072
rect 66130 128020 68816 128072
rect 66130 128016 68202 128020
rect 66069 128014 68202 128016
rect 66069 128011 66135 128014
rect 214741 127530 214807 127533
rect 217182 127530 217242 128044
rect 231669 127938 231735 127941
rect 228968 127936 231735 127938
rect 228968 127880 231674 127936
rect 231730 127880 231735 127936
rect 427862 127908 427922 128284
rect 228968 127878 231735 127880
rect 231669 127875 231735 127878
rect 249006 127604 249012 127668
rect 249076 127666 249082 127668
rect 268150 127666 268210 127908
rect 281625 127802 281691 127805
rect 279956 127800 281691 127802
rect 279956 127744 281630 127800
rect 281686 127744 281691 127800
rect 279956 127742 281691 127744
rect 281625 127739 281691 127742
rect 249076 127606 268210 127666
rect 249076 127604 249082 127606
rect 214741 127528 217242 127530
rect 214741 127472 214746 127528
rect 214802 127472 217242 127528
rect 214741 127470 217242 127472
rect 214741 127467 214807 127470
rect 231209 127394 231275 127397
rect 228968 127392 231275 127394
rect 170438 127196 170444 127260
rect 170508 127258 170514 127260
rect 170508 127198 200130 127258
rect 170508 127196 170514 127198
rect 200070 127122 200130 127198
rect 217366 127122 217426 127364
rect 228968 127336 231214 127392
rect 231270 127336 231275 127392
rect 228968 127334 231275 127336
rect 231209 127331 231275 127334
rect 265893 127258 265959 127261
rect 268518 127260 268578 127500
rect 347957 127394 348023 127397
rect 348877 127394 348943 127397
rect 347957 127392 350060 127394
rect 347957 127336 347962 127392
rect 348018 127336 348882 127392
rect 348938 127336 350060 127392
rect 347957 127334 350060 127336
rect 347957 127331 348023 127334
rect 348877 127331 348943 127334
rect 265893 127256 268210 127258
rect 265893 127200 265898 127256
rect 265954 127200 268210 127256
rect 265893 127198 268210 127200
rect 265893 127195 265959 127198
rect 200070 127062 217426 127122
rect 268150 127092 268210 127198
rect 268510 127196 268516 127260
rect 268580 127196 268586 127260
rect 282269 127122 282335 127125
rect 279956 127120 282335 127122
rect 279956 127064 282274 127120
rect 282330 127064 282335 127120
rect 279956 127062 282335 127064
rect 282269 127059 282335 127062
rect 231761 126986 231827 126989
rect 429142 126986 429148 126988
rect 228968 126984 231827 126986
rect 228968 126928 231766 126984
rect 231822 126928 231827 126984
rect 228968 126926 231827 126928
rect 231761 126923 231827 126926
rect 428230 126926 429148 126986
rect 264421 126850 264487 126853
rect 268510 126850 268516 126852
rect 264421 126848 268516 126850
rect 264421 126792 264426 126848
rect 264482 126792 268516 126848
rect 264421 126790 268516 126792
rect 264421 126787 264487 126790
rect 268510 126788 268516 126790
rect 268580 126788 268586 126852
rect 428230 126820 428290 126926
rect 429142 126924 429148 126926
rect 429212 126924 429218 126988
rect 65149 126306 65215 126309
rect 68142 126306 68816 126312
rect 65149 126304 68816 126306
rect 65149 126248 65154 126304
rect 65210 126252 68816 126304
rect 65210 126248 68202 126252
rect 65149 126246 68202 126248
rect 65149 126243 65215 126246
rect 214005 126170 214071 126173
rect 217182 126170 217242 126684
rect 231669 126442 231735 126445
rect 228968 126440 231735 126442
rect 228968 126384 231674 126440
rect 231730 126384 231735 126440
rect 228968 126382 231735 126384
rect 231669 126379 231735 126382
rect 260046 126380 260052 126444
rect 260116 126442 260122 126444
rect 268150 126442 268210 126684
rect 260116 126382 268210 126442
rect 260116 126380 260122 126382
rect 282821 126306 282887 126309
rect 428089 126306 428155 126309
rect 279956 126304 282887 126306
rect 214005 126168 217242 126170
rect 214005 126112 214010 126168
rect 214066 126112 217242 126168
rect 214005 126110 217242 126112
rect 214005 126107 214071 126110
rect 231117 126034 231183 126037
rect 228968 126032 231183 126034
rect 213913 125762 213979 125765
rect 217182 125762 217242 126004
rect 228968 125976 231122 126032
rect 231178 125976 231183 126032
rect 228968 125974 231183 125976
rect 231117 125971 231183 125974
rect 265893 126034 265959 126037
rect 268150 126034 268210 126276
rect 279956 126248 282826 126304
rect 282882 126248 282887 126304
rect 279956 126246 282887 126248
rect 282821 126243 282887 126246
rect 428046 126304 428155 126306
rect 428046 126248 428094 126304
rect 428150 126248 428155 126304
rect 428046 126243 428155 126248
rect 265893 126032 268210 126034
rect 265893 125976 265898 126032
rect 265954 125976 268210 126032
rect 265893 125974 268210 125976
rect 265893 125971 265959 125974
rect 232446 125836 232452 125900
rect 232516 125898 232522 125900
rect 232516 125838 258090 125898
rect 232516 125836 232522 125838
rect 213913 125760 217242 125762
rect 213913 125704 213918 125760
rect 213974 125704 217242 125760
rect 213913 125702 217242 125704
rect 213913 125699 213979 125702
rect 258030 125626 258090 125838
rect 268150 125626 268210 125868
rect 428046 125732 428106 126243
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 258030 125566 268210 125626
rect 347681 125626 347747 125629
rect 347681 125624 350060 125626
rect 347681 125568 347686 125624
rect 347742 125568 350060 125624
rect 347681 125566 350060 125568
rect 347681 125563 347747 125566
rect 231577 125490 231643 125493
rect 282821 125490 282887 125493
rect 228968 125488 231643 125490
rect 228968 125432 231582 125488
rect 231638 125432 231643 125488
rect 228968 125430 231643 125432
rect 279956 125488 282887 125490
rect 279956 125432 282826 125488
rect 282882 125432 282887 125488
rect 279956 125430 282887 125432
rect 231577 125427 231643 125430
rect 282821 125427 282887 125430
rect 67633 125218 67699 125221
rect 68142 125218 68816 125224
rect 67633 125216 68816 125218
rect 67633 125160 67638 125216
rect 67694 125164 68816 125216
rect 67694 125160 68202 125164
rect 67633 125158 68202 125160
rect 67633 125155 67699 125158
rect 214005 124810 214071 124813
rect 217182 124810 217242 125324
rect 231301 125082 231367 125085
rect 228968 125080 231367 125082
rect 228968 125024 231306 125080
rect 231362 125024 231367 125080
rect 228968 125022 231367 125024
rect 231301 125019 231367 125022
rect 267273 125082 267339 125085
rect 268150 125082 268210 125324
rect 430573 125082 430639 125085
rect 267273 125080 268210 125082
rect 267273 125024 267278 125080
rect 267334 125024 268210 125080
rect 267273 125022 268210 125024
rect 428230 125080 430639 125082
rect 428230 125024 430578 125080
rect 430634 125024 430639 125080
rect 428230 125022 430639 125024
rect 267273 125019 267339 125022
rect 214005 124808 217242 124810
rect 214005 124752 214010 124808
rect 214066 124752 217242 124808
rect 214005 124750 217242 124752
rect 231761 124810 231827 124813
rect 239254 124810 239260 124812
rect 231761 124808 239260 124810
rect 231761 124752 231766 124808
rect 231822 124752 239260 124808
rect 231761 124750 239260 124752
rect 214005 124747 214071 124750
rect 231761 124747 231827 124750
rect 239254 124748 239260 124750
rect 239324 124748 239330 124812
rect 264421 124674 264487 124677
rect 268150 124674 268210 124916
rect 285622 124810 285628 124812
rect 279956 124750 285628 124810
rect 285622 124748 285628 124750
rect 285692 124748 285698 124812
rect 264421 124672 268210 124674
rect 213913 124402 213979 124405
rect 217182 124402 217242 124644
rect 264421 124616 264426 124672
rect 264482 124616 268210 124672
rect 264421 124614 268210 124616
rect 264421 124611 264487 124614
rect 231669 124538 231735 124541
rect 228968 124536 231735 124538
rect 228968 124480 231674 124536
rect 231730 124480 231735 124536
rect 428230 124508 428290 125022
rect 430573 125019 430639 125022
rect 228968 124478 231735 124480
rect 231669 124475 231735 124478
rect 213913 124400 217242 124402
rect 213913 124344 213918 124400
rect 213974 124344 217242 124400
rect 213913 124342 217242 124344
rect 213913 124339 213979 124342
rect 265893 124266 265959 124269
rect 268150 124266 268210 124508
rect 265893 124264 268210 124266
rect 265893 124208 265898 124264
rect 265954 124208 268210 124264
rect 265893 124206 268210 124208
rect 265893 124203 265959 124206
rect 231761 124130 231827 124133
rect 228968 124128 231827 124130
rect -960 123572 480 123812
rect 67541 123586 67607 123589
rect 68142 123586 68816 123592
rect 67541 123584 68816 123586
rect 67541 123528 67546 123584
rect 67602 123532 68816 123584
rect 214005 123586 214071 123589
rect 217182 123586 217242 124100
rect 228968 124072 231766 124128
rect 231822 124072 231827 124128
rect 228968 124070 231827 124072
rect 231761 124067 231827 124070
rect 265985 123858 266051 123861
rect 268150 123858 268210 124100
rect 285806 123994 285812 123996
rect 279956 123934 285812 123994
rect 285806 123932 285812 123934
rect 285876 123932 285882 123996
rect 348969 123994 349035 123997
rect 348969 123992 350060 123994
rect 348969 123936 348974 123992
rect 349030 123936 350060 123992
rect 348969 123934 350060 123936
rect 348969 123931 349035 123934
rect 430573 123858 430639 123861
rect 265985 123856 268210 123858
rect 265985 123800 265990 123856
rect 266046 123800 268210 123856
rect 265985 123798 268210 123800
rect 428230 123856 430639 123858
rect 428230 123800 430578 123856
rect 430634 123800 430639 123856
rect 428230 123798 430639 123800
rect 265985 123795 266051 123798
rect 231301 123586 231367 123589
rect 214005 123584 217242 123586
rect 67602 123528 68202 123532
rect 67541 123526 68202 123528
rect 214005 123528 214010 123584
rect 214066 123528 217242 123584
rect 214005 123526 217242 123528
rect 228968 123584 231367 123586
rect 228968 123528 231306 123584
rect 231362 123528 231367 123584
rect 228968 123526 231367 123528
rect 67541 123523 67607 123526
rect 214005 123523 214071 123526
rect 231301 123523 231367 123526
rect 265893 123450 265959 123453
rect 268150 123450 268210 123692
rect 265893 123448 268210 123450
rect 213913 122906 213979 122909
rect 217182 122906 217242 123420
rect 265893 123392 265898 123448
rect 265954 123392 268210 123448
rect 428230 123420 428290 123798
rect 430573 123795 430639 123798
rect 265893 123390 268210 123392
rect 265893 123387 265959 123390
rect 231485 123178 231551 123181
rect 228968 123176 231551 123178
rect 228968 123120 231490 123176
rect 231546 123120 231551 123176
rect 228968 123118 231551 123120
rect 231485 123115 231551 123118
rect 265893 123042 265959 123045
rect 268518 123044 268578 123284
rect 282177 123178 282243 123181
rect 279956 123176 282243 123178
rect 279956 123120 282182 123176
rect 282238 123120 282243 123176
rect 279956 123118 282243 123120
rect 282177 123115 282243 123118
rect 265893 123040 268210 123042
rect 265893 122984 265898 123040
rect 265954 122984 268210 123040
rect 265893 122982 268210 122984
rect 265893 122979 265959 122982
rect 213913 122904 217242 122906
rect 213913 122848 213918 122904
rect 213974 122848 217242 122904
rect 268150 122876 268210 122982
rect 268510 122980 268516 123044
rect 268580 122980 268586 123044
rect 213913 122846 217242 122848
rect 213913 122843 213979 122846
rect 67357 122634 67423 122637
rect 68142 122634 68816 122640
rect 67357 122632 68816 122634
rect 67357 122576 67362 122632
rect 67418 122580 68816 122632
rect 67418 122576 68202 122580
rect 67357 122574 68202 122576
rect 67357 122571 67423 122574
rect 214005 122226 214071 122229
rect 217182 122226 217242 122740
rect 298686 122708 298692 122772
rect 298756 122770 298762 122772
rect 349061 122770 349127 122773
rect 298756 122768 350090 122770
rect 298756 122712 349066 122768
rect 349122 122712 350090 122768
rect 298756 122710 350090 122712
rect 298756 122708 298762 122710
rect 349061 122707 349127 122710
rect 231577 122634 231643 122637
rect 228968 122632 231643 122634
rect 228968 122576 231582 122632
rect 231638 122576 231643 122632
rect 228968 122574 231643 122576
rect 231577 122571 231643 122574
rect 263133 122634 263199 122637
rect 268510 122634 268516 122636
rect 263133 122632 268516 122634
rect 263133 122576 263138 122632
rect 263194 122576 268516 122632
rect 263133 122574 268516 122576
rect 263133 122571 263199 122574
rect 268510 122572 268516 122574
rect 268580 122572 268586 122636
rect 283005 122498 283071 122501
rect 279956 122496 283071 122498
rect 279956 122440 283010 122496
rect 283066 122440 283071 122496
rect 279956 122438 283071 122440
rect 283005 122435 283071 122438
rect 231761 122226 231827 122229
rect 214005 122224 217242 122226
rect 214005 122168 214010 122224
rect 214066 122168 217242 122224
rect 214005 122166 217242 122168
rect 228968 122224 231827 122226
rect 228968 122168 231766 122224
rect 231822 122168 231827 122224
rect 228968 122166 231827 122168
rect 214005 122163 214071 122166
rect 231761 122163 231827 122166
rect 265985 122090 266051 122093
rect 268150 122090 268210 122332
rect 350030 122196 350090 122710
rect 430573 122634 430639 122637
rect 428230 122632 430639 122634
rect 428230 122576 430578 122632
rect 430634 122576 430639 122632
rect 428230 122574 430639 122576
rect 428230 122332 428290 122574
rect 430573 122571 430639 122574
rect 265985 122088 268210 122090
rect 213913 121818 213979 121821
rect 217182 121818 217242 122060
rect 265985 122032 265990 122088
rect 266046 122032 268210 122088
rect 265985 122030 268210 122032
rect 265985 122027 266051 122030
rect 213913 121816 217242 121818
rect 213913 121760 213918 121816
rect 213974 121760 217242 121816
rect 213913 121758 217242 121760
rect 213913 121755 213979 121758
rect 231485 121682 231551 121685
rect 228968 121680 231551 121682
rect 228968 121624 231490 121680
rect 231546 121624 231551 121680
rect 228968 121622 231551 121624
rect 231485 121619 231551 121622
rect 265893 121682 265959 121685
rect 268518 121684 268578 121924
rect 265893 121680 268210 121682
rect 265893 121624 265898 121680
rect 265954 121624 268210 121680
rect 265893 121622 268210 121624
rect 265893 121619 265959 121622
rect 268150 121516 268210 121622
rect 268510 121620 268516 121684
rect 268580 121620 268586 121684
rect 282821 121682 282887 121685
rect 279956 121680 282887 121682
rect 279956 121624 282826 121680
rect 282882 121624 282887 121680
rect 279956 121622 282887 121624
rect 282821 121619 282887 121622
rect 430573 121410 430639 121413
rect 428230 121408 430639 121410
rect 67449 120866 67515 120869
rect 68142 120866 68816 120872
rect 67449 120864 68816 120866
rect 67449 120808 67454 120864
rect 67510 120812 68816 120864
rect 214005 120866 214071 120869
rect 217182 120866 217242 121380
rect 428230 121352 430578 121408
rect 430634 121352 430639 121408
rect 428230 121350 430639 121352
rect 231761 121274 231827 121277
rect 228968 121272 231827 121274
rect 228968 121216 231766 121272
rect 231822 121216 231827 121272
rect 228968 121214 231827 121216
rect 231761 121211 231827 121214
rect 264237 121274 264303 121277
rect 268510 121274 268516 121276
rect 264237 121272 268516 121274
rect 264237 121216 264242 121272
rect 264298 121216 268516 121272
rect 264237 121214 268516 121216
rect 264237 121211 264303 121214
rect 268510 121212 268516 121214
rect 268580 121212 268586 121276
rect 428230 121244 428290 121350
rect 430573 121347 430639 121350
rect 214005 120864 217242 120866
rect 67510 120808 68202 120812
rect 67449 120806 68202 120808
rect 214005 120808 214010 120864
rect 214066 120808 217242 120864
rect 214005 120806 217242 120808
rect 265617 120866 265683 120869
rect 268150 120866 268210 121108
rect 281901 120866 281967 120869
rect 265617 120864 268210 120866
rect 265617 120808 265622 120864
rect 265678 120808 268210 120864
rect 265617 120806 268210 120808
rect 279956 120864 281967 120866
rect 279956 120808 281906 120864
rect 281962 120808 281967 120864
rect 279956 120806 281967 120808
rect 67449 120803 67515 120806
rect 214005 120803 214071 120806
rect 265617 120803 265683 120806
rect 281901 120803 281967 120806
rect 231117 120730 231183 120733
rect 228968 120728 231183 120730
rect 213913 120186 213979 120189
rect 217182 120186 217242 120700
rect 228968 120672 231122 120728
rect 231178 120672 231183 120728
rect 228968 120670 231183 120672
rect 231117 120667 231183 120670
rect 265525 120458 265591 120461
rect 268150 120458 268210 120700
rect 430573 120594 430639 120597
rect 428230 120592 430639 120594
rect 265525 120456 268210 120458
rect 265525 120400 265530 120456
rect 265586 120400 268210 120456
rect 265525 120398 268210 120400
rect 265525 120395 265591 120398
rect 231485 120322 231551 120325
rect 228968 120320 231551 120322
rect 228968 120264 231490 120320
rect 231546 120264 231551 120320
rect 228968 120262 231551 120264
rect 231485 120259 231551 120262
rect 213913 120184 217242 120186
rect 213913 120128 213918 120184
rect 213974 120128 217242 120184
rect 213913 120126 217242 120128
rect 265709 120186 265775 120189
rect 265709 120184 267842 120186
rect 265709 120128 265714 120184
rect 265770 120128 267842 120184
rect 265709 120126 267842 120128
rect 213913 120123 213979 120126
rect 265709 120123 265775 120126
rect 267782 120050 267842 120126
rect 268334 120050 268394 120292
rect 281625 120186 281691 120189
rect 279956 120184 281691 120186
rect 279956 120128 281630 120184
rect 281686 120128 281691 120184
rect 279956 120126 281691 120128
rect 281625 120123 281691 120126
rect 291878 120124 291884 120188
rect 291948 120186 291954 120188
rect 349102 120186 349108 120188
rect 291948 120126 349108 120186
rect 291948 120124 291954 120126
rect 349102 120124 349108 120126
rect 349172 120186 349178 120188
rect 350030 120186 350090 120564
rect 349172 120126 350090 120186
rect 428230 120536 430578 120592
rect 430634 120536 430639 120592
rect 428230 120534 430639 120536
rect 428230 120156 428290 120534
rect 430573 120531 430639 120534
rect 349172 120124 349178 120126
rect 214005 119642 214071 119645
rect 217182 119642 217242 120020
rect 267782 119990 268394 120050
rect 231301 119778 231367 119781
rect 228968 119776 231367 119778
rect 228968 119720 231306 119776
rect 231362 119720 231367 119776
rect 228968 119718 231367 119720
rect 231301 119715 231367 119718
rect 214005 119640 217242 119642
rect 214005 119584 214010 119640
rect 214066 119584 217242 119640
rect 214005 119582 217242 119584
rect 214005 119579 214071 119582
rect 265617 119506 265683 119509
rect 268150 119506 268210 119748
rect 430573 119506 430639 119509
rect 265617 119504 268210 119506
rect 213913 118962 213979 118965
rect 217182 118962 217242 119476
rect 265617 119448 265622 119504
rect 265678 119448 268210 119504
rect 265617 119446 268210 119448
rect 428230 119504 430639 119506
rect 428230 119448 430578 119504
rect 430634 119448 430639 119504
rect 428230 119446 430639 119448
rect 265617 119443 265683 119446
rect 231393 119370 231459 119373
rect 282085 119370 282151 119373
rect 228968 119368 231459 119370
rect 228968 119312 231398 119368
rect 231454 119312 231459 119368
rect 279956 119368 282151 119370
rect 228968 119310 231459 119312
rect 231393 119307 231459 119310
rect 262070 119036 262076 119100
rect 262140 119098 262146 119100
rect 268150 119098 268210 119340
rect 279956 119312 282090 119368
rect 282146 119312 282151 119368
rect 279956 119310 282151 119312
rect 282085 119307 282151 119310
rect 262140 119038 268210 119098
rect 262140 119036 262146 119038
rect 231761 118962 231827 118965
rect 213913 118960 217242 118962
rect 213913 118904 213918 118960
rect 213974 118904 217242 118960
rect 213913 118902 217242 118904
rect 228968 118960 231827 118962
rect 228968 118904 231766 118960
rect 231822 118904 231827 118960
rect 428230 118932 428290 119446
rect 430573 119443 430639 119446
rect 228968 118902 231827 118904
rect 213913 118899 213979 118902
rect 231761 118899 231827 118902
rect 214097 118826 214163 118829
rect 265709 118826 265775 118829
rect 214097 118824 216874 118826
rect 214097 118768 214102 118824
rect 214158 118768 216874 118824
rect 265709 118824 267842 118826
rect 214097 118766 216874 118768
rect 214097 118763 214163 118766
rect 216814 118554 216874 118766
rect 217366 118554 217426 118796
rect 265709 118768 265714 118824
rect 265770 118768 267842 118824
rect 265709 118766 267842 118768
rect 265709 118763 265775 118766
rect 267782 118690 267842 118766
rect 268334 118690 268394 118932
rect 347037 118826 347103 118829
rect 347037 118824 350060 118826
rect 347037 118768 347042 118824
rect 347098 118768 350060 118824
rect 347037 118766 350060 118768
rect 347037 118763 347103 118766
rect 267782 118630 268394 118690
rect 282821 118554 282887 118557
rect 216814 118494 217426 118554
rect 279956 118552 282887 118554
rect 231761 118418 231827 118421
rect 228968 118416 231827 118418
rect 228968 118360 231766 118416
rect 231822 118360 231827 118416
rect 228968 118358 231827 118360
rect 231761 118355 231827 118358
rect 265985 118282 266051 118285
rect 268150 118282 268210 118524
rect 279956 118496 282826 118552
rect 282882 118496 282887 118552
rect 279956 118494 282887 118496
rect 282821 118491 282887 118494
rect 265985 118280 268210 118282
rect 265985 118224 265990 118280
rect 266046 118224 268210 118280
rect 265985 118222 268210 118224
rect 265985 118219 266051 118222
rect 430573 118146 430639 118149
rect 428230 118144 430639 118146
rect 214005 117602 214071 117605
rect 217182 117602 217242 118116
rect 231117 118010 231183 118013
rect 228968 118008 231183 118010
rect 228968 117952 231122 118008
rect 231178 117952 231183 118008
rect 228968 117950 231183 117952
rect 231117 117947 231183 117950
rect 265341 117874 265407 117877
rect 268150 117874 268210 118116
rect 428230 118088 430578 118144
rect 430634 118088 430639 118144
rect 428230 118086 430639 118088
rect 282453 117874 282519 117877
rect 265341 117872 268210 117874
rect 265341 117816 265346 117872
rect 265402 117816 268210 117872
rect 265341 117814 268210 117816
rect 279956 117872 282519 117874
rect 279956 117816 282458 117872
rect 282514 117816 282519 117872
rect 428230 117844 428290 118086
rect 430573 118083 430639 118086
rect 279956 117814 282519 117816
rect 265341 117811 265407 117814
rect 282453 117811 282519 117814
rect 214005 117600 217242 117602
rect 214005 117544 214010 117600
rect 214066 117544 217242 117600
rect 214005 117542 217242 117544
rect 214005 117539 214071 117542
rect 231485 117466 231551 117469
rect 228968 117464 231551 117466
rect 213913 117330 213979 117333
rect 213913 117328 216874 117330
rect 213913 117272 213918 117328
rect 213974 117272 216874 117328
rect 213913 117270 216874 117272
rect 213913 117267 213979 117270
rect 216814 117194 216874 117270
rect 217366 117194 217426 117436
rect 228968 117408 231490 117464
rect 231546 117408 231551 117464
rect 228968 117406 231551 117408
rect 231485 117403 231551 117406
rect 265709 117466 265775 117469
rect 268150 117466 268210 117708
rect 265709 117464 268210 117466
rect 265709 117408 265714 117464
rect 265770 117408 268210 117464
rect 265709 117406 268210 117408
rect 265709 117403 265775 117406
rect 265617 117330 265683 117333
rect 268510 117330 268516 117332
rect 265617 117328 268516 117330
rect 265617 117272 265622 117328
rect 265678 117272 268516 117328
rect 265617 117270 268516 117272
rect 265617 117267 265683 117270
rect 268510 117268 268516 117270
rect 268580 117268 268586 117332
rect 216814 117134 217426 117194
rect 347313 117194 347379 117197
rect 347313 117192 350060 117194
rect 231158 117058 231164 117060
rect 228968 116998 231164 117058
rect 231158 116996 231164 116998
rect 231228 116996 231234 117060
rect 266077 116922 266143 116925
rect 268150 116922 268210 117164
rect 347313 117136 347318 117192
rect 347374 117136 350060 117192
rect 347313 117134 350060 117136
rect 347313 117131 347379 117134
rect 280286 117058 280292 117060
rect 279956 116998 280292 117058
rect 280286 116996 280292 116998
rect 280356 116996 280362 117060
rect 430573 117058 430639 117061
rect 428230 117056 430639 117058
rect 428230 117000 430578 117056
rect 430634 117000 430639 117056
rect 428230 116998 430639 117000
rect 266077 116920 268210 116922
rect 266077 116864 266082 116920
rect 266138 116864 268210 116920
rect 266077 116862 268210 116864
rect 266077 116859 266143 116862
rect 428230 116756 428290 116998
rect 430573 116995 430639 116998
rect 214005 116242 214071 116245
rect 217182 116242 217242 116756
rect 231485 116514 231551 116517
rect 228968 116512 231551 116514
rect 228968 116456 231490 116512
rect 231546 116456 231551 116512
rect 228968 116454 231551 116456
rect 231485 116451 231551 116454
rect 265985 116514 266051 116517
rect 268150 116514 268210 116756
rect 265985 116512 268210 116514
rect 265985 116456 265990 116512
rect 266046 116456 268210 116512
rect 265985 116454 268210 116456
rect 265985 116451 266051 116454
rect 268510 116452 268516 116516
rect 268580 116452 268586 116516
rect 268518 116348 268578 116452
rect 282545 116378 282611 116381
rect 279956 116376 282611 116378
rect 279956 116320 282550 116376
rect 282606 116320 282611 116376
rect 279956 116318 282611 116320
rect 282545 116315 282611 116318
rect 214005 116240 217242 116242
rect 214005 116184 214010 116240
rect 214066 116184 217242 116240
rect 214005 116182 217242 116184
rect 214005 116179 214071 116182
rect 231669 116106 231735 116109
rect 228968 116104 231735 116106
rect 213913 115970 213979 115973
rect 213913 115968 216874 115970
rect 213913 115912 213918 115968
rect 213974 115912 216874 115968
rect 213913 115910 216874 115912
rect 213913 115907 213979 115910
rect 216814 115834 216874 115910
rect 217366 115834 217426 116076
rect 228968 116048 231674 116104
rect 231730 116048 231735 116104
rect 228968 116046 231735 116048
rect 231669 116043 231735 116046
rect 265709 116106 265775 116109
rect 265709 116104 268210 116106
rect 265709 116048 265714 116104
rect 265770 116048 268210 116104
rect 265709 116046 268210 116048
rect 265709 116043 265775 116046
rect 268150 115940 268210 116046
rect 430573 115834 430639 115837
rect 216814 115774 217426 115834
rect 428230 115832 430639 115834
rect 428230 115776 430578 115832
rect 430634 115776 430639 115832
rect 428230 115774 430639 115776
rect 428230 115668 428290 115774
rect 430573 115771 430639 115774
rect 230657 115562 230723 115565
rect 282821 115562 282887 115565
rect 228968 115560 230723 115562
rect 228968 115504 230662 115560
rect 230718 115504 230723 115560
rect 279956 115560 282887 115562
rect 228968 115502 230723 115504
rect 230657 115499 230723 115502
rect 214005 115018 214071 115021
rect 217182 115018 217242 115396
rect 265249 115290 265315 115293
rect 268150 115290 268210 115532
rect 279956 115504 282826 115560
rect 282882 115504 282887 115560
rect 279956 115502 282887 115504
rect 282821 115499 282887 115502
rect 347497 115426 347563 115429
rect 347497 115424 350060 115426
rect 347497 115368 347502 115424
rect 347558 115368 350060 115424
rect 347497 115366 350060 115368
rect 347497 115363 347563 115366
rect 265249 115288 268210 115290
rect 265249 115232 265254 115288
rect 265310 115232 268210 115288
rect 265249 115230 268210 115232
rect 265249 115227 265315 115230
rect 231669 115154 231735 115157
rect 228968 115152 231735 115154
rect 228968 115096 231674 115152
rect 231730 115096 231735 115152
rect 228968 115094 231735 115096
rect 231669 115091 231735 115094
rect 214005 115016 217242 115018
rect 214005 114960 214010 115016
rect 214066 114960 217242 115016
rect 214005 114958 217242 114960
rect 214005 114955 214071 114958
rect 265985 114882 266051 114885
rect 268150 114882 268210 115124
rect 265985 114880 268210 114882
rect 213913 114610 213979 114613
rect 217366 114610 217426 114852
rect 265985 114824 265990 114880
rect 266046 114824 268210 114880
rect 265985 114822 268210 114824
rect 265985 114819 266051 114822
rect 265709 114746 265775 114749
rect 282545 114746 282611 114749
rect 265709 114744 268210 114746
rect 265709 114688 265714 114744
rect 265770 114688 268210 114744
rect 265709 114686 268210 114688
rect 279956 114744 282611 114746
rect 279956 114688 282550 114744
rect 282606 114688 282611 114744
rect 279956 114686 282611 114688
rect 265709 114683 265775 114686
rect 230565 114610 230631 114613
rect 213913 114608 217426 114610
rect 213913 114552 213918 114608
rect 213974 114552 217426 114608
rect 213913 114550 217426 114552
rect 228968 114608 230631 114610
rect 228968 114552 230570 114608
rect 230626 114552 230631 114608
rect 268150 114580 268210 114686
rect 282545 114683 282611 114686
rect 228968 114550 230631 114552
rect 213913 114547 213979 114550
rect 230565 114547 230631 114550
rect 231117 114202 231183 114205
rect 228968 114200 231183 114202
rect 214005 113658 214071 113661
rect 217182 113658 217242 114172
rect 228968 114144 231122 114200
rect 231178 114144 231183 114200
rect 428046 114202 428106 114444
rect 430573 114202 430639 114205
rect 428046 114200 430639 114202
rect 228968 114142 231183 114144
rect 231117 114139 231183 114142
rect 265249 113930 265315 113933
rect 268150 113930 268210 114172
rect 428046 114144 430578 114200
rect 430634 114144 430639 114200
rect 428046 114142 430639 114144
rect 430573 114139 430639 114142
rect 281625 114066 281691 114069
rect 279956 114064 281691 114066
rect 279956 114008 281630 114064
rect 281686 114008 281691 114064
rect 279956 114006 281691 114008
rect 281625 114003 281691 114006
rect 430849 113930 430915 113933
rect 265249 113928 268210 113930
rect 265249 113872 265254 113928
rect 265310 113872 268210 113928
rect 265249 113870 268210 113872
rect 428230 113928 430915 113930
rect 428230 113872 430854 113928
rect 430910 113872 430915 113928
rect 428230 113870 430915 113872
rect 265249 113867 265315 113870
rect 231761 113658 231827 113661
rect 214005 113656 217242 113658
rect 214005 113600 214010 113656
rect 214066 113600 217242 113656
rect 214005 113598 217242 113600
rect 228968 113656 231827 113658
rect 228968 113600 231766 113656
rect 231822 113600 231827 113656
rect 228968 113598 231827 113600
rect 214005 113595 214071 113598
rect 231761 113595 231827 113598
rect 265709 113522 265775 113525
rect 268150 113522 268210 113764
rect 265709 113520 268210 113522
rect 213913 113250 213979 113253
rect 217366 113250 217426 113492
rect 265709 113464 265714 113520
rect 265770 113464 268210 113520
rect 265709 113462 268210 113464
rect 265709 113459 265775 113462
rect 230565 113250 230631 113253
rect 213913 113248 217426 113250
rect 213913 113192 213918 113248
rect 213974 113192 217426 113248
rect 213913 113190 217426 113192
rect 228968 113248 230631 113250
rect 228968 113192 230570 113248
rect 230626 113192 230631 113248
rect 228968 113190 230631 113192
rect 213913 113187 213979 113190
rect 230565 113187 230631 113190
rect 265709 113250 265775 113253
rect 265709 113248 267842 113250
rect 265709 113192 265714 113248
rect 265770 113192 267842 113248
rect 265709 113190 267842 113192
rect 265709 113187 265775 113190
rect 267782 113114 267842 113190
rect 268334 113114 268394 113356
rect 280245 113250 280311 113253
rect 279956 113248 280311 113250
rect 279956 113192 280250 113248
rect 280306 113192 280311 113248
rect 279956 113190 280311 113192
rect 280245 113187 280311 113190
rect 302734 113188 302740 113252
rect 302804 113250 302810 113252
rect 350030 113250 350090 113764
rect 428230 113356 428290 113870
rect 430849 113867 430915 113870
rect 302804 113190 350090 113250
rect 302804 113188 302810 113190
rect 267782 113054 268394 113114
rect 214005 112298 214071 112301
rect 217182 112298 217242 112812
rect 231761 112706 231827 112709
rect 228968 112704 231827 112706
rect 228968 112648 231766 112704
rect 231822 112648 231827 112704
rect 228968 112646 231827 112648
rect 231761 112643 231827 112646
rect 262990 112644 262996 112708
rect 263060 112706 263066 112708
rect 268150 112706 268210 112948
rect 580349 112842 580415 112845
rect 583520 112842 584960 112932
rect 580349 112840 584960 112842
rect 580349 112784 580354 112840
rect 580410 112784 584960 112840
rect 580349 112782 584960 112784
rect 580349 112779 580415 112782
rect 430757 112706 430823 112709
rect 263060 112646 268210 112706
rect 428230 112704 430823 112706
rect 428230 112648 430762 112704
rect 430818 112648 430823 112704
rect 583520 112692 584960 112782
rect 428230 112646 430823 112648
rect 263060 112644 263066 112646
rect 231209 112298 231275 112301
rect 214005 112296 217242 112298
rect 214005 112240 214010 112296
rect 214066 112240 217242 112296
rect 214005 112238 217242 112240
rect 228968 112296 231275 112298
rect 228968 112240 231214 112296
rect 231270 112240 231275 112296
rect 228968 112238 231275 112240
rect 214005 112235 214071 112238
rect 231209 112235 231275 112238
rect 264237 112162 264303 112165
rect 268150 112162 268210 112540
rect 282085 112434 282151 112437
rect 279956 112432 282151 112434
rect 279956 112376 282090 112432
rect 282146 112376 282151 112432
rect 279956 112374 282151 112376
rect 282085 112371 282151 112374
rect 428230 112268 428290 112646
rect 430757 112643 430823 112646
rect 264237 112160 268210 112162
rect 213913 111890 213979 111893
rect 217366 111890 217426 112132
rect 264237 112104 264242 112160
rect 264298 112104 268210 112160
rect 264237 112102 268210 112104
rect 264237 112099 264303 112102
rect 213913 111888 217426 111890
rect 213913 111832 213918 111888
rect 213974 111832 217426 111888
rect 213913 111830 217426 111832
rect 265709 111890 265775 111893
rect 265709 111888 267842 111890
rect 265709 111832 265714 111888
rect 265770 111832 267842 111888
rect 265709 111830 267842 111832
rect 213913 111827 213979 111830
rect 265709 111827 265775 111830
rect 167913 111754 167979 111757
rect 237966 111754 237972 111756
rect 164694 111752 167979 111754
rect 164694 111696 167918 111752
rect 167974 111696 167979 111752
rect 164694 111694 167979 111696
rect 228968 111694 237972 111754
rect 167913 111691 167979 111694
rect 237966 111692 237972 111694
rect 238036 111692 238042 111756
rect 267782 111754 267842 111830
rect 268334 111754 268394 111996
rect 293166 111828 293172 111892
rect 293236 111890 293242 111892
rect 350030 111890 350090 112132
rect 293236 111830 350090 111890
rect 293236 111828 293242 111830
rect 267782 111694 268394 111754
rect 214005 110938 214071 110941
rect 217182 110938 217242 111452
rect 231761 111346 231827 111349
rect 228968 111344 231827 111346
rect 228968 111288 231766 111344
rect 231822 111288 231827 111344
rect 228968 111286 231827 111288
rect 231761 111283 231827 111286
rect 265985 111346 266051 111349
rect 268150 111346 268210 111588
rect 265985 111344 268210 111346
rect 265985 111288 265990 111344
rect 266046 111288 268210 111344
rect 265985 111286 268210 111288
rect 265985 111283 266051 111286
rect 214005 110936 217242 110938
rect 214005 110880 214010 110936
rect 214066 110880 217242 110936
rect 214005 110878 217242 110880
rect 264329 110938 264395 110941
rect 268150 110938 268210 111180
rect 279926 111074 279986 111724
rect 430573 111482 430639 111485
rect 428230 111480 430639 111482
rect 428230 111424 430578 111480
rect 430634 111424 430639 111480
rect 428230 111422 430639 111424
rect 428230 111180 428290 111422
rect 430573 111419 430639 111422
rect 279926 111014 287070 111074
rect 282821 110938 282887 110941
rect 264329 110936 268210 110938
rect 264329 110880 264334 110936
rect 264390 110880 268210 110936
rect 264329 110878 268210 110880
rect 279956 110936 282887 110938
rect 279956 110880 282826 110936
rect 282882 110880 282887 110936
rect 279956 110878 282887 110880
rect 214005 110875 214071 110878
rect 264329 110875 264395 110878
rect 282821 110875 282887 110878
rect 231485 110802 231551 110805
rect 228968 110800 231551 110802
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 213913 110530 213979 110533
rect 217182 110530 217242 110772
rect 228968 110744 231490 110800
rect 231546 110744 231551 110800
rect 228968 110742 231551 110744
rect 231485 110739 231551 110742
rect 213913 110528 217242 110530
rect 213913 110472 213918 110528
rect 213974 110472 217242 110528
rect 213913 110470 217242 110472
rect 265709 110530 265775 110533
rect 268150 110530 268210 110772
rect 265709 110528 268210 110530
rect 265709 110472 265714 110528
rect 265770 110472 268210 110528
rect 265709 110470 268210 110472
rect 287010 110530 287070 111014
rect 290590 110530 290596 110532
rect 287010 110470 290596 110530
rect 213913 110467 213979 110470
rect 265709 110467 265775 110470
rect 290590 110468 290596 110470
rect 290660 110468 290666 110532
rect 231761 110394 231827 110397
rect 228968 110392 231827 110394
rect 228968 110336 231766 110392
rect 231822 110336 231827 110392
rect 347037 110394 347103 110397
rect 431861 110394 431927 110397
rect 347037 110392 350060 110394
rect 228968 110334 231827 110336
rect 231761 110331 231827 110334
rect 168097 110122 168163 110125
rect 164694 110120 168163 110122
rect 164694 110064 168102 110120
rect 168158 110064 168163 110120
rect 164694 110062 168163 110064
rect 168097 110059 168163 110062
rect 214005 109714 214071 109717
rect 217182 109714 217242 110228
rect 265709 110122 265775 110125
rect 268150 110122 268210 110364
rect 347037 110336 347042 110392
rect 347098 110336 350060 110392
rect 347037 110334 350060 110336
rect 428230 110392 431927 110394
rect 428230 110336 431866 110392
rect 431922 110336 431927 110392
rect 428230 110334 431927 110336
rect 347037 110331 347103 110334
rect 265709 110120 268210 110122
rect 265709 110064 265714 110120
rect 265770 110064 268210 110120
rect 265709 110062 268210 110064
rect 265709 110059 265775 110062
rect 231761 109850 231827 109853
rect 228968 109848 231827 109850
rect 228968 109792 231766 109848
rect 231822 109792 231827 109848
rect 228968 109790 231827 109792
rect 231761 109787 231827 109790
rect 214005 109712 217242 109714
rect 214005 109656 214010 109712
rect 214066 109656 217242 109712
rect 214005 109654 217242 109656
rect 265157 109714 265223 109717
rect 268150 109714 268210 109956
rect 265157 109712 268210 109714
rect 265157 109656 265162 109712
rect 265218 109656 268210 109712
rect 265157 109654 268210 109656
rect 214005 109651 214071 109654
rect 265157 109651 265223 109654
rect 279926 109578 279986 110092
rect 428230 109956 428290 110334
rect 431861 110331 431927 110334
rect 213913 109306 213979 109309
rect 217182 109306 217242 109548
rect 230657 109442 230723 109445
rect 228968 109440 230723 109442
rect 228968 109384 230662 109440
rect 230718 109384 230723 109440
rect 228968 109382 230723 109384
rect 230657 109379 230723 109382
rect 213913 109304 217242 109306
rect 213913 109248 213918 109304
rect 213974 109248 217242 109304
rect 213913 109246 217242 109248
rect 265525 109306 265591 109309
rect 268150 109306 268210 109548
rect 279926 109518 287070 109578
rect 282269 109442 282335 109445
rect 279956 109440 282335 109442
rect 279956 109384 282274 109440
rect 282330 109384 282335 109440
rect 279956 109382 282335 109384
rect 282269 109379 282335 109382
rect 265525 109304 268210 109306
rect 265525 109248 265530 109304
rect 265586 109248 268210 109304
rect 265525 109246 268210 109248
rect 213913 109243 213979 109246
rect 265525 109243 265591 109246
rect 287010 109170 287070 109518
rect 298134 109170 298140 109172
rect 287010 109110 298140 109170
rect 298134 109108 298140 109110
rect 298204 109108 298210 109172
rect 430573 109034 430639 109037
rect 428230 109032 430639 109034
rect 231761 108898 231827 108901
rect 228968 108896 231827 108898
rect 167913 108762 167979 108765
rect 164694 108760 167979 108762
rect 164694 108704 167918 108760
rect 167974 108704 167979 108760
rect 164694 108702 167979 108704
rect 167913 108699 167979 108702
rect 214005 108354 214071 108357
rect 217182 108354 217242 108868
rect 228968 108840 231766 108896
rect 231822 108840 231827 108896
rect 228968 108838 231827 108840
rect 231761 108835 231827 108838
rect 265157 108762 265223 108765
rect 268150 108762 268210 109004
rect 428230 108976 430578 109032
rect 430634 108976 430639 109032
rect 428230 108974 430639 108976
rect 428230 108868 428290 108974
rect 430573 108971 430639 108974
rect 265157 108760 268210 108762
rect 265157 108704 265162 108760
rect 265218 108704 268210 108760
rect 265157 108702 268210 108704
rect 347497 108762 347563 108765
rect 347497 108760 350060 108762
rect 347497 108704 347502 108760
rect 347558 108704 350060 108760
rect 347497 108702 350060 108704
rect 265157 108699 265223 108702
rect 347497 108699 347563 108702
rect 280153 108626 280219 108629
rect 279956 108624 280219 108626
rect 231669 108490 231735 108493
rect 228968 108488 231735 108490
rect 228968 108432 231674 108488
rect 231730 108432 231735 108488
rect 228968 108430 231735 108432
rect 231669 108427 231735 108430
rect 214005 108352 217242 108354
rect 214005 108296 214010 108352
rect 214066 108296 217242 108352
rect 214005 108294 217242 108296
rect 265985 108354 266051 108357
rect 268150 108354 268210 108596
rect 279956 108568 280158 108624
rect 280214 108568 280219 108624
rect 279956 108566 280219 108568
rect 280153 108563 280219 108566
rect 265985 108352 268210 108354
rect 265985 108296 265990 108352
rect 266046 108296 268210 108352
rect 265985 108294 268210 108296
rect 214005 108291 214071 108294
rect 265985 108291 266051 108294
rect 213913 107946 213979 107949
rect 217182 107946 217242 108188
rect 230565 107946 230631 107949
rect 213913 107944 217242 107946
rect 213913 107888 213918 107944
rect 213974 107888 217242 107944
rect 213913 107886 217242 107888
rect 228968 107944 230631 107946
rect 228968 107888 230570 107944
rect 230626 107888 230631 107944
rect 228968 107886 230631 107888
rect 213913 107883 213979 107886
rect 230565 107883 230631 107886
rect 265709 107946 265775 107949
rect 268150 107946 268210 108188
rect 436134 107946 436140 107948
rect 265709 107944 268210 107946
rect 265709 107888 265714 107944
rect 265770 107888 268210 107944
rect 265709 107886 268210 107888
rect 428230 107886 436140 107946
rect 265709 107883 265775 107886
rect 281533 107810 281599 107813
rect 279956 107808 281599 107810
rect 265709 107674 265775 107677
rect 265709 107672 267842 107674
rect 265709 107616 265714 107672
rect 265770 107616 267842 107672
rect 265709 107614 267842 107616
rect 265709 107611 265775 107614
rect 231761 107538 231827 107541
rect 228968 107536 231827 107538
rect 214005 106994 214071 106997
rect 217182 106994 217242 107508
rect 228968 107480 231766 107536
rect 231822 107480 231827 107536
rect 228968 107478 231827 107480
rect 267782 107538 267842 107614
rect 268334 107538 268394 107780
rect 279956 107752 281538 107808
rect 281594 107752 281599 107808
rect 428230 107780 428290 107886
rect 436134 107884 436140 107886
rect 436204 107884 436210 107948
rect 279956 107750 281599 107752
rect 281533 107747 281599 107750
rect 267782 107478 268394 107538
rect 231761 107475 231827 107478
rect 231669 107130 231735 107133
rect 228968 107128 231735 107130
rect 228968 107072 231674 107128
rect 231730 107072 231735 107128
rect 228968 107070 231735 107072
rect 231669 107067 231735 107070
rect 264278 107068 264284 107132
rect 264348 107130 264354 107132
rect 268150 107130 268210 107372
rect 282821 107130 282887 107133
rect 430573 107130 430639 107133
rect 264348 107070 268210 107130
rect 279956 107128 282887 107130
rect 279956 107072 282826 107128
rect 282882 107072 282887 107128
rect 279956 107070 282887 107072
rect 264348 107068 264354 107070
rect 282821 107067 282887 107070
rect 428230 107128 430639 107130
rect 428230 107072 430578 107128
rect 430634 107072 430639 107128
rect 428230 107070 430639 107072
rect 214005 106992 217242 106994
rect 214005 106936 214010 106992
rect 214066 106936 217242 106992
rect 347497 106994 347563 106997
rect 347497 106992 350060 106994
rect 214005 106934 217242 106936
rect 214005 106931 214071 106934
rect 213913 106586 213979 106589
rect 217182 106586 217242 106828
rect 265525 106722 265591 106725
rect 268150 106722 268210 106964
rect 347497 106936 347502 106992
rect 347558 106936 350060 106992
rect 347497 106934 350060 106936
rect 347497 106931 347563 106934
rect 265525 106720 268210 106722
rect 265525 106664 265530 106720
rect 265586 106664 268210 106720
rect 428230 106692 428290 107070
rect 430573 107067 430639 107070
rect 265525 106662 268210 106664
rect 265525 106659 265591 106662
rect 231761 106586 231827 106589
rect 213913 106584 217242 106586
rect 213913 106528 213918 106584
rect 213974 106528 217242 106584
rect 213913 106526 217242 106528
rect 228968 106584 231827 106586
rect 228968 106528 231766 106584
rect 231822 106528 231827 106584
rect 228968 106526 231827 106528
rect 213913 106523 213979 106526
rect 231761 106523 231827 106526
rect 265709 106586 265775 106589
rect 265709 106584 268210 106586
rect 265709 106528 265714 106584
rect 265770 106528 268210 106584
rect 265709 106526 268210 106528
rect 265709 106523 265775 106526
rect 268150 106420 268210 106526
rect 284334 106314 284340 106316
rect 279956 106254 284340 106314
rect 284334 106252 284340 106254
rect 284404 106252 284410 106316
rect 231761 106178 231827 106181
rect 228968 106176 231827 106178
rect 213453 105770 213519 105773
rect 217182 105770 217242 106148
rect 228968 106120 231766 106176
rect 231822 106120 231827 106176
rect 228968 106118 231827 106120
rect 231761 106115 231827 106118
rect 213453 105768 217242 105770
rect 213453 105712 213458 105768
rect 213514 105712 217242 105768
rect 213453 105710 217242 105712
rect 265525 105770 265591 105773
rect 268150 105770 268210 106012
rect 430573 105906 430639 105909
rect 265525 105768 268210 105770
rect 265525 105712 265530 105768
rect 265586 105712 268210 105768
rect 265525 105710 268210 105712
rect 428230 105904 430639 105906
rect 428230 105848 430578 105904
rect 430634 105848 430639 105904
rect 428230 105846 430639 105848
rect 213453 105707 213519 105710
rect 265525 105707 265591 105710
rect 233734 105634 233740 105636
rect 214005 105362 214071 105365
rect 217182 105362 217242 105604
rect 228968 105574 233740 105634
rect 233734 105572 233740 105574
rect 233804 105572 233810 105636
rect 214005 105360 217242 105362
rect 214005 105304 214010 105360
rect 214066 105304 217242 105360
rect 214005 105302 217242 105304
rect 265709 105362 265775 105365
rect 268150 105362 268210 105604
rect 428230 105468 428290 105846
rect 430573 105843 430639 105846
rect 265709 105360 268210 105362
rect 265709 105304 265714 105360
rect 265770 105304 268210 105360
rect 265709 105302 268210 105304
rect 214005 105299 214071 105302
rect 265709 105299 265775 105302
rect 231669 105226 231735 105229
rect 228968 105224 231735 105226
rect 228968 105168 231674 105224
rect 231730 105168 231735 105224
rect 228968 105166 231735 105168
rect 231669 105163 231735 105166
rect 213913 105090 213979 105093
rect 213913 105088 217242 105090
rect 213913 105032 213918 105088
rect 213974 105032 217242 105088
rect 213913 105030 217242 105032
rect 213913 105027 213979 105030
rect 217182 104924 217242 105030
rect 265985 104954 266051 104957
rect 268334 104954 268394 105196
rect 265985 104952 268394 104954
rect 265985 104896 265990 104952
rect 266046 104896 268394 104952
rect 265985 104894 268394 104896
rect 279926 104954 279986 105468
rect 287094 104954 287100 104956
rect 279926 104894 287100 104954
rect 265985 104891 266051 104894
rect 287094 104892 287100 104894
rect 287164 104892 287170 104956
rect 304206 104892 304212 104956
rect 304276 104954 304282 104956
rect 350030 104954 350090 105332
rect 304276 104894 350090 104954
rect 304276 104892 304282 104894
rect 280337 104818 280403 104821
rect 279956 104816 280403 104818
rect 231669 104682 231735 104685
rect 228968 104680 231735 104682
rect 228968 104624 231674 104680
rect 231730 104624 231735 104680
rect 228968 104622 231735 104624
rect 231669 104619 231735 104622
rect 264513 104546 264579 104549
rect 268150 104546 268210 104788
rect 279956 104760 280342 104816
rect 280398 104760 280403 104816
rect 279956 104758 280403 104760
rect 280337 104755 280403 104758
rect 430573 104682 430639 104685
rect 264513 104544 268210 104546
rect 264513 104488 264518 104544
rect 264574 104488 268210 104544
rect 264513 104486 268210 104488
rect 428230 104680 430639 104682
rect 428230 104624 430578 104680
rect 430634 104624 430639 104680
rect 428230 104622 430639 104624
rect 264513 104483 264579 104486
rect 428230 104380 428290 104622
rect 430573 104619 430639 104622
rect 231761 104274 231827 104277
rect 228968 104272 231827 104274
rect 214005 104002 214071 104005
rect 217182 104002 217242 104244
rect 228968 104216 231766 104272
rect 231822 104216 231827 104272
rect 228968 104214 231827 104216
rect 231761 104211 231827 104214
rect 265985 104138 266051 104141
rect 268150 104138 268210 104380
rect 265985 104136 268210 104138
rect 265985 104080 265990 104136
rect 266046 104080 268210 104136
rect 265985 104078 268210 104080
rect 265985 104075 266051 104078
rect 214005 104000 217242 104002
rect 214005 103944 214010 104000
rect 214066 103944 217242 104000
rect 214005 103942 217242 103944
rect 265709 104002 265775 104005
rect 281993 104002 282059 104005
rect 265709 104000 268210 104002
rect 265709 103944 265714 104000
rect 265770 103944 268210 104000
rect 265709 103942 268210 103944
rect 279956 104000 282059 104002
rect 279956 103944 281998 104000
rect 282054 103944 282059 104000
rect 279956 103942 282059 103944
rect 214005 103939 214071 103942
rect 265709 103939 265775 103942
rect 268150 103836 268210 103942
rect 281993 103939 282059 103942
rect 213913 103730 213979 103733
rect 231485 103730 231551 103733
rect 213913 103728 217242 103730
rect 213913 103672 213918 103728
rect 213974 103672 217242 103728
rect 213913 103670 217242 103672
rect 228968 103728 231551 103730
rect 228968 103672 231490 103728
rect 231546 103672 231551 103728
rect 228968 103670 231551 103672
rect 213913 103667 213979 103670
rect 217182 103564 217242 103670
rect 231485 103667 231551 103670
rect 347037 103594 347103 103597
rect 347037 103592 350060 103594
rect 347037 103536 347042 103592
rect 347098 103536 350060 103592
rect 347037 103534 350060 103536
rect 347037 103531 347103 103534
rect 430573 103458 430639 103461
rect 428230 103456 430639 103458
rect 231117 103322 231183 103325
rect 228968 103320 231183 103322
rect 228968 103264 231122 103320
rect 231178 103264 231183 103320
rect 228968 103262 231183 103264
rect 231117 103259 231183 103262
rect 266077 103186 266143 103189
rect 268150 103186 268210 103428
rect 428230 103400 430578 103456
rect 430634 103400 430639 103456
rect 428230 103398 430639 103400
rect 428230 103292 428290 103398
rect 430573 103395 430639 103398
rect 266077 103184 268210 103186
rect 266077 103128 266082 103184
rect 266138 103128 268210 103184
rect 266077 103126 268210 103128
rect 266077 103123 266143 103126
rect 213913 102642 213979 102645
rect 217182 102642 217242 102884
rect 230565 102778 230631 102781
rect 228968 102776 230631 102778
rect 228968 102720 230570 102776
rect 230626 102720 230631 102776
rect 228968 102718 230631 102720
rect 230565 102715 230631 102718
rect 265157 102778 265223 102781
rect 268150 102778 268210 103020
rect 265157 102776 268210 102778
rect 265157 102720 265162 102776
rect 265218 102720 268210 102776
rect 265157 102718 268210 102720
rect 265157 102715 265223 102718
rect 213913 102640 217242 102642
rect 213913 102584 213918 102640
rect 213974 102584 217242 102640
rect 279926 102642 279986 103156
rect 430757 102778 430823 102781
rect 428230 102776 430823 102778
rect 428230 102720 430762 102776
rect 430818 102720 430823 102776
rect 428230 102718 430823 102720
rect 287278 102642 287284 102644
rect 213913 102582 217242 102584
rect 213913 102579 213979 102582
rect 214414 102444 214420 102508
rect 214484 102506 214490 102508
rect 214484 102446 217426 102506
rect 214484 102444 214490 102446
rect 65977 102370 66043 102373
rect 68142 102370 68816 102376
rect 65977 102368 68816 102370
rect 65977 102312 65982 102368
rect 66038 102316 68816 102368
rect 66038 102312 68202 102316
rect 65977 102310 68202 102312
rect 65977 102307 66043 102310
rect 217366 102204 217426 102446
rect 230974 102370 230980 102372
rect 228968 102310 230980 102370
rect 230974 102308 230980 102310
rect 231044 102308 231050 102372
rect 265709 102370 265775 102373
rect 268518 102372 268578 102612
rect 279926 102582 287284 102642
rect 287278 102580 287284 102582
rect 287348 102580 287354 102644
rect 281533 102506 281599 102509
rect 279956 102504 281599 102506
rect 279956 102448 281538 102504
rect 281594 102448 281599 102504
rect 279956 102446 281599 102448
rect 281533 102443 281599 102446
rect 265709 102368 268210 102370
rect 265709 102312 265714 102368
rect 265770 102312 268210 102368
rect 265709 102310 268210 102312
rect 265709 102307 265775 102310
rect 268150 102204 268210 102310
rect 268510 102308 268516 102372
rect 268580 102308 268586 102372
rect 428230 102204 428290 102718
rect 430757 102715 430823 102718
rect 264605 101962 264671 101965
rect 268510 101962 268516 101964
rect 264605 101960 268516 101962
rect 264605 101904 264610 101960
rect 264666 101904 268516 101960
rect 264605 101902 268516 101904
rect 264605 101899 264671 101902
rect 268510 101900 268516 101902
rect 268580 101900 268586 101964
rect 347221 101962 347287 101965
rect 347221 101960 350060 101962
rect 347221 101904 347226 101960
rect 347282 101904 350060 101960
rect 347221 101902 350060 101904
rect 347221 101899 347287 101902
rect 231485 101826 231551 101829
rect 228968 101824 231551 101826
rect 228968 101768 231490 101824
rect 231546 101768 231551 101824
rect 228968 101766 231551 101768
rect 231485 101763 231551 101766
rect 214833 101146 214899 101149
rect 217182 101146 217242 101524
rect 231577 101418 231643 101421
rect 228968 101416 231643 101418
rect 228968 101360 231582 101416
rect 231638 101360 231643 101416
rect 228968 101358 231643 101360
rect 231577 101355 231643 101358
rect 265341 101418 265407 101421
rect 268150 101418 268210 101796
rect 282821 101690 282887 101693
rect 279956 101688 282887 101690
rect 279956 101632 282826 101688
rect 282882 101632 282887 101688
rect 279956 101630 282887 101632
rect 282821 101627 282887 101630
rect 430573 101554 430639 101557
rect 265341 101416 268210 101418
rect 265341 101360 265346 101416
rect 265402 101360 268210 101416
rect 265341 101358 268210 101360
rect 428230 101552 430639 101554
rect 428230 101496 430578 101552
rect 430634 101496 430639 101552
rect 428230 101494 430639 101496
rect 265341 101355 265407 101358
rect 214833 101144 217242 101146
rect 214833 101088 214838 101144
rect 214894 101088 217242 101144
rect 214833 101086 217242 101088
rect 214833 101083 214899 101086
rect 265709 101010 265775 101013
rect 268150 101010 268210 101252
rect 265709 101008 268210 101010
rect 213913 100874 213979 100877
rect 213913 100872 216874 100874
rect 213913 100816 213918 100872
rect 213974 100816 216874 100872
rect 213913 100814 216874 100816
rect 213913 100811 213979 100814
rect 67725 100738 67791 100741
rect 68142 100738 68816 100744
rect 67725 100736 68816 100738
rect 67725 100680 67730 100736
rect 67786 100684 68816 100736
rect 216814 100738 216874 100814
rect 217366 100738 217426 100980
rect 265709 100952 265714 101008
rect 265770 100952 268210 101008
rect 428230 100980 428290 101494
rect 430573 101491 430639 101494
rect 265709 100950 268210 100952
rect 265709 100947 265775 100950
rect 231761 100874 231827 100877
rect 228968 100872 231827 100874
rect 228968 100816 231766 100872
rect 231822 100816 231827 100872
rect 228968 100814 231827 100816
rect 231761 100811 231827 100814
rect 265525 100874 265591 100877
rect 281717 100874 281783 100877
rect 265525 100872 267842 100874
rect 265525 100816 265530 100872
rect 265586 100816 267842 100872
rect 279956 100872 281783 100874
rect 265525 100814 267842 100816
rect 265525 100811 265591 100814
rect 67786 100680 68202 100684
rect 67725 100678 68202 100680
rect 216814 100678 217426 100738
rect 67725 100675 67791 100678
rect 267782 100602 267842 100814
rect 268334 100602 268394 100844
rect 279956 100816 281722 100872
rect 281778 100816 281783 100872
rect 279956 100814 281783 100816
rect 281717 100811 281783 100814
rect 267782 100542 268394 100602
rect 231669 100466 231735 100469
rect 228968 100464 231735 100466
rect 228968 100408 231674 100464
rect 231730 100408 231735 100464
rect 228968 100406 231735 100408
rect 231669 100403 231735 100406
rect 214005 99786 214071 99789
rect 217182 99786 217242 100300
rect 265709 100194 265775 100197
rect 268150 100194 268210 100436
rect 281717 100194 281783 100197
rect 265709 100192 268210 100194
rect 265709 100136 265714 100192
rect 265770 100136 268210 100192
rect 265709 100134 268210 100136
rect 279956 100192 281783 100194
rect 279956 100136 281722 100192
rect 281778 100136 281783 100192
rect 279956 100134 281783 100136
rect 265709 100131 265775 100134
rect 281717 100131 281783 100134
rect 347497 100194 347563 100197
rect 347497 100192 350060 100194
rect 347497 100136 347502 100192
rect 347558 100136 350060 100192
rect 347497 100134 350060 100136
rect 347497 100131 347563 100134
rect 231393 99922 231459 99925
rect 228968 99920 231459 99922
rect 228968 99864 231398 99920
rect 231454 99864 231459 99920
rect 228968 99862 231459 99864
rect 231393 99859 231459 99862
rect 214005 99784 217242 99786
rect 214005 99728 214010 99784
rect 214066 99728 217242 99784
rect 214005 99726 217242 99728
rect 265985 99786 266051 99789
rect 268150 99786 268210 100028
rect 265985 99784 268210 99786
rect 265985 99728 265990 99784
rect 266046 99728 268210 99784
rect 265985 99726 268210 99728
rect 214005 99723 214071 99726
rect 265985 99723 266051 99726
rect 213913 99514 213979 99517
rect 213913 99512 216874 99514
rect 213913 99456 213918 99512
rect 213974 99456 216874 99512
rect 213913 99454 216874 99456
rect 213913 99451 213979 99454
rect 216814 99378 216874 99454
rect 217366 99378 217426 99620
rect 231761 99514 231827 99517
rect 228968 99512 231827 99514
rect 228968 99456 231766 99512
rect 231822 99456 231827 99512
rect 228968 99454 231827 99456
rect 231761 99451 231827 99454
rect 265525 99514 265591 99517
rect 265525 99512 267842 99514
rect 265525 99456 265530 99512
rect 265586 99456 267842 99512
rect 265525 99454 267842 99456
rect 265525 99451 265591 99454
rect 216814 99318 217426 99378
rect 267782 99378 267842 99454
rect 268334 99378 268394 99620
rect 428046 99381 428106 99892
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 281574 99378 281580 99380
rect 267782 99318 268394 99378
rect 279956 99318 281580 99378
rect 281574 99316 281580 99318
rect 281644 99316 281650 99380
rect 428046 99376 428155 99381
rect 428046 99320 428094 99376
rect 428150 99320 428155 99376
rect 583520 99364 584960 99454
rect 428046 99318 428155 99320
rect 428089 99315 428155 99318
rect 230013 98970 230079 98973
rect 228968 98968 230079 98970
rect 214005 98426 214071 98429
rect 217182 98426 217242 98940
rect 228968 98912 230018 98968
rect 230074 98912 230079 98968
rect 228968 98910 230079 98912
rect 230013 98907 230079 98910
rect 266077 98834 266143 98837
rect 268150 98834 268210 99212
rect 266077 98832 268210 98834
rect 266077 98776 266082 98832
rect 266138 98776 268210 98832
rect 266077 98774 268210 98776
rect 266077 98771 266143 98774
rect 231301 98562 231367 98565
rect 228968 98560 231367 98562
rect 228968 98504 231306 98560
rect 231362 98504 231367 98560
rect 228968 98502 231367 98504
rect 231301 98499 231367 98502
rect 214005 98424 217242 98426
rect 214005 98368 214010 98424
rect 214066 98368 217242 98424
rect 214005 98366 217242 98368
rect 265617 98426 265683 98429
rect 268150 98426 268210 98668
rect 265617 98424 268210 98426
rect 265617 98368 265622 98424
rect 265678 98368 268210 98424
rect 265617 98366 268210 98368
rect 214005 98363 214071 98366
rect 265617 98363 265683 98366
rect 264605 98290 264671 98293
rect 279374 98292 279434 98532
rect 264605 98288 268026 98290
rect 213913 98018 213979 98021
rect 217366 98018 217426 98260
rect 264605 98232 264610 98288
rect 264666 98232 268026 98288
rect 264605 98230 268026 98232
rect 264605 98227 264671 98230
rect 267966 98188 268026 98230
rect 268334 98188 268394 98260
rect 279366 98228 279372 98292
rect 279436 98228 279442 98292
rect 267966 98128 268394 98188
rect 230473 98018 230539 98021
rect 213913 98016 217426 98018
rect 213913 97960 213918 98016
rect 213974 97960 217426 98016
rect 213913 97958 217426 97960
rect 228968 98016 230539 98018
rect 228968 97960 230478 98016
rect 230534 97960 230539 98016
rect 228968 97958 230539 97960
rect 213913 97955 213979 97958
rect 230473 97955 230539 97958
rect 267966 97958 268210 98018
rect 261385 97882 261451 97885
rect 267966 97882 268026 97958
rect 261385 97880 268026 97882
rect 261385 97824 261390 97880
rect 261446 97824 268026 97880
rect 268150 97852 268210 97958
rect 295926 97956 295932 98020
rect 295996 98018 296002 98020
rect 350030 98018 350090 98532
rect 428230 98293 428290 98804
rect 428181 98288 428290 98293
rect 428181 98232 428186 98288
rect 428242 98232 428290 98288
rect 428181 98230 428290 98232
rect 428181 98227 428247 98230
rect 295996 97958 350090 98018
rect 295996 97956 296002 97958
rect 281901 97882 281967 97885
rect 430573 97882 430639 97885
rect 279956 97880 281967 97882
rect 261385 97822 268026 97824
rect 279956 97824 281906 97880
rect 281962 97824 281967 97880
rect 279956 97822 281967 97824
rect 261385 97819 261451 97822
rect 281901 97819 281967 97822
rect 428230 97880 430639 97882
rect 428230 97824 430578 97880
rect 430634 97824 430639 97880
rect 428230 97822 430639 97824
rect 428230 97716 428290 97822
rect 430573 97819 430639 97822
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect 230933 97610 230999 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect 228968 97608 230999 97610
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 213913 97066 213979 97069
rect 217182 97066 217242 97580
rect 228968 97552 230938 97608
rect 230994 97552 230999 97608
rect 228968 97550 230999 97552
rect 230933 97547 230999 97550
rect 267966 97550 268210 97610
rect 264605 97474 264671 97477
rect 267966 97474 268026 97550
rect 264605 97472 268026 97474
rect 264605 97416 264610 97472
rect 264666 97416 268026 97472
rect 268150 97444 268210 97550
rect 264605 97414 268026 97416
rect 264605 97411 264671 97414
rect 229134 97140 229140 97204
rect 229204 97202 229210 97204
rect 229204 97142 258090 97202
rect 229204 97140 229210 97142
rect 230473 97066 230539 97069
rect 213913 97064 217242 97066
rect 213913 97008 213918 97064
rect 213974 97008 217242 97064
rect 213913 97006 217242 97008
rect 228968 97064 230539 97066
rect 228968 97008 230478 97064
rect 230534 97008 230539 97064
rect 228968 97006 230539 97008
rect 213913 97003 213979 97006
rect 230473 97003 230539 97006
rect 214925 96658 214991 96661
rect 217182 96658 217242 96900
rect 258030 96794 258090 97142
rect 267966 97142 268210 97202
rect 265617 97066 265683 97069
rect 267966 97066 268026 97142
rect 265617 97064 268026 97066
rect 265617 97008 265622 97064
rect 265678 97008 268026 97064
rect 268150 97036 268210 97142
rect 265617 97006 268026 97008
rect 265617 97003 265683 97006
rect 258030 96734 268210 96794
rect 229134 96658 229140 96660
rect 214925 96656 217242 96658
rect 214925 96600 214930 96656
rect 214986 96600 217242 96656
rect 214925 96598 217242 96600
rect 228968 96598 229140 96658
rect 214925 96595 214991 96598
rect 229134 96596 229140 96598
rect 229204 96658 229210 96660
rect 231761 96658 231827 96661
rect 229204 96656 231827 96658
rect 229204 96600 231766 96656
rect 231822 96600 231827 96656
rect 268150 96628 268210 96734
rect 279374 96661 279434 97036
rect 347497 96930 347563 96933
rect 347497 96928 350060 96930
rect 347497 96872 347502 96928
rect 347558 96872 350060 96928
rect 347497 96870 350060 96872
rect 347497 96867 347563 96870
rect 279325 96656 279434 96661
rect 229204 96598 231827 96600
rect 229204 96596 229210 96598
rect 231761 96595 231827 96598
rect 279325 96600 279330 96656
rect 279386 96600 279434 96656
rect 279325 96598 279434 96600
rect 279325 96595 279391 96598
rect 213913 95842 213979 95845
rect 217182 95842 217242 96356
rect 213913 95840 217242 95842
rect 213913 95784 213918 95840
rect 213974 95784 217242 95840
rect 213913 95782 217242 95784
rect 213913 95779 213979 95782
rect 228774 95706 228834 96220
rect 230565 95706 230631 95709
rect 228774 95704 230631 95706
rect 228774 95648 230570 95704
rect 230626 95648 230631 95704
rect 228774 95646 230631 95648
rect 230565 95643 230631 95646
rect 265525 95706 265591 95709
rect 268150 95706 268210 96220
rect 265525 95704 268210 95706
rect 265525 95648 265530 95704
rect 265586 95648 268210 95704
rect 265525 95646 268210 95648
rect 265525 95643 265591 95646
rect 170254 95508 170260 95572
rect 170324 95570 170330 95572
rect 279374 95570 279434 96356
rect 427678 95981 427738 96628
rect 427629 95976 427738 95981
rect 427629 95920 427634 95976
rect 427690 95920 427738 95976
rect 427629 95918 427738 95920
rect 427629 95915 427695 95918
rect 170324 95510 279434 95570
rect 170324 95508 170330 95510
rect 227662 95236 227668 95300
rect 227732 95298 227738 95300
rect 228950 95298 228956 95300
rect 227732 95238 228956 95298
rect 227732 95236 227738 95238
rect 228950 95236 228956 95238
rect 229020 95236 229026 95300
rect 177246 95100 177252 95164
rect 177316 95162 177322 95164
rect 279325 95162 279391 95165
rect 177316 95160 279391 95162
rect 177316 95104 279330 95160
rect 279386 95104 279391 95160
rect 177316 95102 279391 95104
rect 177316 95100 177322 95102
rect 279325 95099 279391 95102
rect 213177 95026 213243 95029
rect 281574 95026 281580 95028
rect 213177 95024 281580 95026
rect 213177 94968 213182 95024
rect 213238 94968 281580 95024
rect 213177 94966 281580 94968
rect 213177 94963 213243 94966
rect 281574 94964 281580 94966
rect 281644 94964 281650 95028
rect 66069 94890 66135 94893
rect 205081 94890 205147 94893
rect 66069 94888 205147 94890
rect 66069 94832 66074 94888
rect 66130 94832 205086 94888
rect 205142 94832 205147 94888
rect 66069 94830 205147 94832
rect 66069 94827 66135 94830
rect 205081 94827 205147 94830
rect 93853 94756 93919 94757
rect 106641 94756 106707 94757
rect 118233 94756 118299 94757
rect 120625 94756 120691 94757
rect 93824 94692 93830 94756
rect 93894 94754 93919 94756
rect 93894 94752 93986 94754
rect 93914 94696 93986 94752
rect 93894 94694 93986 94696
rect 93894 94692 93919 94694
rect 106608 94692 106614 94756
rect 106678 94754 106707 94756
rect 106678 94752 106770 94754
rect 106702 94696 106770 94752
rect 106678 94694 106770 94696
rect 106678 94692 106707 94694
rect 118168 94692 118174 94756
rect 118238 94754 118299 94756
rect 118238 94752 118330 94754
rect 118294 94696 118330 94752
rect 118238 94694 118330 94696
rect 118238 94692 118299 94694
rect 120616 94692 120622 94756
rect 120686 94754 120692 94756
rect 120686 94694 120778 94754
rect 120686 94692 120692 94694
rect 151486 94692 151492 94756
rect 151556 94754 151562 94756
rect 151760 94754 151766 94756
rect 151556 94694 151766 94754
rect 151556 94692 151562 94694
rect 151760 94692 151766 94694
rect 151830 94692 151836 94756
rect 93853 94691 93919 94692
rect 106641 94691 106707 94692
rect 118233 94691 118299 94692
rect 120625 94691 120691 94692
rect 66161 93802 66227 93805
rect 192569 93802 192635 93805
rect 66161 93800 192635 93802
rect 66161 93744 66166 93800
rect 66222 93744 192574 93800
rect 192630 93744 192635 93800
rect 66161 93742 192635 93744
rect 66161 93739 66227 93742
rect 192569 93739 192635 93742
rect 199469 93802 199535 93805
rect 278814 93802 278820 93804
rect 199469 93800 278820 93802
rect 199469 93744 199474 93800
rect 199530 93744 278820 93800
rect 199469 93742 278820 93744
rect 199469 93739 199535 93742
rect 278814 93740 278820 93742
rect 278884 93740 278890 93804
rect 331949 93802 332015 93805
rect 390645 93802 390711 93805
rect 331949 93800 390711 93802
rect 331949 93744 331954 93800
rect 332010 93744 390650 93800
rect 390706 93744 390711 93800
rect 331949 93742 390711 93744
rect 331949 93739 332015 93742
rect 390645 93739 390711 93742
rect 114369 93668 114435 93669
rect 151721 93668 151787 93669
rect 114318 93666 114324 93668
rect 114278 93606 114324 93666
rect 114388 93664 114435 93668
rect 151670 93666 151676 93668
rect 114430 93608 114435 93664
rect 114318 93604 114324 93606
rect 114388 93604 114435 93608
rect 151630 93606 151676 93666
rect 151740 93664 151787 93668
rect 151782 93608 151787 93664
rect 151670 93604 151676 93606
rect 151740 93604 151787 93608
rect 114369 93603 114435 93604
rect 151721 93603 151787 93604
rect 113817 93532 113883 93533
rect 129457 93532 129523 93533
rect 113766 93530 113772 93532
rect 113726 93470 113772 93530
rect 113836 93528 113883 93532
rect 129406 93530 129412 93532
rect 113878 93472 113883 93528
rect 113766 93468 113772 93470
rect 113836 93468 113883 93472
rect 129366 93470 129412 93530
rect 129476 93528 129523 93532
rect 129518 93472 129523 93528
rect 129406 93468 129412 93470
rect 129476 93468 129523 93472
rect 113817 93467 113883 93468
rect 129457 93467 129523 93468
rect 103278 93196 103284 93260
rect 103348 93258 103354 93260
rect 103421 93258 103487 93261
rect 110137 93260 110203 93261
rect 110086 93258 110092 93260
rect 103348 93256 103487 93258
rect 103348 93200 103426 93256
rect 103482 93200 103487 93256
rect 103348 93198 103487 93200
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 110198 93200 110203 93256
rect 103348 93196 103354 93198
rect 103421 93195 103487 93198
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 110137 93195 110203 93196
rect 74809 92444 74875 92445
rect 84377 92444 84443 92445
rect 88977 92444 89043 92445
rect 98177 92444 98243 92445
rect 74758 92442 74764 92444
rect 74718 92382 74764 92442
rect 74828 92440 74875 92444
rect 84326 92442 84332 92444
rect 74870 92384 74875 92440
rect 74758 92380 74764 92382
rect 74828 92380 74875 92384
rect 84286 92382 84332 92442
rect 84396 92440 84443 92444
rect 88926 92442 88932 92444
rect 84438 92384 84443 92440
rect 84326 92380 84332 92382
rect 84396 92380 84443 92384
rect 88886 92382 88932 92442
rect 88996 92440 89043 92444
rect 98126 92442 98132 92444
rect 89038 92384 89043 92440
rect 88926 92380 88932 92382
rect 88996 92380 89043 92384
rect 98086 92382 98132 92442
rect 98196 92440 98243 92444
rect 98238 92384 98243 92440
rect 98126 92380 98132 92382
rect 98196 92380 98243 92384
rect 105670 92380 105676 92444
rect 105740 92442 105746 92444
rect 105905 92442 105971 92445
rect 105740 92440 105971 92442
rect 105740 92384 105910 92440
rect 105966 92384 105971 92440
rect 105740 92382 105971 92384
rect 105740 92380 105746 92382
rect 74809 92379 74875 92380
rect 84377 92379 84443 92380
rect 88977 92379 89043 92380
rect 98177 92379 98243 92380
rect 105905 92379 105971 92382
rect 111190 92380 111196 92444
rect 111260 92442 111266 92444
rect 111609 92442 111675 92445
rect 111260 92440 111675 92442
rect 111260 92384 111614 92440
rect 111670 92384 111675 92440
rect 111260 92382 111675 92384
rect 111260 92380 111266 92382
rect 111609 92379 111675 92382
rect 115422 92380 115428 92444
rect 115492 92442 115498 92444
rect 115841 92442 115907 92445
rect 115492 92440 115907 92442
rect 115492 92384 115846 92440
rect 115902 92384 115907 92440
rect 115492 92382 115907 92384
rect 115492 92380 115498 92382
rect 115841 92379 115907 92382
rect 124438 92380 124444 92444
rect 124508 92442 124514 92444
rect 124581 92442 124647 92445
rect 125961 92444 126027 92445
rect 126513 92444 126579 92445
rect 133137 92444 133203 92445
rect 136081 92444 136147 92445
rect 151537 92444 151603 92445
rect 152089 92444 152155 92445
rect 125910 92442 125916 92444
rect 124508 92440 124647 92442
rect 124508 92384 124586 92440
rect 124642 92384 124647 92440
rect 124508 92382 124647 92384
rect 125870 92382 125916 92442
rect 125980 92440 126027 92444
rect 126462 92442 126468 92444
rect 126022 92384 126027 92440
rect 124508 92380 124514 92382
rect 124581 92379 124647 92382
rect 125910 92380 125916 92382
rect 125980 92380 126027 92384
rect 126422 92382 126468 92442
rect 126532 92440 126579 92444
rect 133086 92442 133092 92444
rect 126574 92384 126579 92440
rect 126462 92380 126468 92382
rect 126532 92380 126579 92384
rect 133046 92382 133092 92442
rect 133156 92440 133203 92444
rect 136030 92442 136036 92444
rect 133198 92384 133203 92440
rect 133086 92380 133092 92382
rect 133156 92380 133203 92384
rect 135990 92382 136036 92442
rect 136100 92440 136147 92444
rect 151486 92442 151492 92444
rect 136142 92384 136147 92440
rect 136030 92380 136036 92382
rect 136100 92380 136147 92384
rect 151446 92382 151492 92442
rect 151556 92440 151603 92444
rect 152038 92442 152044 92444
rect 151598 92384 151603 92440
rect 151486 92380 151492 92382
rect 151556 92380 151603 92384
rect 151998 92382 152044 92442
rect 152108 92440 152155 92444
rect 152150 92384 152155 92440
rect 152038 92380 152044 92382
rect 152108 92380 152155 92384
rect 125961 92379 126027 92380
rect 126513 92379 126579 92380
rect 133137 92379 133203 92380
rect 136081 92379 136147 92380
rect 151537 92379 151603 92380
rect 152089 92379 152155 92380
rect 113214 92244 113220 92308
rect 113284 92306 113290 92308
rect 166533 92306 166599 92309
rect 113284 92304 166599 92306
rect 113284 92248 166538 92304
rect 166594 92248 166599 92304
rect 113284 92246 166599 92248
rect 113284 92244 113290 92246
rect 166533 92243 166599 92246
rect 119286 92108 119292 92172
rect 119356 92170 119362 92172
rect 174629 92170 174695 92173
rect 119356 92168 174695 92170
rect 119356 92112 174634 92168
rect 174690 92112 174695 92168
rect 119356 92110 174695 92112
rect 119356 92108 119362 92110
rect 174629 92107 174695 92110
rect 120206 91836 120212 91900
rect 120276 91898 120282 91900
rect 121085 91898 121151 91901
rect 120276 91896 121151 91898
rect 120276 91840 121090 91896
rect 121146 91840 121151 91896
rect 120276 91838 121151 91840
rect 120276 91836 120282 91838
rect 121085 91835 121151 91838
rect 99966 91700 99972 91764
rect 100036 91762 100042 91764
rect 100569 91762 100635 91765
rect 100036 91760 100635 91762
rect 100036 91704 100574 91760
rect 100630 91704 100635 91760
rect 100036 91702 100635 91704
rect 100036 91700 100042 91702
rect 100569 91699 100635 91702
rect 102726 91700 102732 91764
rect 102796 91762 102802 91764
rect 102869 91762 102935 91765
rect 102796 91760 102935 91762
rect 102796 91704 102874 91760
rect 102930 91704 102935 91760
rect 102796 91702 102935 91704
rect 102796 91700 102802 91702
rect 102869 91699 102935 91702
rect 114870 91564 114876 91628
rect 114940 91626 114946 91628
rect 115841 91626 115907 91629
rect 132401 91628 132467 91629
rect 132350 91626 132356 91628
rect 114940 91624 115907 91626
rect 114940 91568 115846 91624
rect 115902 91568 115907 91624
rect 114940 91566 115907 91568
rect 132310 91566 132356 91626
rect 132420 91624 132467 91628
rect 132462 91568 132467 91624
rect 114940 91564 114946 91566
rect 115841 91563 115907 91566
rect 132350 91564 132356 91566
rect 132420 91564 132467 91568
rect 132401 91563 132467 91564
rect 101949 91492 102015 91493
rect 101949 91488 101996 91492
rect 102060 91490 102066 91492
rect 101949 91432 101954 91488
rect 101949 91428 101996 91432
rect 102060 91430 102106 91490
rect 102060 91428 102066 91430
rect 101949 91427 102015 91428
rect 96654 91292 96660 91356
rect 96724 91354 96730 91356
rect 97809 91354 97875 91357
rect 96724 91352 97875 91354
rect 96724 91296 97814 91352
rect 97870 91296 97875 91352
rect 96724 91294 97875 91296
rect 96724 91292 96730 91294
rect 97809 91291 97875 91294
rect 98494 91292 98500 91356
rect 98564 91354 98570 91356
rect 99189 91354 99255 91357
rect 101857 91356 101923 91357
rect 101806 91354 101812 91356
rect 98564 91352 99255 91354
rect 98564 91296 99194 91352
rect 99250 91296 99255 91352
rect 98564 91294 99255 91296
rect 101766 91294 101812 91354
rect 101876 91352 101923 91356
rect 101918 91296 101923 91352
rect 98564 91292 98570 91294
rect 99189 91291 99255 91294
rect 101806 91292 101812 91294
rect 101876 91292 101923 91296
rect 104198 91292 104204 91356
rect 104268 91354 104274 91356
rect 104709 91354 104775 91357
rect 104268 91352 104775 91354
rect 104268 91296 104714 91352
rect 104770 91296 104775 91352
rect 104268 91294 104775 91296
rect 104268 91292 104274 91294
rect 101857 91291 101923 91292
rect 104709 91291 104775 91294
rect 107694 91292 107700 91356
rect 107764 91354 107770 91356
rect 108941 91354 109007 91357
rect 107764 91352 109007 91354
rect 107764 91296 108946 91352
rect 109002 91296 109007 91352
rect 107764 91294 109007 91296
rect 107764 91292 107770 91294
rect 108941 91291 109007 91294
rect 109166 91292 109172 91356
rect 109236 91354 109242 91356
rect 110321 91354 110387 91357
rect 109236 91352 110387 91354
rect 109236 91296 110326 91352
rect 110382 91296 110387 91352
rect 109236 91294 110387 91296
rect 109236 91292 109242 91294
rect 110321 91291 110387 91294
rect 111926 91292 111932 91356
rect 111996 91354 112002 91356
rect 113081 91354 113147 91357
rect 117129 91356 117195 91357
rect 117078 91354 117084 91356
rect 111996 91352 113147 91354
rect 111996 91296 113086 91352
rect 113142 91296 113147 91352
rect 111996 91294 113147 91296
rect 117038 91294 117084 91354
rect 117148 91352 117195 91356
rect 117190 91296 117195 91352
rect 111996 91292 112002 91294
rect 113081 91291 113147 91294
rect 117078 91292 117084 91294
rect 117148 91292 117195 91296
rect 121678 91292 121684 91356
rect 121748 91354 121754 91356
rect 122741 91354 122807 91357
rect 121748 91352 122807 91354
rect 121748 91296 122746 91352
rect 122802 91296 122807 91352
rect 121748 91294 122807 91296
rect 121748 91292 121754 91294
rect 117129 91291 117195 91292
rect 122741 91291 122807 91294
rect 123150 91292 123156 91356
rect 123220 91354 123226 91356
rect 124029 91354 124095 91357
rect 123220 91352 124095 91354
rect 123220 91296 124034 91352
rect 124090 91296 124095 91352
rect 123220 91294 124095 91296
rect 123220 91292 123226 91294
rect 124029 91291 124095 91294
rect 85849 91220 85915 91221
rect 85798 91218 85804 91220
rect 85758 91158 85804 91218
rect 85868 91216 85915 91220
rect 85910 91160 85915 91216
rect 85798 91156 85804 91158
rect 85868 91156 85915 91160
rect 86718 91156 86724 91220
rect 86788 91218 86794 91220
rect 86861 91218 86927 91221
rect 88057 91220 88123 91221
rect 88006 91218 88012 91220
rect 86788 91216 86927 91218
rect 86788 91160 86866 91216
rect 86922 91160 86927 91216
rect 86788 91158 86927 91160
rect 87966 91158 88012 91218
rect 88076 91216 88123 91220
rect 88118 91160 88123 91216
rect 86788 91156 86794 91158
rect 85849 91155 85915 91156
rect 86861 91155 86927 91158
rect 88006 91156 88012 91158
rect 88076 91156 88123 91160
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 90633 91218 90699 91221
rect 90284 91216 90699 91218
rect 90284 91160 90638 91216
rect 90694 91160 90699 91216
rect 90284 91158 90699 91160
rect 90284 91156 90290 91158
rect 88057 91155 88123 91156
rect 90633 91155 90699 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 92289 91218 92355 91221
rect 91388 91216 92355 91218
rect 91388 91160 92294 91216
rect 92350 91160 92355 91216
rect 91388 91158 92355 91160
rect 91388 91156 91394 91158
rect 92289 91155 92355 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 94998 91156 95004 91220
rect 95068 91218 95074 91220
rect 95141 91218 95207 91221
rect 95068 91216 95207 91218
rect 95068 91160 95146 91216
rect 95202 91160 95207 91216
rect 95068 91158 95207 91160
rect 95068 91156 95074 91158
rect 95141 91155 95207 91158
rect 96286 91156 96292 91220
rect 96356 91218 96362 91220
rect 96521 91218 96587 91221
rect 96356 91216 96587 91218
rect 96356 91160 96526 91216
rect 96582 91160 96587 91216
rect 96356 91158 96587 91160
rect 96356 91156 96362 91158
rect 96521 91155 96587 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97901 91218 97967 91221
rect 97276 91216 97967 91218
rect 97276 91160 97906 91216
rect 97962 91160 97967 91216
rect 97276 91158 97967 91160
rect 97276 91156 97282 91158
rect 97901 91155 97967 91158
rect 99046 91156 99052 91220
rect 99116 91218 99122 91220
rect 99281 91218 99347 91221
rect 99116 91216 99347 91218
rect 99116 91160 99286 91216
rect 99342 91160 99347 91216
rect 99116 91158 99347 91160
rect 99116 91156 99122 91158
rect 99281 91155 99347 91158
rect 100518 91156 100524 91220
rect 100588 91218 100594 91220
rect 100661 91218 100727 91221
rect 100588 91216 100727 91218
rect 100588 91160 100666 91216
rect 100722 91160 100727 91216
rect 100588 91158 100727 91160
rect 100588 91156 100594 91158
rect 100661 91155 100727 91158
rect 100886 91156 100892 91220
rect 100956 91218 100962 91220
rect 102041 91218 102107 91221
rect 100956 91216 102107 91218
rect 100956 91160 102046 91216
rect 102102 91160 102107 91216
rect 100956 91158 102107 91160
rect 100956 91156 100962 91158
rect 102041 91155 102107 91158
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104801 91218 104867 91221
rect 104636 91216 104867 91218
rect 104636 91160 104806 91216
rect 104862 91160 104867 91216
rect 104636 91158 104867 91160
rect 104636 91156 104642 91158
rect 104801 91155 104867 91158
rect 105486 91156 105492 91220
rect 105556 91218 105562 91220
rect 106089 91218 106155 91221
rect 105556 91216 106155 91218
rect 105556 91160 106094 91216
rect 106150 91160 106155 91216
rect 105556 91158 106155 91160
rect 105556 91156 105562 91158
rect 106089 91155 106155 91158
rect 106406 91156 106412 91220
rect 106476 91218 106482 91220
rect 107193 91218 107259 91221
rect 106476 91216 107259 91218
rect 106476 91160 107198 91216
rect 107254 91160 107259 91216
rect 106476 91158 107259 91160
rect 106476 91156 106482 91158
rect 107193 91155 107259 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108849 91218 108915 91221
rect 108132 91216 108915 91218
rect 108132 91160 108854 91216
rect 108910 91160 108915 91216
rect 108132 91158 108915 91160
rect 108132 91156 108138 91158
rect 108849 91155 108915 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110229 91218 110295 91221
rect 109604 91216 110295 91218
rect 109604 91160 110234 91216
rect 110290 91160 110295 91216
rect 109604 91158 110295 91160
rect 109604 91156 109610 91158
rect 110229 91155 110295 91158
rect 110638 91156 110644 91220
rect 110708 91218 110714 91220
rect 110781 91218 110847 91221
rect 110708 91216 110847 91218
rect 110708 91160 110786 91216
rect 110842 91160 110847 91216
rect 110708 91158 110847 91160
rect 110708 91156 110714 91158
rect 110781 91155 110847 91158
rect 112294 91156 112300 91220
rect 112364 91218 112370 91220
rect 112989 91218 113055 91221
rect 112364 91216 113055 91218
rect 112364 91160 112994 91216
rect 113050 91160 113055 91216
rect 112364 91158 113055 91160
rect 112364 91156 112370 91158
rect 112989 91155 113055 91158
rect 115749 91220 115815 91221
rect 115749 91216 115796 91220
rect 115860 91218 115866 91220
rect 115749 91160 115754 91216
rect 115749 91156 115796 91160
rect 115860 91158 115906 91218
rect 115860 91156 115866 91158
rect 116710 91156 116716 91220
rect 116780 91218 116786 91220
rect 117221 91218 117287 91221
rect 116780 91216 117287 91218
rect 116780 91160 117226 91216
rect 117282 91160 117287 91216
rect 116780 91158 117287 91160
rect 116780 91156 116786 91158
rect 115749 91155 115815 91156
rect 117221 91155 117287 91158
rect 117998 91156 118004 91220
rect 118068 91218 118074 91220
rect 118233 91218 118299 91221
rect 118068 91216 118299 91218
rect 118068 91160 118238 91216
rect 118294 91160 118299 91216
rect 118068 91158 118299 91160
rect 118068 91156 118074 91158
rect 118233 91155 118299 91158
rect 119654 91156 119660 91220
rect 119724 91218 119730 91220
rect 119981 91218 120047 91221
rect 119724 91216 120047 91218
rect 119724 91160 119986 91216
rect 120042 91160 120047 91216
rect 119724 91158 120047 91160
rect 119724 91156 119730 91158
rect 119981 91155 120047 91158
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122649 91218 122715 91221
rect 122833 91220 122899 91221
rect 124121 91220 124187 91221
rect 125409 91220 125475 91221
rect 122116 91216 122715 91218
rect 122116 91160 122654 91216
rect 122710 91160 122715 91216
rect 122116 91158 122715 91160
rect 122116 91156 122122 91158
rect 122649 91155 122715 91158
rect 122782 91156 122788 91220
rect 122852 91218 122899 91220
rect 124070 91218 124076 91220
rect 122852 91216 122944 91218
rect 122894 91160 122944 91216
rect 122852 91158 122944 91160
rect 124030 91158 124076 91218
rect 124140 91216 124187 91220
rect 125358 91218 125364 91220
rect 124182 91160 124187 91216
rect 122852 91156 122899 91158
rect 124070 91156 124076 91158
rect 124140 91156 124187 91160
rect 125318 91158 125364 91218
rect 125428 91216 125475 91220
rect 125470 91160 125475 91216
rect 125358 91156 125364 91158
rect 125428 91156 125475 91160
rect 126646 91156 126652 91220
rect 126716 91218 126722 91220
rect 126881 91218 126947 91221
rect 126716 91216 126947 91218
rect 126716 91160 126886 91216
rect 126942 91160 126947 91216
rect 126716 91158 126947 91160
rect 126716 91156 126722 91158
rect 122833 91155 122899 91156
rect 124121 91155 124187 91156
rect 125409 91155 125475 91156
rect 126881 91155 126947 91158
rect 127566 91156 127572 91220
rect 127636 91218 127642 91220
rect 128169 91218 128235 91221
rect 127636 91216 128235 91218
rect 127636 91160 128174 91216
rect 128230 91160 128235 91216
rect 127636 91158 128235 91160
rect 127636 91156 127642 91158
rect 128169 91155 128235 91158
rect 130694 91156 130700 91220
rect 130764 91218 130770 91220
rect 131021 91218 131087 91221
rect 130764 91216 131087 91218
rect 130764 91160 131026 91216
rect 131082 91160 131087 91216
rect 130764 91158 131087 91160
rect 130764 91156 130770 91158
rect 131021 91155 131087 91158
rect 134374 91156 134380 91220
rect 134444 91218 134450 91220
rect 135069 91218 135135 91221
rect 134444 91216 135135 91218
rect 134444 91160 135074 91216
rect 135130 91160 135135 91216
rect 134444 91158 135135 91160
rect 134444 91156 134450 91158
rect 135069 91155 135135 91158
rect 151302 91156 151308 91220
rect 151372 91218 151378 91220
rect 151629 91218 151695 91221
rect 151372 91216 151695 91218
rect 151372 91160 151634 91216
rect 151690 91160 151695 91216
rect 151372 91158 151695 91160
rect 151372 91156 151378 91158
rect 151629 91155 151695 91158
rect 67357 91082 67423 91085
rect 214414 91082 214420 91084
rect 67357 91080 214420 91082
rect 67357 91024 67362 91080
rect 67418 91024 214420 91080
rect 67357 91022 214420 91024
rect 67357 91019 67423 91022
rect 214414 91020 214420 91022
rect 214484 91020 214490 91084
rect 214557 90402 214623 90405
rect 265750 90402 265756 90404
rect 214557 90400 265756 90402
rect 214557 90344 214562 90400
rect 214618 90344 265756 90400
rect 214557 90342 265756 90344
rect 214557 90339 214623 90342
rect 265750 90340 265756 90342
rect 265820 90340 265826 90404
rect 388437 90402 388503 90405
rect 430798 90402 430804 90404
rect 388437 90400 430804 90402
rect 388437 90344 388442 90400
rect 388498 90344 430804 90400
rect 388437 90342 430804 90344
rect 388437 90339 388503 90342
rect 430798 90340 430804 90342
rect 430868 90340 430874 90404
rect 121085 89722 121151 89725
rect 168230 89722 168236 89724
rect 121085 89720 168236 89722
rect 121085 89664 121090 89720
rect 121146 89664 168236 89720
rect 121085 89662 168236 89664
rect 121085 89659 121151 89662
rect 168230 89660 168236 89662
rect 168300 89660 168306 89724
rect 110781 88226 110847 88229
rect 166390 88226 166396 88228
rect 110781 88224 166396 88226
rect 110781 88168 110786 88224
rect 110842 88168 166396 88224
rect 110781 88166 166396 88168
rect 110781 88163 110847 88166
rect 166390 88164 166396 88166
rect 166460 88164 166466 88228
rect 295374 86940 295380 87004
rect 295444 87002 295450 87004
rect 298093 87002 298159 87005
rect 295444 87000 298159 87002
rect 295444 86944 298098 87000
rect 298154 86944 298159 87000
rect 295444 86942 298159 86944
rect 295444 86940 295450 86942
rect 298093 86939 298159 86942
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 101949 85506 102015 85509
rect 169150 85506 169156 85508
rect 101949 85504 169156 85506
rect 101949 85448 101954 85504
rect 102010 85448 169156 85504
rect 101949 85446 169156 85448
rect 101949 85443 102015 85446
rect 169150 85444 169156 85446
rect 169220 85444 169226 85508
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 103421 82786 103487 82789
rect 166206 82786 166212 82788
rect 103421 82784 166212 82786
rect 103421 82728 103426 82784
rect 103482 82728 166212 82784
rect 103421 82726 166212 82728
rect 103421 82723 103487 82726
rect 166206 82724 166212 82726
rect 166276 82724 166282 82788
rect 117221 82650 117287 82653
rect 168966 82650 168972 82652
rect 117221 82648 168972 82650
rect 117221 82592 117226 82648
rect 117282 82592 168972 82648
rect 117221 82590 168972 82592
rect 117221 82587 117287 82590
rect 168966 82588 168972 82590
rect 169036 82588 169042 82652
rect 97809 81426 97875 81429
rect 170438 81426 170444 81428
rect 97809 81424 170444 81426
rect 97809 81368 97814 81424
rect 97870 81368 170444 81424
rect 97809 81366 170444 81368
rect 97809 81363 97875 81366
rect 170438 81364 170444 81366
rect 170508 81364 170514 81428
rect 104801 81290 104867 81293
rect 173014 81290 173020 81292
rect 104801 81288 173020 81290
rect 104801 81232 104806 81288
rect 104862 81232 173020 81288
rect 104801 81230 173020 81232
rect 104801 81227 104867 81230
rect 173014 81228 173020 81230
rect 173084 81228 173090 81292
rect 9673 73810 9739 73813
rect 260046 73810 260052 73812
rect 9673 73808 260052 73810
rect 9673 73752 9678 73808
rect 9734 73752 260052 73808
rect 9673 73750 260052 73752
rect 9673 73747 9739 73750
rect 260046 73748 260052 73750
rect 260116 73748 260122 73812
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect 49693 72450 49759 72453
rect 257286 72450 257292 72452
rect 49693 72448 257292 72450
rect 49693 72392 49698 72448
rect 49754 72392 257292 72448
rect 49693 72390 257292 72392
rect 49693 72387 49759 72390
rect 257286 72388 257292 72390
rect 257356 72388 257362 72452
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 182909 70274 182975 70277
rect 227662 70274 227668 70276
rect 182909 70272 227668 70274
rect 182909 70216 182914 70272
rect 182970 70216 227668 70272
rect 182909 70214 227668 70216
rect 182909 70211 182975 70214
rect 227662 70212 227668 70214
rect 227732 70212 227738 70276
rect 13 69594 79 69597
rect 182173 69594 182239 69597
rect 182909 69594 182975 69597
rect 13 69592 182975 69594
rect 13 69536 18 69592
rect 74 69536 182178 69592
rect 182234 69536 182914 69592
rect 182970 69536 182975 69592
rect 13 69534 182975 69536
rect 13 69531 79 69534
rect 182173 69531 182239 69534
rect 182909 69531 182975 69534
rect 61878 68852 61884 68916
rect 61948 68914 61954 68916
rect 332593 68914 332659 68917
rect 333237 68914 333303 68917
rect 61948 68912 333303 68914
rect 61948 68856 332598 68912
rect 332654 68856 333242 68912
rect 333298 68856 333303 68912
rect 61948 68854 333303 68856
rect 61948 68852 61954 68854
rect 332593 68851 332659 68854
rect 333237 68851 333303 68854
rect 299657 66876 299723 66877
rect 299606 66812 299612 66876
rect 299676 66874 299723 66876
rect 299676 66872 299768 66874
rect 299718 66816 299768 66872
rect 299676 66814 299768 66816
rect 299676 66812 299723 66814
rect 299657 66811 299723 66812
rect 580257 59666 580323 59669
rect 583520 59666 584960 59756
rect 580257 59664 584960 59666
rect 580257 59608 580262 59664
rect 580318 59608 584960 59664
rect 580257 59606 584960 59608
rect 580257 59603 580323 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 78673 50282 78739 50285
rect 264278 50282 264284 50284
rect 78673 50280 264284 50282
rect 78673 50224 78678 50280
rect 78734 50224 264284 50280
rect 78673 50222 264284 50224
rect 78673 50219 78739 50222
rect 264278 50220 264284 50222
rect 264348 50220 264354 50284
rect 309225 49060 309291 49061
rect 309174 48996 309180 49060
rect 309244 49058 309291 49060
rect 309244 49056 309336 49058
rect 309286 49000 309336 49056
rect 309244 48998 309336 49000
rect 309244 48996 309291 48998
rect 309225 48995 309291 48996
rect 247718 48316 247724 48380
rect 247788 48378 247794 48380
rect 248505 48378 248571 48381
rect 247788 48376 248571 48378
rect 247788 48320 248510 48376
rect 248566 48320 248571 48376
rect 247788 48318 248571 48320
rect 247788 48316 247794 48318
rect 248505 48315 248571 48318
rect 343633 47562 343699 47565
rect 434846 47562 434852 47564
rect 343633 47560 434852 47562
rect 343633 47504 343638 47560
rect 343694 47504 434852 47560
rect 343633 47502 434852 47504
rect 343633 47499 343699 47502
rect 434846 47500 434852 47502
rect 434916 47500 434922 47564
rect 242934 46276 242940 46340
rect 243004 46338 243010 46340
rect 244273 46338 244339 46341
rect 243004 46336 244339 46338
rect 243004 46280 244278 46336
rect 244334 46280 244339 46336
rect 243004 46278 244339 46280
rect 243004 46276 243010 46278
rect 244273 46275 244339 46278
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 240409 43620 240475 43621
rect 240358 43556 240364 43620
rect 240428 43618 240475 43620
rect 240428 43616 240520 43618
rect 240470 43560 240520 43616
rect 240428 43558 240520 43560
rect 240428 43556 240475 43558
rect 240409 43555 240475 43556
rect 23473 42122 23539 42125
rect 249006 42122 249012 42124
rect 23473 42120 249012 42122
rect 23473 42064 23478 42120
rect 23534 42064 249012 42120
rect 23473 42062 249012 42064
rect 23473 42059 23539 42062
rect 249006 42060 249012 42062
rect 249076 42060 249082 42124
rect 255313 39404 255379 39405
rect 255262 39340 255268 39404
rect 255332 39402 255379 39404
rect 255332 39400 255424 39402
rect 255374 39344 255424 39400
rect 255332 39342 255424 39344
rect 255332 39340 255379 39342
rect 255313 39339 255379 39340
rect 248505 37908 248571 37909
rect 248454 37844 248460 37908
rect 248524 37906 248571 37908
rect 248524 37904 248616 37906
rect 248566 37848 248616 37904
rect 248524 37846 248616 37848
rect 248524 37844 248571 37846
rect 248505 37843 248571 37844
rect 8293 36546 8359 36549
rect 262990 36546 262996 36548
rect 8293 36544 262996 36546
rect 8293 36488 8298 36544
rect 8354 36488 262996 36544
rect 8293 36486 262996 36488
rect 8293 36483 8359 36486
rect 262990 36484 262996 36486
rect 263060 36484 263066 36548
rect 241881 35188 241947 35189
rect 241830 35124 241836 35188
rect 241900 35186 241947 35188
rect 241900 35184 241992 35186
rect 241942 35128 241992 35184
rect 241900 35126 241992 35128
rect 241900 35124 241947 35126
rect 241881 35123 241947 35124
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3233 32466 3299 32469
rect -960 32464 3299 32466
rect -960 32408 3238 32464
rect 3294 32408 3299 32464
rect -960 32406 3299 32408
rect -960 32316 480 32406
rect 3233 32403 3299 32406
rect 38653 32466 38719 32469
rect 244774 32466 244780 32468
rect 38653 32464 244780 32466
rect 38653 32408 38658 32464
rect 38714 32408 244780 32464
rect 38653 32406 244780 32408
rect 38653 32403 38719 32406
rect 244774 32404 244780 32406
rect 244844 32404 244850 32468
rect 291694 31044 291700 31108
rect 291764 31106 291770 31108
rect 294137 31106 294203 31109
rect 291764 31104 294203 31106
rect 291764 31048 294142 31104
rect 294198 31048 294203 31104
rect 291764 31046 294203 31048
rect 291764 31044 291770 31046
rect 294137 31043 294203 31046
rect 42793 26890 42859 26893
rect 262806 26890 262812 26892
rect 42793 26888 262812 26890
rect 42793 26832 42798 26888
rect 42854 26832 262812 26888
rect 42793 26830 262812 26832
rect 42793 26827 42859 26830
rect 262806 26828 262812 26830
rect 262876 26828 262882 26892
rect 120073 25530 120139 25533
rect 264094 25530 264100 25532
rect 120073 25528 264100 25530
rect 120073 25472 120078 25528
rect 120134 25472 264100 25528
rect 120073 25470 264100 25472
rect 120073 25467 120139 25470
rect 264094 25468 264100 25470
rect 264164 25468 264170 25532
rect 252921 24308 252987 24309
rect 252870 24244 252876 24308
rect 252940 24306 252987 24308
rect 252940 24304 253032 24306
rect 252982 24248 253032 24304
rect 252940 24246 253032 24248
rect 252940 24244 252987 24246
rect 252921 24243 252987 24244
rect 245745 22676 245811 22677
rect 245694 22612 245700 22676
rect 245764 22674 245811 22676
rect 245764 22672 245856 22674
rect 245806 22616 245856 22672
rect 245764 22614 245856 22616
rect 245764 22612 245811 22614
rect 245745 22611 245811 22612
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 2865 17234 2931 17237
rect 228214 17234 228220 17236
rect 2865 17232 228220 17234
rect 2865 17176 2870 17232
rect 2926 17176 228220 17232
rect 2865 17174 228220 17176
rect 2865 17171 2931 17174
rect 228214 17172 228220 17174
rect 228284 17172 228290 17236
rect 248454 15540 248460 15604
rect 248524 15602 248530 15604
rect 249701 15602 249767 15605
rect 248524 15600 249767 15602
rect 248524 15544 249706 15600
rect 249762 15544 249767 15600
rect 248524 15542 249767 15544
rect 248524 15540 248530 15542
rect 249701 15539 249767 15542
rect 119889 14514 119955 14517
rect 232446 14514 232452 14516
rect 119889 14512 232452 14514
rect 119889 14456 119894 14512
rect 119950 14456 232452 14512
rect 119889 14454 232452 14456
rect 119889 14451 119955 14454
rect 232446 14452 232452 14454
rect 232516 14452 232522 14516
rect 240358 11732 240364 11796
rect 240428 11794 240434 11796
rect 241329 11794 241395 11797
rect 240428 11792 241395 11794
rect 240428 11736 241334 11792
rect 241390 11736 241395 11792
rect 240428 11734 241395 11736
rect 240428 11732 240434 11734
rect 241329 11731 241395 11734
rect 241830 11732 241836 11796
rect 241900 11794 241906 11796
rect 242801 11794 242867 11797
rect 241900 11792 242867 11794
rect 241900 11736 242806 11792
rect 242862 11736 242867 11792
rect 241900 11734 242867 11736
rect 241900 11732 241906 11734
rect 242801 11731 242867 11734
rect 242934 11732 242940 11796
rect 243004 11794 243010 11796
rect 245101 11794 245167 11797
rect 243004 11792 245167 11794
rect 243004 11736 245106 11792
rect 245162 11736 245167 11792
rect 243004 11734 245167 11736
rect 243004 11732 243010 11734
rect 245101 11731 245167 11734
rect 245694 11732 245700 11796
rect 245764 11794 245770 11796
rect 246941 11794 247007 11797
rect 245764 11792 247007 11794
rect 245764 11736 246946 11792
rect 247002 11736 247007 11792
rect 245764 11734 247007 11736
rect 245764 11732 245770 11734
rect 246941 11731 247007 11734
rect 252870 11732 252876 11796
rect 252940 11794 252946 11796
rect 253841 11794 253907 11797
rect 252940 11792 253907 11794
rect 252940 11736 253846 11792
rect 253902 11736 253907 11792
rect 252940 11734 253907 11736
rect 252940 11732 252946 11734
rect 253841 11731 253907 11734
rect 255262 11732 255268 11796
rect 255332 11794 255338 11796
rect 256325 11794 256391 11797
rect 255332 11792 256391 11794
rect 255332 11736 256330 11792
rect 256386 11736 256391 11792
rect 255332 11734 256391 11736
rect 255332 11732 255338 11734
rect 256325 11731 256391 11734
rect 309174 11732 309180 11796
rect 309244 11794 309250 11796
rect 310237 11794 310303 11797
rect 309244 11792 310303 11794
rect 309244 11736 310242 11792
rect 310298 11736 310303 11792
rect 309244 11734 310303 11736
rect 309244 11732 309250 11734
rect 310237 11731 310303 11734
rect 258441 10980 258507 10981
rect 258390 10916 258396 10980
rect 258460 10978 258507 10980
rect 258460 10976 258552 10978
rect 258502 10920 258552 10976
rect 258460 10918 258552 10920
rect 258460 10916 258507 10918
rect 258441 10915 258507 10916
rect 251265 8260 251331 8261
rect 251214 8196 251220 8260
rect 251284 8258 251331 8260
rect 251284 8256 251376 8258
rect 251326 8200 251376 8256
rect 251284 8198 251376 8200
rect 251284 8196 251331 8198
rect 306414 8196 306420 8260
rect 306484 8258 306490 8260
rect 306741 8258 306807 8261
rect 306484 8256 306807 8258
rect 306484 8200 306746 8256
rect 306802 8200 306807 8256
rect 306484 8198 306807 8200
rect 306484 8196 306490 8198
rect 251265 8195 251331 8196
rect 306741 8195 306807 8198
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 268326 3980 268332 4044
rect 268396 4042 268402 4044
rect 286593 4042 286659 4045
rect 268396 4040 286659 4042
rect 268396 3984 286598 4040
rect 286654 3984 286659 4040
rect 268396 3982 286659 3984
rect 268396 3980 268402 3982
rect 286593 3979 286659 3982
rect 250294 3844 250300 3908
rect 250364 3906 250370 3908
rect 264973 3906 265039 3909
rect 250364 3904 265039 3906
rect 250364 3848 264978 3904
rect 265034 3848 265039 3904
rect 250364 3846 265039 3848
rect 250364 3844 250370 3846
rect 264973 3843 265039 3846
rect 240501 3498 240567 3501
rect 241329 3498 241395 3501
rect 240501 3496 241395 3498
rect 240501 3440 240506 3496
rect 240562 3440 241334 3496
rect 241390 3440 241395 3496
rect 240501 3438 241395 3440
rect 240501 3435 240567 3438
rect 241329 3435 241395 3438
rect 241697 3498 241763 3501
rect 242801 3498 242867 3501
rect 241697 3496 242867 3498
rect 241697 3440 241702 3496
rect 241758 3440 242806 3496
rect 242862 3440 242867 3496
rect 241697 3438 242867 3440
rect 241697 3435 241763 3438
rect 242801 3435 242867 3438
rect 246389 3498 246455 3501
rect 246941 3498 247007 3501
rect 246389 3496 247007 3498
rect 246389 3440 246394 3496
rect 246450 3440 246946 3496
rect 247002 3440 247007 3496
rect 246389 3438 247007 3440
rect 246389 3435 246455 3438
rect 246941 3435 247007 3438
rect 247585 3498 247651 3501
rect 247718 3498 247724 3500
rect 247585 3496 247724 3498
rect 247585 3440 247590 3496
rect 247646 3440 247724 3496
rect 247585 3438 247724 3440
rect 247585 3435 247651 3438
rect 247718 3436 247724 3438
rect 247788 3436 247794 3500
rect 248781 3498 248847 3501
rect 249701 3498 249767 3501
rect 248781 3496 249767 3498
rect 248781 3440 248786 3496
rect 248842 3440 249706 3496
rect 249762 3440 249767 3496
rect 248781 3438 249767 3440
rect 248781 3435 248847 3438
rect 249701 3435 249767 3438
rect 258257 3498 258323 3501
rect 259361 3498 259427 3501
rect 258257 3496 259427 3498
rect 258257 3440 258262 3496
rect 258318 3440 259366 3496
rect 259422 3440 259427 3496
rect 258257 3438 259427 3440
rect 258257 3435 258323 3438
rect 259361 3435 259427 3438
rect 295374 3436 295380 3500
rect 295444 3498 295450 3500
rect 296069 3498 296135 3501
rect 295444 3496 296135 3498
rect 295444 3440 296074 3496
rect 296130 3440 296135 3496
rect 295444 3438 296135 3440
rect 295444 3436 295450 3438
rect 296069 3435 296135 3438
rect 299606 3436 299612 3500
rect 299676 3498 299682 3500
rect 300761 3498 300827 3501
rect 299676 3496 300827 3498
rect 299676 3440 300766 3496
rect 300822 3440 300827 3496
rect 299676 3438 300827 3440
rect 299676 3436 299682 3438
rect 300761 3435 300827 3438
rect 305545 3498 305611 3501
rect 306230 3498 306236 3500
rect 305545 3496 306236 3498
rect 305545 3440 305550 3496
rect 305606 3440 306236 3496
rect 305545 3438 306236 3440
rect 305545 3435 305611 3438
rect 306230 3436 306236 3438
rect 306300 3436 306306 3500
rect 66713 2002 66779 2005
rect 262070 2002 262076 2004
rect 66713 2000 262076 2002
rect 66713 1944 66718 2000
rect 66774 1944 262076 2000
rect 66713 1942 262076 1944
rect 66713 1939 66779 1942
rect 262070 1940 262076 1942
rect 262140 1940 262146 2004
<< via3 >>
rect 115060 702476 115124 702540
rect 436140 701660 436204 701724
rect 111564 620196 111628 620260
rect 124260 583748 124324 583812
rect 118740 582388 118804 582452
rect 123340 575996 123404 576060
rect 64644 574228 64708 574292
rect 126100 572792 126164 572796
rect 126100 572736 126150 572792
rect 126150 572736 126164 572792
rect 126100 572732 126164 572736
rect 66116 570284 66180 570348
rect 106412 564436 106476 564500
rect 107700 563076 107764 563140
rect 62988 557500 63052 557564
rect 69980 557364 70044 557428
rect 68876 553964 68940 554028
rect 111564 553964 111628 554028
rect 106044 552604 106108 552668
rect 106780 552196 106844 552260
rect 68140 548524 68204 548588
rect 61884 546620 61948 546684
rect 66668 545124 66732 545188
rect 115980 544308 116044 544372
rect 108252 542676 108316 542740
rect 115060 538052 115124 538116
rect 101996 537916 102060 537980
rect 98500 536828 98564 536892
rect 110644 531932 110708 531996
rect 57836 498748 57900 498812
rect 111748 497388 111812 497452
rect 111932 496164 111996 496228
rect 124260 496028 124324 496092
rect 118924 494668 118988 494732
rect 54892 493308 54956 493372
rect 118740 493308 118804 493372
rect 57652 492628 57716 492692
rect 100708 490588 100772 490652
rect 48084 489092 48148 489156
rect 99328 487188 99392 487252
rect 114324 487248 114388 487252
rect 114324 487192 114374 487248
rect 114374 487192 114388 487248
rect 114324 487188 114388 487192
rect 124444 485692 124508 485756
rect 70532 484604 70596 484668
rect 126100 484332 126164 484396
rect 123340 483652 123404 483716
rect 58572 482972 58636 483036
rect 106044 481476 106108 481540
rect 53604 480796 53668 480860
rect 65932 480524 65996 480588
rect 118004 479436 118068 479500
rect 61516 478484 61580 478548
rect 64644 477396 64708 477460
rect 106412 473996 106476 474060
rect 107700 471820 107764 471884
rect 66116 471548 66180 471612
rect 60596 470732 60660 470796
rect 66116 470732 66180 470796
rect 104756 468420 104820 468484
rect 59124 467876 59188 467940
rect 64460 466380 64524 466444
rect 104756 466516 104820 466580
rect 64828 466108 64892 466172
rect 110644 465700 110708 465764
rect 104020 464068 104084 464132
rect 106780 462164 106844 462228
rect 133828 461076 133892 461140
rect 64828 460804 64892 460868
rect 62988 458764 63052 458828
rect 68876 454548 68940 454612
rect 129780 454004 129844 454068
rect 57652 453928 57716 453932
rect 57652 453872 57702 453928
rect 57702 453872 57716 453928
rect 57652 453868 57716 453872
rect 69060 451964 69124 452028
rect 115980 452024 116044 452028
rect 115980 451968 115994 452024
rect 115994 451968 116044 452024
rect 115980 451964 116044 451968
rect 64828 451420 64892 451484
rect 69060 451284 69124 451348
rect 108988 451284 109052 451348
rect 62620 451148 62684 451212
rect 64828 451208 64892 451212
rect 64828 451152 64842 451208
rect 64842 451152 64892 451208
rect 64828 451148 64892 451152
rect 108988 450468 109052 450532
rect 68140 450060 68204 450124
rect 68140 448564 68204 448628
rect 61884 447340 61948 447404
rect 111932 447204 111996 447268
rect 64828 447128 64892 447132
rect 64828 447072 64842 447128
rect 64842 447072 64892 447128
rect 64828 447068 64892 447072
rect 66668 446388 66732 446452
rect 61700 445768 61764 445772
rect 61700 445712 61750 445768
rect 61750 445712 61764 445768
rect 61700 445708 61764 445712
rect 128860 445028 128924 445092
rect 66668 442988 66732 443052
rect 58572 442444 58636 442508
rect 70348 442308 70412 442372
rect 101996 441900 102060 441964
rect 120028 442172 120092 442236
rect 125732 439452 125796 439516
rect 65932 438908 65996 438972
rect 121684 438908 121748 438972
rect 111748 438636 111812 438700
rect 98500 437820 98564 437884
rect 64828 437548 64892 437612
rect 57836 437412 57900 437476
rect 69244 436460 69308 436524
rect 70348 436112 70412 436116
rect 70348 436056 70398 436112
rect 70398 436056 70412 436112
rect 70348 436052 70412 436056
rect 48084 434556 48148 434620
rect 64828 431972 64892 432036
rect 64828 431836 64892 431900
rect 69060 428436 69124 428500
rect 64828 422316 64892 422380
rect 64828 412524 64892 412588
rect 59124 406948 59188 407012
rect 64828 403004 64892 403068
rect 61516 402188 61580 402252
rect 121868 400964 121932 401028
rect 98500 400828 98564 400892
rect 64460 400344 64524 400348
rect 64460 400288 64510 400344
rect 64510 400288 64524 400344
rect 64460 400284 64524 400288
rect 104020 397972 104084 398036
rect 118740 395252 118804 395316
rect 115428 391172 115492 391236
rect 116164 389948 116228 390012
rect 118924 389812 118988 389876
rect 124260 389812 124324 389876
rect 114324 389328 114388 389332
rect 114324 389272 114338 389328
rect 114338 389272 114388 389328
rect 114324 389268 114388 389272
rect 100708 388860 100772 388924
rect 119292 388452 119356 388516
rect 53604 388316 53668 388380
rect 58572 388376 58636 388380
rect 58572 388320 58586 388376
rect 58586 388320 58636 388376
rect 58572 388316 58636 388320
rect 305500 388316 305564 388380
rect 70900 387908 70964 387972
rect 137140 387908 137204 387972
rect 55076 387772 55140 387836
rect 117268 387696 117332 387700
rect 117268 387640 117318 387696
rect 117318 387640 117332 387696
rect 117268 387636 117332 387640
rect 50844 387092 50908 387156
rect 295380 386956 295444 387020
rect 54892 386608 54956 386612
rect 54892 386552 54942 386608
rect 54942 386552 54956 386608
rect 54892 386548 54956 386552
rect 306420 386412 306484 386476
rect 115612 385868 115676 385932
rect 268332 385324 268396 385388
rect 123524 385188 123588 385252
rect 57836 384236 57900 384300
rect 69244 384236 69308 384300
rect 69980 383148 70044 383212
rect 64644 382196 64708 382260
rect 115612 381788 115676 381852
rect 68876 379612 68940 379676
rect 124444 379672 124508 379676
rect 124444 379616 124494 379672
rect 124494 379616 124508 379672
rect 44036 379476 44100 379540
rect 64460 379476 64524 379540
rect 124444 379612 124508 379616
rect 118004 379476 118068 379540
rect 123340 378932 123404 378996
rect 60596 377980 60660 378044
rect 61884 377980 61948 378044
rect 115428 377844 115492 377908
rect 61884 376892 61948 376956
rect 252876 375940 252940 376004
rect 117268 372676 117332 372740
rect 116164 371316 116228 371380
rect 299612 370500 299676 370564
rect 119844 368324 119908 368388
rect 119292 367644 119356 367708
rect 251220 367644 251284 367708
rect 60596 365876 60660 365940
rect 255268 360844 255332 360908
rect 62620 353364 62684 353428
rect 133828 353636 133892 353700
rect 123524 352548 123588 352612
rect 68692 347380 68756 347444
rect 61700 346972 61764 347036
rect 68692 346972 68756 347036
rect 66668 345884 66732 345948
rect 129780 342892 129844 342956
rect 115980 342348 116044 342412
rect 70532 340988 70596 341052
rect 118740 339764 118804 339828
rect 57836 339356 57900 339420
rect 121684 339356 121748 339420
rect 120028 339220 120092 339284
rect 61700 338812 61764 338876
rect 68876 338676 68940 338740
rect 60596 336092 60660 336156
rect 258396 335956 258460 336020
rect 128860 335336 128924 335340
rect 128860 335280 128874 335336
rect 128874 335280 128924 335336
rect 128860 335276 128924 335280
rect 241836 334596 241900 334660
rect 59124 334052 59188 334116
rect 250300 333236 250364 333300
rect 68692 331740 68756 331804
rect 248460 331740 248524 331804
rect 245700 330380 245764 330444
rect 121868 329700 121932 329764
rect 125732 328340 125796 328404
rect 121684 323580 121748 323644
rect 121868 312564 121932 312628
rect 240364 312428 240428 312492
rect 309180 311068 309244 311132
rect 247724 309708 247788 309772
rect 64644 308348 64708 308412
rect 242940 308348 243004 308412
rect 71084 307124 71148 307188
rect 70900 306988 70964 307052
rect 252692 302228 252756 302292
rect 137140 301412 137204 301476
rect 236500 296924 236564 296988
rect 241652 296788 241716 296852
rect 123340 294204 123404 294268
rect 177252 294068 177316 294132
rect 119108 292088 119172 292092
rect 119108 292032 119122 292088
rect 119122 292032 119172 292088
rect 119108 292028 119172 292032
rect 70532 286724 70596 286788
rect 119292 286452 119356 286516
rect 285628 286452 285692 286516
rect 304212 282100 304276 282164
rect 227668 281828 227732 281892
rect 285812 280468 285876 280532
rect 58572 278972 58636 279036
rect 121868 276796 121932 276860
rect 120028 276252 120092 276316
rect 121868 276040 121932 276044
rect 121868 275984 121918 276040
rect 121918 275984 121932 276040
rect 121868 275980 121932 275984
rect 69060 273532 69124 273596
rect 298692 272444 298756 272508
rect 61700 265644 61764 265708
rect 302740 262788 302804 262852
rect 66116 260884 66180 260948
rect 123340 258708 123404 258772
rect 430620 258708 430684 258772
rect 57100 246876 57164 246940
rect 121684 243476 121748 243540
rect 427860 240756 427924 240820
rect 70532 240212 70596 240276
rect 170260 239396 170324 239460
rect 50844 238580 50908 238644
rect 59124 237220 59188 237284
rect 129780 237220 129844 237284
rect 44036 235860 44100 235924
rect 55076 235724 55140 235788
rect 124260 234500 124324 234564
rect 291884 233820 291948 233884
rect 69060 231100 69124 231164
rect 61700 226884 61764 226948
rect 287100 222804 287164 222868
rect 294460 220084 294524 220148
rect 293172 218588 293236 218652
rect 233188 216004 233252 216068
rect 287284 215868 287348 215932
rect 295932 211788 295996 211852
rect 288388 208932 288452 208996
rect 429148 206212 429212 206276
rect 57100 202132 57164 202196
rect 280292 199276 280356 199340
rect 238524 198052 238588 198116
rect 290596 197916 290660 197980
rect 66116 196556 66180 196620
rect 237420 195196 237484 195260
rect 284340 192476 284404 192540
rect 298140 189620 298204 189684
rect 349108 188260 349172 188324
rect 244228 186900 244292 186964
rect 233372 185540 233436 185604
rect 245884 182820 245948 182884
rect 70900 180100 70964 180164
rect 231900 179964 231964 180028
rect 237604 178604 237668 178668
rect 279004 178604 279068 178668
rect 228956 177788 229020 177852
rect 104572 177652 104636 177716
rect 105676 177652 105740 177716
rect 108068 177652 108132 177716
rect 116900 177712 116964 177716
rect 116900 177656 116950 177712
rect 116950 177656 116964 177712
rect 116900 177652 116964 177656
rect 119476 177712 119540 177716
rect 119476 177656 119526 177712
rect 119526 177656 119540 177712
rect 119476 177652 119540 177656
rect 121868 177652 121932 177716
rect 129412 177652 129476 177716
rect 130700 177652 130764 177716
rect 132356 177712 132420 177716
rect 132356 177656 132406 177712
rect 132406 177656 132420 177712
rect 132356 177652 132420 177656
rect 234660 177380 234724 177444
rect 288572 177380 288636 177444
rect 240548 177244 240612 177308
rect 291700 177244 291764 177308
rect 115796 177168 115860 177172
rect 115796 177112 115846 177168
rect 115846 177112 115860 177168
rect 115796 177108 115860 177112
rect 120764 177108 120828 177172
rect 133092 177168 133156 177172
rect 133092 177112 133142 177168
rect 133142 177112 133156 177168
rect 133092 177108 133156 177112
rect 97028 176972 97092 177036
rect 100708 176972 100772 177036
rect 168236 176972 168300 177036
rect 106964 176836 107028 176900
rect 101996 176760 102060 176764
rect 101996 176704 102046 176760
rect 102046 176704 102060 176760
rect 101996 176700 102060 176704
rect 109540 176700 109604 176764
rect 110644 176760 110708 176764
rect 110644 176704 110694 176760
rect 110694 176704 110708 176760
rect 110644 176700 110708 176704
rect 112116 176836 112180 176900
rect 166212 176836 166276 176900
rect 114324 176760 114388 176764
rect 114324 176704 114374 176760
rect 114374 176704 114388 176760
rect 114324 176700 114388 176704
rect 118372 176760 118436 176764
rect 118372 176704 118422 176760
rect 118422 176704 118436 176760
rect 118372 176700 118436 176704
rect 124444 176760 124508 176764
rect 124444 176704 124494 176760
rect 124494 176704 124508 176760
rect 124444 176700 124508 176704
rect 125732 176760 125796 176764
rect 125732 176704 125782 176760
rect 125782 176704 125796 176760
rect 125732 176700 125796 176704
rect 127020 176760 127084 176764
rect 127020 176704 127070 176760
rect 127070 176704 127084 176760
rect 127020 176700 127084 176704
rect 134380 176760 134444 176764
rect 134380 176704 134430 176760
rect 134430 176704 134444 176760
rect 134380 176700 134444 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 435036 176020 435100 176084
rect 135668 175536 135732 175540
rect 135668 175480 135718 175536
rect 135718 175480 135732 175536
rect 135668 175476 135732 175480
rect 98316 175400 98380 175404
rect 98316 175344 98366 175400
rect 98366 175344 98380 175400
rect 98316 175340 98380 175344
rect 128124 175400 128188 175404
rect 128124 175344 128174 175400
rect 128174 175344 128188 175400
rect 128124 175340 128188 175344
rect 158852 175400 158916 175404
rect 158852 175344 158902 175400
rect 158902 175344 158916 175400
rect 158852 175340 158916 175344
rect 229140 175204 229204 175268
rect 113142 174992 113206 174996
rect 113142 174936 113178 174992
rect 113178 174936 113206 174992
rect 113142 174932 113206 174936
rect 123070 174992 123134 174996
rect 123070 174936 123114 174992
rect 123114 174936 123134 174992
rect 123070 174932 123134 174936
rect 229140 174660 229204 174724
rect 279372 173708 279436 173772
rect 288572 171124 288636 171188
rect 434852 171124 434916 171188
rect 430804 168812 430868 168876
rect 238708 168328 238772 168332
rect 238708 168272 238758 168328
rect 238758 168272 238772 168328
rect 238708 168268 238772 168272
rect 240548 167588 240612 167652
rect 435036 165004 435100 165068
rect 237420 164732 237484 164796
rect 239260 164460 239324 164524
rect 268516 161604 268580 161668
rect 268516 161196 268580 161260
rect 166212 160108 166276 160172
rect 168236 157932 168300 157996
rect 237604 157388 237668 157452
rect 231164 154532 231228 154596
rect 233188 153308 233252 153372
rect 241652 152492 241716 152556
rect 237972 152356 238036 152420
rect 265756 150452 265820 150516
rect 234660 150044 234724 150108
rect 233372 148684 233436 148748
rect 268516 147868 268580 147932
rect 244228 147188 244292 147252
rect 233740 146916 233804 146980
rect 265756 146372 265820 146436
rect 268516 146100 268580 146164
rect 245884 144876 245948 144940
rect 230980 142700 231044 142764
rect 236500 142020 236564 142084
rect 268516 141884 268580 141948
rect 268516 140524 268580 140588
rect 252692 140116 252756 140180
rect 168236 139436 168300 139500
rect 306236 139980 306300 140044
rect 264100 139436 264164 139500
rect 168972 136852 169036 136916
rect 231900 136308 231964 136372
rect 166396 134132 166460 134196
rect 305500 134404 305564 134468
rect 173020 131140 173084 131204
rect 294460 131004 294524 131068
rect 166212 130052 166276 130116
rect 257292 130188 257356 130252
rect 430620 130732 430684 130796
rect 169156 129916 169220 129980
rect 262812 129780 262876 129844
rect 244780 128964 244844 129028
rect 265756 128964 265820 129028
rect 288388 128692 288452 128756
rect 268516 128556 268580 128620
rect 427860 128284 427924 128348
rect 268516 128148 268580 128212
rect 249012 127604 249076 127668
rect 170444 127196 170508 127260
rect 268516 127196 268580 127260
rect 268516 126788 268580 126852
rect 429148 126924 429212 126988
rect 260052 126380 260116 126444
rect 232452 125836 232516 125900
rect 239260 124748 239324 124812
rect 285628 124748 285692 124812
rect 285812 123932 285876 123996
rect 268516 122980 268580 123044
rect 298692 122708 298756 122772
rect 268516 122572 268580 122636
rect 268516 121620 268580 121684
rect 268516 121212 268580 121276
rect 291884 120124 291948 120188
rect 349108 120124 349172 120188
rect 262076 119036 262140 119100
rect 268516 117268 268580 117332
rect 231164 116996 231228 117060
rect 280292 116996 280356 117060
rect 268516 116452 268580 116516
rect 302740 113188 302804 113252
rect 262996 112644 263060 112708
rect 237972 111692 238036 111756
rect 293172 111828 293236 111892
rect 290596 110468 290660 110532
rect 298140 109108 298204 109172
rect 436140 107884 436204 107948
rect 264284 107068 264348 107132
rect 284340 106252 284404 106316
rect 233740 105572 233804 105636
rect 287100 104892 287164 104956
rect 304212 104892 304276 104956
rect 214420 102444 214484 102508
rect 230980 102308 231044 102372
rect 287284 102580 287348 102644
rect 268516 102308 268580 102372
rect 268516 101900 268580 101964
rect 281580 99316 281644 99380
rect 279372 98228 279436 98292
rect 295932 97956 295996 98020
rect 229140 97140 229204 97204
rect 229140 96596 229204 96660
rect 170260 95508 170324 95572
rect 227668 95236 227732 95300
rect 228956 95236 229020 95300
rect 177252 95100 177316 95164
rect 281580 94964 281644 95028
rect 93830 94752 93894 94756
rect 93830 94696 93858 94752
rect 93858 94696 93894 94752
rect 93830 94692 93894 94696
rect 106614 94752 106678 94756
rect 106614 94696 106646 94752
rect 106646 94696 106678 94752
rect 106614 94692 106678 94696
rect 118174 94692 118238 94756
rect 120622 94752 120686 94756
rect 120622 94696 120630 94752
rect 120630 94696 120686 94752
rect 120622 94692 120686 94696
rect 151492 94692 151556 94756
rect 151766 94692 151830 94756
rect 278820 93740 278884 93804
rect 114324 93664 114388 93668
rect 114324 93608 114374 93664
rect 114374 93608 114388 93664
rect 114324 93604 114388 93608
rect 151676 93664 151740 93668
rect 151676 93608 151726 93664
rect 151726 93608 151740 93664
rect 151676 93604 151740 93608
rect 113772 93528 113836 93532
rect 113772 93472 113822 93528
rect 113822 93472 113836 93528
rect 113772 93468 113836 93472
rect 129412 93528 129476 93532
rect 129412 93472 129462 93528
rect 129462 93472 129476 93528
rect 129412 93468 129476 93472
rect 103284 93196 103348 93260
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 74764 92440 74828 92444
rect 74764 92384 74814 92440
rect 74814 92384 74828 92440
rect 74764 92380 74828 92384
rect 84332 92440 84396 92444
rect 84332 92384 84382 92440
rect 84382 92384 84396 92440
rect 84332 92380 84396 92384
rect 88932 92440 88996 92444
rect 88932 92384 88982 92440
rect 88982 92384 88996 92440
rect 88932 92380 88996 92384
rect 98132 92440 98196 92444
rect 98132 92384 98182 92440
rect 98182 92384 98196 92440
rect 98132 92380 98196 92384
rect 105676 92380 105740 92444
rect 111196 92380 111260 92444
rect 115428 92380 115492 92444
rect 124444 92380 124508 92444
rect 125916 92440 125980 92444
rect 125916 92384 125966 92440
rect 125966 92384 125980 92440
rect 125916 92380 125980 92384
rect 126468 92440 126532 92444
rect 126468 92384 126518 92440
rect 126518 92384 126532 92440
rect 126468 92380 126532 92384
rect 133092 92440 133156 92444
rect 133092 92384 133142 92440
rect 133142 92384 133156 92440
rect 133092 92380 133156 92384
rect 136036 92440 136100 92444
rect 136036 92384 136086 92440
rect 136086 92384 136100 92440
rect 136036 92380 136100 92384
rect 151492 92440 151556 92444
rect 151492 92384 151542 92440
rect 151542 92384 151556 92440
rect 151492 92380 151556 92384
rect 152044 92440 152108 92444
rect 152044 92384 152094 92440
rect 152094 92384 152108 92440
rect 152044 92380 152108 92384
rect 113220 92244 113284 92308
rect 119292 92108 119356 92172
rect 120212 91836 120276 91900
rect 99972 91700 100036 91764
rect 102732 91700 102796 91764
rect 114876 91564 114940 91628
rect 132356 91624 132420 91628
rect 132356 91568 132406 91624
rect 132406 91568 132420 91624
rect 132356 91564 132420 91568
rect 101996 91488 102060 91492
rect 101996 91432 102010 91488
rect 102010 91432 102060 91488
rect 101996 91428 102060 91432
rect 96660 91292 96724 91356
rect 98500 91292 98564 91356
rect 101812 91352 101876 91356
rect 101812 91296 101862 91352
rect 101862 91296 101876 91352
rect 101812 91292 101876 91296
rect 104204 91292 104268 91356
rect 107700 91292 107764 91356
rect 109172 91292 109236 91356
rect 111932 91292 111996 91356
rect 117084 91352 117148 91356
rect 117084 91296 117134 91352
rect 117134 91296 117148 91352
rect 117084 91292 117148 91296
rect 121684 91292 121748 91356
rect 123156 91292 123220 91356
rect 85804 91216 85868 91220
rect 85804 91160 85854 91216
rect 85854 91160 85868 91216
rect 85804 91156 85868 91160
rect 86724 91156 86788 91220
rect 88012 91216 88076 91220
rect 88012 91160 88062 91216
rect 88062 91160 88076 91216
rect 88012 91156 88076 91160
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 95004 91156 95068 91220
rect 96292 91156 96356 91220
rect 97212 91156 97276 91220
rect 99052 91156 99116 91220
rect 100524 91156 100588 91220
rect 100892 91156 100956 91220
rect 104572 91156 104636 91220
rect 105492 91156 105556 91220
rect 106412 91156 106476 91220
rect 108068 91156 108132 91220
rect 109540 91156 109604 91220
rect 110644 91156 110708 91220
rect 112300 91156 112364 91220
rect 115796 91216 115860 91220
rect 115796 91160 115810 91216
rect 115810 91160 115860 91216
rect 115796 91156 115860 91160
rect 116716 91156 116780 91220
rect 118004 91156 118068 91220
rect 119660 91156 119724 91220
rect 122052 91156 122116 91220
rect 122788 91216 122852 91220
rect 122788 91160 122838 91216
rect 122838 91160 122852 91216
rect 122788 91156 122852 91160
rect 124076 91216 124140 91220
rect 124076 91160 124126 91216
rect 124126 91160 124140 91216
rect 124076 91156 124140 91160
rect 125364 91216 125428 91220
rect 125364 91160 125414 91216
rect 125414 91160 125428 91216
rect 125364 91156 125428 91160
rect 126652 91156 126716 91220
rect 127572 91156 127636 91220
rect 130700 91156 130764 91220
rect 134380 91156 134444 91220
rect 151308 91156 151372 91220
rect 214420 91020 214484 91084
rect 265756 90340 265820 90404
rect 430804 90340 430868 90404
rect 168236 89660 168300 89724
rect 166396 88164 166460 88228
rect 295380 86940 295444 87004
rect 169156 85444 169220 85508
rect 166212 82724 166276 82788
rect 168972 82588 169036 82652
rect 170444 81364 170508 81428
rect 173020 81228 173084 81292
rect 260052 73748 260116 73812
rect 257292 72388 257356 72452
rect 227668 70212 227732 70276
rect 61884 68852 61948 68916
rect 299612 66872 299676 66876
rect 299612 66816 299662 66872
rect 299662 66816 299676 66872
rect 299612 66812 299676 66816
rect 264284 50220 264348 50284
rect 309180 49056 309244 49060
rect 309180 49000 309230 49056
rect 309230 49000 309244 49056
rect 309180 48996 309244 49000
rect 247724 48316 247788 48380
rect 434852 47500 434916 47564
rect 242940 46276 243004 46340
rect 240364 43616 240428 43620
rect 240364 43560 240414 43616
rect 240414 43560 240428 43616
rect 240364 43556 240428 43560
rect 249012 42060 249076 42124
rect 255268 39400 255332 39404
rect 255268 39344 255318 39400
rect 255318 39344 255332 39400
rect 255268 39340 255332 39344
rect 248460 37904 248524 37908
rect 248460 37848 248510 37904
rect 248510 37848 248524 37904
rect 248460 37844 248524 37848
rect 262996 36484 263060 36548
rect 241836 35184 241900 35188
rect 241836 35128 241886 35184
rect 241886 35128 241900 35184
rect 241836 35124 241900 35128
rect 244780 32404 244844 32468
rect 291700 31044 291764 31108
rect 262812 26828 262876 26892
rect 264100 25468 264164 25532
rect 252876 24304 252940 24308
rect 252876 24248 252926 24304
rect 252926 24248 252940 24304
rect 252876 24244 252940 24248
rect 245700 22672 245764 22676
rect 245700 22616 245750 22672
rect 245750 22616 245764 22672
rect 245700 22612 245764 22616
rect 228220 17172 228284 17236
rect 248460 15540 248524 15604
rect 232452 14452 232516 14516
rect 240364 11732 240428 11796
rect 241836 11732 241900 11796
rect 242940 11732 243004 11796
rect 245700 11732 245764 11796
rect 252876 11732 252940 11796
rect 255268 11732 255332 11796
rect 309180 11732 309244 11796
rect 258396 10976 258460 10980
rect 258396 10920 258446 10976
rect 258446 10920 258460 10976
rect 258396 10916 258460 10920
rect 251220 8256 251284 8260
rect 251220 8200 251270 8256
rect 251270 8200 251284 8256
rect 251220 8196 251284 8200
rect 306420 8196 306484 8260
rect 268332 3980 268396 4044
rect 250300 3844 250364 3908
rect 247724 3436 247788 3500
rect 295380 3436 295444 3500
rect 299612 3436 299676 3500
rect 306236 3436 306300 3500
rect 262076 1940 262140 2004
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48083 489156 48149 489157
rect 48083 489092 48084 489156
rect 48148 489092 48149 489156
rect 48083 489091 48149 489092
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 48086 434621 48146 489091
rect 48954 482614 49574 518058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 54891 493372 54957 493373
rect 54891 493308 54892 493372
rect 54956 493308 54957 493372
rect 54891 493307 54957 493308
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 53603 480860 53669 480861
rect 53603 480796 53604 480860
rect 53668 480796 53669 480860
rect 53603 480795 53669 480796
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48083 434620 48149 434621
rect 48083 434556 48084 434620
rect 48148 434556 48149 434620
rect 48083 434555 48149 434556
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 44035 379540 44101 379541
rect 44035 379476 44036 379540
rect 44100 379476 44101 379540
rect 44035 379475 44101 379476
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 44038 235925 44098 379475
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 44035 235924 44101 235925
rect 44035 235860 44036 235924
rect 44100 235860 44101 235924
rect 44035 235859 44101 235860
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 53606 388381 53666 480795
rect 53603 388380 53669 388381
rect 53603 388316 53604 388380
rect 53668 388316 53669 388380
rect 53603 388315 53669 388316
rect 50843 387156 50909 387157
rect 50843 387092 50844 387156
rect 50908 387092 50909 387156
rect 50843 387091 50909 387092
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 50846 238645 50906 387091
rect 54894 386613 54954 493307
rect 55794 489454 56414 524898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 64643 574292 64709 574293
rect 64643 574228 64644 574292
rect 64708 574228 64709 574292
rect 64643 574227 64709 574228
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 62987 557564 63053 557565
rect 62987 557500 62988 557564
rect 63052 557500 63053 557564
rect 62987 557499 63053 557500
rect 61883 546684 61949 546685
rect 61883 546620 61884 546684
rect 61948 546620 61949 546684
rect 61883 546619 61949 546620
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 57835 498812 57901 498813
rect 57835 498748 57836 498812
rect 57900 498748 57901 498812
rect 57835 498747 57901 498748
rect 57651 492692 57717 492693
rect 57651 492628 57652 492692
rect 57716 492628 57717 492692
rect 57651 492627 57717 492628
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 57654 453933 57714 492627
rect 57651 453932 57717 453933
rect 57651 453868 57652 453932
rect 57716 453868 57717 453932
rect 57651 453867 57717 453868
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 57838 437477 57898 498747
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 58571 483036 58637 483037
rect 58571 482972 58572 483036
rect 58636 482972 58637 483036
rect 58571 482971 58637 482972
rect 58574 442509 58634 482971
rect 59123 467940 59189 467941
rect 59123 467876 59124 467940
rect 59188 467876 59189 467940
rect 59123 467875 59189 467876
rect 58571 442508 58637 442509
rect 58571 442444 58572 442508
rect 58636 442444 58637 442508
rect 58571 442443 58637 442444
rect 57835 437476 57901 437477
rect 57835 437412 57836 437476
rect 57900 437412 57901 437476
rect 57835 437411 57901 437412
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55075 387836 55141 387837
rect 55075 387772 55076 387836
rect 55140 387772 55141 387836
rect 55075 387771 55141 387772
rect 54891 386612 54957 386613
rect 54891 386548 54892 386612
rect 54956 386548 54957 386612
rect 54891 386547 54957 386548
rect 50843 238644 50909 238645
rect 50843 238580 50844 238644
rect 50908 238580 50909 238644
rect 50843 238579 50909 238580
rect 55078 235789 55138 387771
rect 55794 381454 56414 416898
rect 59126 407013 59186 467875
rect 59514 457174 60134 492618
rect 61515 478548 61581 478549
rect 61515 478484 61516 478548
rect 61580 478484 61581 478548
rect 61515 478483 61581 478484
rect 60595 470796 60661 470797
rect 60595 470732 60596 470796
rect 60660 470732 60661 470796
rect 60595 470731 60661 470732
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59123 407012 59189 407013
rect 59123 406948 59124 407012
rect 59188 406948 59189 407012
rect 59123 406947 59189 406948
rect 58571 388380 58637 388381
rect 58571 388316 58572 388380
rect 58636 388316 58637 388380
rect 58571 388315 58637 388316
rect 57835 384300 57901 384301
rect 57835 384236 57836 384300
rect 57900 384236 57901 384300
rect 57835 384235 57901 384236
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 57838 339421 57898 384235
rect 57835 339420 57901 339421
rect 57835 339356 57836 339420
rect 57900 339356 57901 339420
rect 57835 339355 57901 339356
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 58574 279037 58634 388315
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 60598 378045 60658 470731
rect 61518 402253 61578 478483
rect 61886 447405 61946 546619
rect 62990 458829 63050 557499
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 64646 477461 64706 574227
rect 66954 572614 67574 608058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 584000 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 584000 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 584000 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 584000 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 584000 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 584000 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 584000 99854 604338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 584000 103574 608058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 113514 691174 114134 706202
rect 115059 702540 115125 702541
rect 115059 702476 115060 702540
rect 115124 702476 115125 702540
rect 115059 702475 115125 702476
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 111563 620260 111629 620261
rect 111563 620196 111564 620260
rect 111628 620196 111629 620260
rect 111563 620195 111629 620196
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 76576 579454 76896 579486
rect 76576 579218 76618 579454
rect 76854 579218 76896 579454
rect 76576 579134 76896 579218
rect 76576 578898 76618 579134
rect 76854 578898 76896 579134
rect 76576 578866 76896 578898
rect 87840 579454 88160 579486
rect 87840 579218 87882 579454
rect 88118 579218 88160 579454
rect 87840 579134 88160 579218
rect 87840 578898 87882 579134
rect 88118 578898 88160 579134
rect 87840 578866 88160 578898
rect 99104 579454 99424 579486
rect 99104 579218 99146 579454
rect 99382 579218 99424 579454
rect 99104 579134 99424 579218
rect 99104 578898 99146 579134
rect 99382 578898 99424 579134
rect 99104 578866 99424 578898
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66115 570348 66181 570349
rect 66115 570284 66116 570348
rect 66180 570284 66181 570348
rect 66115 570283 66181 570284
rect 65931 480588 65997 480589
rect 65931 480524 65932 480588
rect 65996 480524 65997 480588
rect 65931 480523 65997 480524
rect 64643 477460 64709 477461
rect 64643 477396 64644 477460
rect 64708 477396 64709 477460
rect 64643 477395 64709 477396
rect 64459 466444 64525 466445
rect 64459 466380 64460 466444
rect 64524 466380 64525 466444
rect 64459 466379 64525 466380
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 64462 460950 64522 466379
rect 64827 466172 64893 466173
rect 64827 466170 64828 466172
rect 64646 466110 64828 466170
rect 64646 461410 64706 466110
rect 64827 466108 64828 466110
rect 64892 466108 64893 466172
rect 64827 466107 64893 466108
rect 64646 461350 64890 461410
rect 64462 460890 64706 460950
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 62987 458828 63053 458829
rect 62987 458764 62988 458828
rect 63052 458764 63053 458828
rect 62987 458763 63053 458764
rect 62619 451212 62685 451213
rect 62619 451148 62620 451212
rect 62684 451148 62685 451212
rect 62619 451147 62685 451148
rect 61883 447404 61949 447405
rect 61883 447340 61884 447404
rect 61948 447340 61949 447404
rect 61883 447339 61949 447340
rect 61699 445772 61765 445773
rect 61699 445708 61700 445772
rect 61764 445708 61765 445772
rect 61699 445707 61765 445708
rect 61515 402252 61581 402253
rect 61515 402188 61516 402252
rect 61580 402188 61581 402252
rect 61515 402187 61581 402188
rect 60595 378044 60661 378045
rect 60595 377980 60596 378044
rect 60660 377980 60661 378044
rect 60595 377979 60661 377980
rect 60595 365940 60661 365941
rect 60595 365876 60596 365940
rect 60660 365876 60661 365940
rect 60595 365875 60661 365876
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59123 334116 59189 334117
rect 59123 334052 59124 334116
rect 59188 334052 59189 334116
rect 59123 334051 59189 334052
rect 58571 279036 58637 279037
rect 58571 278972 58572 279036
rect 58636 278972 58637 279036
rect 58571 278971 58637 278972
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 57099 246940 57165 246941
rect 57099 246876 57100 246940
rect 57164 246876 57165 246940
rect 57099 246875 57165 246876
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55075 235788 55141 235789
rect 55075 235724 55076 235788
rect 55140 235724 55141 235788
rect 55075 235723 55141 235724
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 201454 56414 236898
rect 57102 202197 57162 246875
rect 59126 237285 59186 334051
rect 59514 313174 60134 348618
rect 60598 336157 60658 365875
rect 61702 347037 61762 445707
rect 61883 378044 61949 378045
rect 61883 377980 61884 378044
rect 61948 377980 61949 378044
rect 61883 377979 61949 377980
rect 61886 376957 61946 377979
rect 61883 376956 61949 376957
rect 61883 376892 61884 376956
rect 61948 376892 61949 376956
rect 61883 376891 61949 376892
rect 61699 347036 61765 347037
rect 61699 346972 61700 347036
rect 61764 346972 61765 347036
rect 61699 346971 61765 346972
rect 61699 338876 61765 338877
rect 61699 338812 61700 338876
rect 61764 338812 61765 338876
rect 61699 338811 61765 338812
rect 60595 336156 60661 336157
rect 60595 336092 60596 336156
rect 60660 336092 60661 336156
rect 60595 336091 60661 336092
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 61702 265709 61762 338811
rect 61699 265708 61765 265709
rect 61699 265644 61700 265708
rect 61764 265644 61765 265708
rect 61699 265643 61765 265644
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59123 237284 59189 237285
rect 59123 237220 59124 237284
rect 59188 237220 59189 237284
rect 59123 237219 59189 237220
rect 59514 205174 60134 240618
rect 61702 226949 61762 265643
rect 61699 226948 61765 226949
rect 61699 226884 61700 226948
rect 61764 226884 61765 226948
rect 61699 226883 61765 226884
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 57099 202196 57165 202197
rect 57099 202132 57100 202196
rect 57164 202132 57165 202196
rect 57099 202131 57165 202132
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 61886 68917 61946 376891
rect 62622 353429 62682 451147
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 64646 422310 64706 460890
rect 64830 460869 64890 461350
rect 64827 460868 64893 460869
rect 64827 460804 64828 460868
rect 64892 460804 64893 460868
rect 64827 460803 64893 460804
rect 64827 451484 64893 451485
rect 64827 451420 64828 451484
rect 64892 451420 64893 451484
rect 64827 451419 64893 451420
rect 64830 451213 64890 451419
rect 64827 451212 64893 451213
rect 64827 451148 64828 451212
rect 64892 451148 64893 451212
rect 64827 451147 64893 451148
rect 64827 447132 64893 447133
rect 64827 447068 64828 447132
rect 64892 447068 64893 447132
rect 64827 447067 64893 447068
rect 64830 437613 64890 447067
rect 65934 438973 65994 480523
rect 66118 471613 66178 570283
rect 66667 545188 66733 545189
rect 66667 545124 66668 545188
rect 66732 545124 66733 545188
rect 66667 545123 66733 545124
rect 66115 471612 66181 471613
rect 66115 471548 66116 471612
rect 66180 471548 66181 471612
rect 66115 471547 66181 471548
rect 66118 470797 66178 471547
rect 66115 470796 66181 470797
rect 66115 470732 66116 470796
rect 66180 470732 66181 470796
rect 66115 470731 66181 470732
rect 66670 446453 66730 545123
rect 66954 536614 67574 572058
rect 106411 564500 106477 564501
rect 106411 564436 106412 564500
rect 106476 564436 106477 564500
rect 106411 564435 106477 564436
rect 82208 561454 82528 561486
rect 82208 561218 82250 561454
rect 82486 561218 82528 561454
rect 82208 561134 82528 561218
rect 82208 560898 82250 561134
rect 82486 560898 82528 561134
rect 82208 560866 82528 560898
rect 93472 561454 93792 561486
rect 93472 561218 93514 561454
rect 93750 561218 93792 561454
rect 93472 561134 93792 561218
rect 93472 560898 93514 561134
rect 93750 560898 93792 561134
rect 93472 560866 93792 560898
rect 69979 557428 70045 557429
rect 69979 557364 69980 557428
rect 70044 557364 70045 557428
rect 69979 557363 70045 557364
rect 69982 557290 70042 557363
rect 69982 557230 70410 557290
rect 68875 554028 68941 554029
rect 68875 553964 68876 554028
rect 68940 553964 68941 554028
rect 68875 553963 68941 553964
rect 68139 548588 68205 548589
rect 68139 548524 68140 548588
rect 68204 548524 68205 548588
rect 68139 548523 68205 548524
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66667 446452 66733 446453
rect 66667 446388 66668 446452
rect 66732 446388 66733 446452
rect 66667 446387 66733 446388
rect 66667 443052 66733 443053
rect 66667 442988 66668 443052
rect 66732 442988 66733 443052
rect 66667 442987 66733 442988
rect 65931 438972 65997 438973
rect 65931 438908 65932 438972
rect 65996 438908 65997 438972
rect 65931 438907 65997 438908
rect 64827 437612 64893 437613
rect 64827 437548 64828 437612
rect 64892 437548 64893 437612
rect 64827 437547 64893 437548
rect 64827 432036 64893 432037
rect 64827 431972 64828 432036
rect 64892 431972 64893 432036
rect 64827 431971 64893 431972
rect 64830 431901 64890 431971
rect 64827 431900 64893 431901
rect 64827 431836 64828 431900
rect 64892 431836 64893 431900
rect 64827 431835 64893 431836
rect 64827 422380 64893 422381
rect 64827 422316 64828 422380
rect 64892 422316 64893 422380
rect 64827 422315 64893 422316
rect 64462 422250 64706 422310
rect 64462 412650 64522 422250
rect 64830 421970 64890 422315
rect 64646 421910 64890 421970
rect 64646 413130 64706 421910
rect 64646 413070 64890 413130
rect 64462 412590 64706 412650
rect 64646 402990 64706 412590
rect 64830 412589 64890 413070
rect 64827 412588 64893 412589
rect 64827 412524 64828 412588
rect 64892 412524 64893 412588
rect 64827 412523 64893 412524
rect 64827 403068 64893 403069
rect 64827 403004 64828 403068
rect 64892 403004 64893 403068
rect 64827 403003 64893 403004
rect 64462 402930 64706 402990
rect 64830 402930 64890 403003
rect 64462 400349 64522 402930
rect 64830 402870 65074 402930
rect 65014 402250 65074 402870
rect 64646 402190 65074 402250
rect 64459 400348 64525 400349
rect 64459 400284 64460 400348
rect 64524 400284 64525 400348
rect 64459 400283 64525 400284
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 62619 353428 62685 353429
rect 62619 353364 62620 353428
rect 62684 353364 62685 353428
rect 62619 353363 62685 353364
rect 63234 352894 63854 388338
rect 64646 383670 64706 402190
rect 64462 383610 64706 383670
rect 64462 379541 64522 383610
rect 64643 382260 64709 382261
rect 64643 382196 64644 382260
rect 64708 382196 64709 382260
rect 64643 382195 64709 382196
rect 64459 379540 64525 379541
rect 64459 379476 64460 379540
rect 64524 379476 64525 379540
rect 64459 379475 64525 379476
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 64646 308413 64706 382195
rect 66670 345949 66730 442987
rect 66954 428614 67574 464058
rect 68142 450125 68202 548523
rect 68878 454613 68938 553963
rect 70350 485790 70410 557230
rect 106043 552668 106109 552669
rect 106043 552604 106044 552668
rect 106108 552604 106109 552668
rect 106043 552603 106109 552604
rect 76576 543454 76896 543486
rect 76576 543218 76618 543454
rect 76854 543218 76896 543454
rect 76576 543134 76896 543218
rect 76576 542898 76618 543134
rect 76854 542898 76896 543134
rect 76576 542866 76896 542898
rect 87840 543454 88160 543486
rect 87840 543218 87882 543454
rect 88118 543218 88160 543454
rect 87840 543134 88160 543218
rect 87840 542898 87882 543134
rect 88118 542898 88160 543134
rect 87840 542866 88160 542898
rect 99104 543454 99424 543486
rect 99104 543218 99146 543454
rect 99382 543218 99424 543454
rect 99104 543134 99424 543218
rect 99104 542898 99146 543134
rect 99382 542898 99424 543134
rect 99104 542866 99424 542898
rect 73794 507454 74414 538000
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 492000 74414 506898
rect 77514 511174 78134 538000
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 492000 78134 510618
rect 81234 514894 81854 538000
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 492000 81854 514338
rect 84954 518614 85574 538000
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 492000 85574 518058
rect 91794 525454 92414 538000
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 492000 92414 524898
rect 95514 529174 96134 538000
rect 98499 536892 98565 536893
rect 98499 536828 98500 536892
rect 98564 536828 98565 536892
rect 98499 536827 98565 536828
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 492000 96134 492618
rect 98502 487250 98562 536827
rect 99234 532894 99854 538000
rect 101995 537980 102061 537981
rect 101995 537916 101996 537980
rect 102060 537916 102061 537980
rect 101995 537915 102061 537916
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 492000 99854 496338
rect 100707 490652 100773 490653
rect 100707 490588 100708 490652
rect 100772 490588 100773 490652
rect 100707 490587 100773 490588
rect 99327 487252 99393 487253
rect 99327 487250 99328 487252
rect 98502 487190 99328 487250
rect 99327 487188 99328 487190
rect 99392 487188 99393 487252
rect 99327 487187 99393 487188
rect 70350 485730 70594 485790
rect 70534 484669 70594 485730
rect 70531 484668 70597 484669
rect 70531 484604 70532 484668
rect 70596 484604 70597 484668
rect 70531 484603 70597 484604
rect 75576 471454 75896 471486
rect 75576 471218 75618 471454
rect 75854 471218 75896 471454
rect 75576 471134 75896 471218
rect 75576 470898 75618 471134
rect 75854 470898 75896 471134
rect 75576 470866 75896 470898
rect 84840 471454 85160 471486
rect 84840 471218 84882 471454
rect 85118 471218 85160 471454
rect 84840 471134 85160 471218
rect 84840 470898 84882 471134
rect 85118 470898 85160 471134
rect 84840 470866 85160 470898
rect 94104 471454 94424 471486
rect 94104 471218 94146 471454
rect 94382 471218 94424 471454
rect 94104 471134 94424 471218
rect 94104 470898 94146 471134
rect 94382 470898 94424 471134
rect 94104 470866 94424 470898
rect 68875 454612 68941 454613
rect 68875 454548 68876 454612
rect 68940 454548 68941 454612
rect 68875 454547 68941 454548
rect 80208 453454 80528 453486
rect 80208 453218 80250 453454
rect 80486 453218 80528 453454
rect 80208 453134 80528 453218
rect 80208 452898 80250 453134
rect 80486 452898 80528 453134
rect 80208 452866 80528 452898
rect 89472 453454 89792 453486
rect 89472 453218 89514 453454
rect 89750 453218 89792 453454
rect 89472 453134 89792 453218
rect 89472 452898 89514 453134
rect 89750 452898 89792 453134
rect 89472 452866 89792 452898
rect 69059 452028 69125 452029
rect 69059 451964 69060 452028
rect 69124 451964 69125 452028
rect 69059 451963 69125 451964
rect 69062 451349 69122 451963
rect 69059 451348 69125 451349
rect 69059 451284 69060 451348
rect 69124 451284 69125 451348
rect 69059 451283 69125 451284
rect 68139 450124 68205 450125
rect 68139 450060 68140 450124
rect 68204 450060 68205 450124
rect 68139 450059 68205 450060
rect 68142 448629 68202 450059
rect 68139 448628 68205 448629
rect 68139 448564 68140 448628
rect 68204 448564 68205 448628
rect 68139 448563 68205 448564
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 69062 428501 69122 451283
rect 70347 442372 70413 442373
rect 70347 442308 70348 442372
rect 70412 442370 70413 442372
rect 70412 442310 70594 442370
rect 70412 442308 70413 442310
rect 70347 442307 70413 442308
rect 70534 437490 70594 442310
rect 70534 437430 70962 437490
rect 69243 436524 69309 436525
rect 69243 436460 69244 436524
rect 69308 436460 69309 436524
rect 69243 436459 69309 436460
rect 69059 428500 69125 428501
rect 69059 428436 69060 428500
rect 69124 428436 69125 428500
rect 69059 428435 69125 428436
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 69246 384301 69306 436459
rect 70347 436116 70413 436117
rect 70347 436052 70348 436116
rect 70412 436052 70413 436116
rect 70347 436051 70413 436052
rect 70350 389190 70410 436051
rect 70350 389130 70594 389190
rect 69243 384300 69309 384301
rect 69243 384236 69244 384300
rect 69308 384236 69309 384300
rect 69243 384235 69309 384236
rect 69979 383212 70045 383213
rect 69979 383148 69980 383212
rect 70044 383210 70045 383212
rect 70534 383210 70594 389130
rect 70902 387973 70962 437430
rect 73794 435454 74414 438000
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 388000 74414 398898
rect 77514 403174 78134 438000
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 388000 78134 402618
rect 81234 406894 81854 438000
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 388000 81854 406338
rect 84954 410614 85574 438000
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 388000 85574 410058
rect 91794 417454 92414 438000
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 388000 92414 416898
rect 95514 421174 96134 438000
rect 98499 437884 98565 437885
rect 98499 437820 98500 437884
rect 98564 437820 98565 437884
rect 98499 437819 98565 437820
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 388000 96134 420618
rect 98502 400893 98562 437819
rect 99234 424894 99854 438000
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 98499 400892 98565 400893
rect 98499 400828 98500 400892
rect 98564 400828 98565 400892
rect 98499 400827 98565 400828
rect 99234 388894 99854 424338
rect 100710 388925 100770 490587
rect 101998 441965 102058 537915
rect 102954 536614 103574 538000
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 106046 481541 106106 552603
rect 106043 481540 106109 481541
rect 106043 481476 106044 481540
rect 106108 481476 106109 481540
rect 106043 481475 106109 481476
rect 106414 474061 106474 564435
rect 107699 563140 107765 563141
rect 107699 563076 107700 563140
rect 107764 563076 107765 563140
rect 107699 563075 107765 563076
rect 106779 552260 106845 552261
rect 106779 552196 106780 552260
rect 106844 552196 106845 552260
rect 106779 552195 106845 552196
rect 106411 474060 106477 474061
rect 106411 473996 106412 474060
rect 106476 473996 106477 474060
rect 106411 473995 106477 473996
rect 104755 468484 104821 468485
rect 104755 468420 104756 468484
rect 104820 468420 104821 468484
rect 104755 468419 104821 468420
rect 104758 466581 104818 468419
rect 104755 466580 104821 466581
rect 104755 466516 104756 466580
rect 104820 466516 104821 466580
rect 104755 466515 104821 466516
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 104019 464132 104085 464133
rect 104019 464068 104020 464132
rect 104084 464068 104085 464132
rect 104019 464067 104085 464068
rect 101995 441964 102061 441965
rect 101995 441900 101996 441964
rect 102060 441900 102061 441964
rect 101995 441899 102061 441900
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 104022 398037 104082 464067
rect 106782 462229 106842 552195
rect 107702 471885 107762 563075
rect 109794 543454 110414 578898
rect 111566 554029 111626 620195
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 111563 554028 111629 554029
rect 111563 553964 111564 554028
rect 111628 553964 111629 554028
rect 111563 553963 111629 553964
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 108251 542740 108317 542741
rect 108251 542676 108252 542740
rect 108316 542676 108317 542740
rect 108251 542675 108317 542676
rect 107699 471884 107765 471885
rect 107699 471820 107700 471884
rect 107764 471820 107765 471884
rect 107699 471819 107765 471820
rect 106779 462228 106845 462229
rect 106779 462164 106780 462228
rect 106844 462164 106845 462228
rect 106779 462163 106845 462164
rect 108254 451290 108314 542675
rect 109794 507454 110414 542898
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 110643 531996 110709 531997
rect 110643 531932 110644 531996
rect 110708 531932 110709 531996
rect 110643 531931 110709 531932
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 108987 451348 109053 451349
rect 108987 451290 108988 451348
rect 108254 451284 108988 451290
rect 109052 451284 109053 451348
rect 108254 451283 109053 451284
rect 108254 451230 109050 451283
rect 108990 450533 109050 451230
rect 108987 450532 109053 450533
rect 108987 450468 108988 450532
rect 109052 450468 109053 450532
rect 108987 450467 109053 450468
rect 109794 435454 110414 470898
rect 110646 465765 110706 531931
rect 113514 511174 114134 546618
rect 115062 538117 115122 702475
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 118739 582452 118805 582453
rect 118739 582388 118740 582452
rect 118804 582388 118805 582452
rect 118739 582387 118805 582388
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 115979 544372 116045 544373
rect 115979 544308 115980 544372
rect 116044 544308 116045 544372
rect 115979 544307 116045 544308
rect 115059 538116 115125 538117
rect 115059 538052 115060 538116
rect 115124 538052 115125 538116
rect 115059 538051 115125 538052
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 111747 497452 111813 497453
rect 111747 497388 111748 497452
rect 111812 497388 111813 497452
rect 111747 497387 111813 497388
rect 110643 465764 110709 465765
rect 110643 465700 110644 465764
rect 110708 465700 110709 465764
rect 110643 465699 110709 465700
rect 111750 438701 111810 497387
rect 111931 496228 111997 496229
rect 111931 496164 111932 496228
rect 111996 496164 111997 496228
rect 111931 496163 111997 496164
rect 111934 447269 111994 496163
rect 113514 475174 114134 510618
rect 114323 487252 114389 487253
rect 114323 487188 114324 487252
rect 114388 487188 114389 487252
rect 114323 487187 114389 487188
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 111931 447268 111997 447269
rect 111931 447204 111932 447268
rect 111996 447204 111997 447268
rect 111931 447203 111997 447204
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 111747 438700 111813 438701
rect 111747 438636 111748 438700
rect 111812 438636 111813 438700
rect 111747 438635 111813 438636
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 104019 398036 104085 398037
rect 104019 397972 104020 398036
rect 104084 397972 104085 398036
rect 104019 397971 104085 397972
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 100707 388924 100773 388925
rect 100707 388860 100708 388924
rect 100772 388860 100773 388924
rect 100707 388859 100773 388860
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 388000 99854 388338
rect 102954 388000 103574 392058
rect 109794 388000 110414 398898
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 388000 114134 402618
rect 114326 389333 114386 487187
rect 115982 452029 116042 544307
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 118742 493373 118802 582387
rect 120954 554614 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 124259 583812 124325 583813
rect 124259 583748 124260 583812
rect 124324 583748 124325 583812
rect 124259 583747 124325 583748
rect 123339 576060 123405 576061
rect 123339 575996 123340 576060
rect 123404 575996 123405 576060
rect 123339 575995 123405 575996
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 118923 494732 118989 494733
rect 118923 494668 118924 494732
rect 118988 494668 118989 494732
rect 118923 494667 118989 494668
rect 118739 493372 118805 493373
rect 118739 493308 118740 493372
rect 118804 493308 118805 493372
rect 118739 493307 118805 493308
rect 118003 479500 118069 479501
rect 118003 479436 118004 479500
rect 118068 479436 118069 479500
rect 118003 479435 118069 479436
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 115979 452028 116045 452029
rect 115979 451964 115980 452028
rect 116044 451964 116045 452028
rect 115979 451963 116045 451964
rect 115427 391236 115493 391237
rect 115427 391172 115428 391236
rect 115492 391172 115493 391236
rect 115427 391171 115493 391172
rect 114323 389332 114389 389333
rect 114323 389268 114324 389332
rect 114388 389268 114389 389332
rect 114323 389267 114389 389268
rect 70899 387972 70965 387973
rect 70899 387908 70900 387972
rect 70964 387908 70965 387972
rect 70899 387907 70965 387908
rect 70044 383150 70594 383210
rect 70044 383148 70045 383150
rect 69979 383147 70045 383148
rect 89568 381454 89888 381486
rect 89568 381218 89610 381454
rect 89846 381218 89888 381454
rect 89568 381134 89888 381218
rect 89568 380898 89610 381134
rect 89846 380898 89888 381134
rect 89568 380866 89888 380898
rect 68875 379676 68941 379677
rect 68875 379612 68876 379676
rect 68940 379612 68941 379676
rect 68875 379611 68941 379612
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66667 345948 66733 345949
rect 66667 345884 66668 345948
rect 66732 345884 66733 345948
rect 66667 345883 66733 345884
rect 66954 320614 67574 356058
rect 68691 347444 68757 347445
rect 68691 347380 68692 347444
rect 68756 347380 68757 347444
rect 68691 347379 68757 347380
rect 68694 347037 68754 347379
rect 68691 347036 68757 347037
rect 68691 346972 68692 347036
rect 68756 346972 68757 347036
rect 68691 346971 68757 346972
rect 68694 331805 68754 346971
rect 68878 338741 68938 379611
rect 115430 377909 115490 391171
rect 115611 385932 115677 385933
rect 115611 385868 115612 385932
rect 115676 385868 115677 385932
rect 115611 385867 115677 385868
rect 115614 381853 115674 385867
rect 115611 381852 115677 381853
rect 115611 381788 115612 381852
rect 115676 381788 115677 381852
rect 115611 381787 115677 381788
rect 115427 377908 115493 377909
rect 115427 377844 115428 377908
rect 115492 377844 115493 377908
rect 115427 377843 115493 377844
rect 74208 363454 74528 363486
rect 74208 363218 74250 363454
rect 74486 363218 74528 363454
rect 74208 363134 74528 363218
rect 74208 362898 74250 363134
rect 74486 362898 74528 363134
rect 74208 362866 74528 362898
rect 104928 363454 105248 363486
rect 104928 363218 104970 363454
rect 105206 363218 105248 363454
rect 104928 363134 105248 363218
rect 104928 362898 104970 363134
rect 105206 362898 105248 363134
rect 104928 362866 105248 362898
rect 89568 345454 89888 345486
rect 89568 345218 89610 345454
rect 89846 345218 89888 345454
rect 89568 345134 89888 345218
rect 89568 344898 89610 345134
rect 89846 344898 89888 345134
rect 89568 344866 89888 344898
rect 115982 342413 116042 451963
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 116163 390012 116229 390013
rect 116163 389948 116164 390012
rect 116228 389948 116229 390012
rect 116163 389947 116229 389948
rect 116166 371381 116226 389947
rect 117234 388000 117854 406338
rect 117267 387700 117333 387701
rect 117267 387636 117268 387700
rect 117332 387636 117333 387700
rect 117267 387635 117333 387636
rect 117270 372741 117330 387635
rect 118006 379541 118066 479435
rect 118739 395316 118805 395317
rect 118739 395252 118740 395316
rect 118804 395252 118805 395316
rect 118739 395251 118805 395252
rect 118003 379540 118069 379541
rect 118003 379476 118004 379540
rect 118068 379476 118069 379540
rect 118003 379475 118069 379476
rect 117267 372740 117333 372741
rect 117267 372676 117268 372740
rect 117332 372676 117333 372740
rect 117267 372675 117333 372676
rect 116163 371380 116229 371381
rect 116163 371316 116164 371380
rect 116228 371316 116229 371380
rect 116163 371315 116229 371316
rect 115979 342412 116045 342413
rect 115979 342348 115980 342412
rect 116044 342348 116045 342412
rect 115979 342347 116045 342348
rect 70531 341052 70597 341053
rect 70531 340988 70532 341052
rect 70596 340988 70597 341052
rect 70531 340987 70597 340988
rect 68875 338740 68941 338741
rect 68875 338676 68876 338740
rect 68940 338676 68941 338740
rect 68875 338675 68941 338676
rect 70534 335370 70594 340987
rect 118742 339829 118802 395251
rect 118926 389877 118986 494667
rect 120954 482614 121574 518058
rect 123342 483717 123402 575995
rect 124262 496093 124322 583747
rect 126099 572796 126165 572797
rect 126099 572732 126100 572796
rect 126164 572732 126165 572796
rect 126099 572731 126165 572732
rect 124259 496092 124325 496093
rect 124259 496028 124260 496092
rect 124324 496028 124325 496092
rect 124259 496027 124325 496028
rect 124443 485756 124509 485757
rect 124443 485692 124444 485756
rect 124508 485692 124509 485756
rect 124443 485691 124509 485692
rect 123339 483716 123405 483717
rect 123339 483652 123340 483716
rect 123404 483652 123405 483716
rect 123339 483651 123405 483652
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120027 442236 120093 442237
rect 120027 442172 120028 442236
rect 120092 442172 120093 442236
rect 120027 442171 120093 442172
rect 118923 389876 118989 389877
rect 118923 389812 118924 389876
rect 118988 389812 118989 389876
rect 118923 389811 118989 389812
rect 119291 388516 119357 388517
rect 119291 388452 119292 388516
rect 119356 388452 119357 388516
rect 119291 388451 119357 388452
rect 119294 367709 119354 388451
rect 119843 368388 119909 368389
rect 119843 368324 119844 368388
rect 119908 368324 119909 368388
rect 119843 368323 119909 368324
rect 119291 367708 119357 367709
rect 119291 367644 119292 367708
rect 119356 367644 119357 367708
rect 119291 367643 119357 367644
rect 118739 339828 118805 339829
rect 118739 339764 118740 339828
rect 118804 339764 118805 339828
rect 118739 339763 118805 339764
rect 70534 335310 70962 335370
rect 68691 331804 68757 331805
rect 68691 331740 68692 331804
rect 68756 331740 68757 331804
rect 68691 331739 68757 331740
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 64643 308412 64709 308413
rect 64643 308348 64644 308412
rect 64708 308348 64709 308412
rect 64643 308347 64709 308348
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 66954 284614 67574 320058
rect 70902 307053 70962 335310
rect 73794 327454 74414 338000
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 71083 307188 71149 307189
rect 71083 307124 71084 307188
rect 71148 307124 71149 307188
rect 71083 307123 71149 307124
rect 70899 307052 70965 307053
rect 70899 306988 70900 307052
rect 70964 306988 70965 307052
rect 70899 306987 70965 306988
rect 71086 287070 71146 307123
rect 73794 294000 74414 326898
rect 77514 331174 78134 338000
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 294000 78134 294618
rect 81234 334894 81854 338000
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 294000 81854 298338
rect 84954 302614 85574 338000
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 294000 85574 302058
rect 91794 309454 92414 338000
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 95514 313174 96134 338000
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 294000 96134 312618
rect 99234 316894 99854 338000
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 294000 99854 316338
rect 102954 320614 103574 338000
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 294000 103574 320058
rect 109794 327454 110414 338000
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 113514 331174 114134 338000
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 294000 114134 294618
rect 117234 334894 117854 338000
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 294000 117854 298338
rect 119107 292092 119173 292093
rect 119107 292028 119108 292092
rect 119172 292028 119173 292092
rect 119107 292027 119173 292028
rect 70534 287010 71146 287070
rect 119110 287070 119170 292027
rect 119846 287070 119906 368323
rect 120030 339285 120090 442171
rect 120954 410614 121574 446058
rect 121683 438972 121749 438973
rect 121683 438908 121684 438972
rect 121748 438908 121749 438972
rect 121683 438907 121749 438908
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120027 339284 120093 339285
rect 120027 339220 120028 339284
rect 120092 339220 120093 339284
rect 120027 339219 120093 339220
rect 120954 338614 121574 374058
rect 121686 339421 121746 438907
rect 121867 401028 121933 401029
rect 121867 400964 121868 401028
rect 121932 400964 121933 401028
rect 121867 400963 121933 400964
rect 121683 339420 121749 339421
rect 121683 339356 121684 339420
rect 121748 339356 121749 339420
rect 121683 339355 121749 339356
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 121870 329765 121930 400963
rect 123342 378997 123402 483651
rect 124259 389876 124325 389877
rect 124259 389812 124260 389876
rect 124324 389812 124325 389876
rect 124259 389811 124325 389812
rect 123523 385252 123589 385253
rect 123523 385188 123524 385252
rect 123588 385188 123589 385252
rect 123523 385187 123589 385188
rect 123339 378996 123405 378997
rect 123339 378932 123340 378996
rect 123404 378932 123405 378996
rect 123339 378931 123405 378932
rect 123526 352613 123586 385187
rect 123523 352612 123589 352613
rect 123523 352548 123524 352612
rect 123588 352548 123589 352612
rect 123523 352547 123589 352548
rect 121867 329764 121933 329765
rect 121867 329700 121868 329764
rect 121932 329700 121933 329764
rect 121867 329699 121933 329700
rect 121683 323644 121749 323645
rect 121683 323580 121684 323644
rect 121748 323580 121749 323644
rect 121683 323579 121749 323580
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 294000 121574 302058
rect 119110 287010 119354 287070
rect 119846 287010 120090 287070
rect 70534 286789 70594 287010
rect 70531 286788 70597 286789
rect 70531 286724 70532 286788
rect 70596 286724 70597 286788
rect 70531 286723 70597 286724
rect 119294 286517 119354 287010
rect 119291 286516 119357 286517
rect 119291 286452 119292 286516
rect 119356 286452 119357 286516
rect 119291 286451 119357 286452
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66115 260948 66181 260949
rect 66115 260884 66116 260948
rect 66180 260884 66181 260948
rect 66115 260883 66181 260884
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 66118 196621 66178 260883
rect 66954 248614 67574 284058
rect 120030 276317 120090 287010
rect 120027 276316 120093 276317
rect 120027 276252 120028 276316
rect 120092 276252 120093 276316
rect 120027 276251 120093 276252
rect 69059 273596 69125 273597
rect 69059 273532 69060 273596
rect 69124 273532 69125 273596
rect 69059 273531 69125 273532
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 69062 231165 69122 273531
rect 89568 273454 89888 273486
rect 89568 273218 89610 273454
rect 89846 273218 89888 273454
rect 89568 273134 89888 273218
rect 89568 272898 89610 273134
rect 89846 272898 89888 273134
rect 89568 272866 89888 272898
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 121686 243541 121746 323579
rect 121867 312628 121933 312629
rect 121867 312564 121868 312628
rect 121932 312564 121933 312628
rect 121867 312563 121933 312564
rect 121870 276861 121930 312563
rect 123339 294268 123405 294269
rect 123339 294204 123340 294268
rect 123404 294204 123405 294268
rect 123339 294203 123405 294204
rect 121867 276860 121933 276861
rect 121867 276796 121868 276860
rect 121932 276796 121933 276860
rect 121867 276795 121933 276796
rect 121870 276045 121930 276795
rect 121867 276044 121933 276045
rect 121867 275980 121868 276044
rect 121932 275980 121933 276044
rect 121867 275979 121933 275980
rect 123342 258773 123402 294203
rect 123339 258772 123405 258773
rect 123339 258708 123340 258772
rect 123404 258708 123405 258772
rect 123339 258707 123405 258708
rect 121683 243540 121749 243541
rect 121683 243476 121684 243540
rect 121748 243476 121749 243540
rect 121683 243475 121749 243476
rect 70531 240276 70597 240277
rect 70531 240212 70532 240276
rect 70596 240212 70597 240276
rect 70531 240211 70597 240212
rect 70534 238770 70594 240211
rect 70534 238710 70962 238770
rect 69059 231164 69125 231165
rect 69059 231100 69060 231164
rect 69124 231100 69125 231164
rect 69059 231099 69125 231100
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66115 196620 66181 196621
rect 66115 196556 66116 196620
rect 66180 196556 66181 196620
rect 66115 196555 66181 196556
rect 66954 176600 67574 212058
rect 70902 180165 70962 238710
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 70899 180164 70965 180165
rect 70899 180100 70900 180164
rect 70964 180100 70965 180164
rect 70899 180099 70965 180100
rect 73794 176600 74414 182898
rect 77514 223174 78134 238000
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 238000
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 230614 85574 238000
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 238000
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 238000
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 177036 97093 177037
rect 97027 176972 97028 177036
rect 97092 176972 97093 177036
rect 97027 176971 97093 176972
rect 97030 175130 97090 176971
rect 99234 176600 99854 208338
rect 102954 212614 103574 238000
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 100707 177036 100773 177037
rect 100707 176972 100708 177036
rect 100772 176972 100773 177036
rect 100707 176971 100773 176972
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 98315 175404 98381 175405
rect 98315 175340 98316 175404
rect 98380 175340 98381 175404
rect 98315 175339 98381 175340
rect 96960 175070 97090 175130
rect 98318 175130 98378 175339
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 176971
rect 101995 176764 102061 176765
rect 101995 176700 101996 176764
rect 102060 176700 102061 176764
rect 101995 176699 102061 176700
rect 101998 175130 102058 176699
rect 102954 176600 103574 212058
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 104571 177716 104637 177717
rect 104571 177652 104572 177716
rect 104636 177652 104637 177716
rect 104571 177651 104637 177652
rect 105675 177716 105741 177717
rect 105675 177652 105676 177716
rect 105740 177652 105741 177716
rect 105675 177651 105741 177652
rect 108067 177716 108133 177717
rect 108067 177652 108068 177716
rect 108132 177652 108133 177716
rect 108067 177651 108133 177652
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 177651
rect 105678 175130 105738 177651
rect 106963 176900 107029 176901
rect 106963 176836 106964 176900
rect 107028 176836 107029 176900
rect 106963 176835 107029 176836
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 176835
rect 108070 175130 108130 177651
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109542 174994 109602 176699
rect 109794 176600 110414 182898
rect 113514 223174 114134 238000
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 112115 176900 112181 176901
rect 112115 176836 112116 176900
rect 112180 176836 112181 176900
rect 112115 176835 112181 176836
rect 110643 176764 110709 176765
rect 110643 176700 110644 176764
rect 110708 176700 110709 176764
rect 110643 176699 110709 176700
rect 110646 175130 110706 176699
rect 112118 175130 112178 176835
rect 113514 176600 114134 186618
rect 117234 226894 117854 238000
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 116899 177716 116965 177717
rect 116899 177652 116900 177716
rect 116964 177652 116965 177716
rect 116899 177651 116965 177652
rect 115795 177172 115861 177173
rect 115795 177108 115796 177172
rect 115860 177108 115861 177172
rect 115795 177107 115861 177108
rect 114323 176764 114389 176765
rect 114323 176700 114324 176764
rect 114388 176700 114389 176764
rect 114323 176699 114389 176700
rect 110646 175070 110756 175130
rect 109472 174934 109602 174994
rect 109472 174494 109532 174934
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 114326 175130 114386 176699
rect 115798 175130 115858 177107
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113141 174996 113207 174997
rect 113141 174932 113142 174996
rect 113206 174932 113207 174996
rect 113141 174931 113207 174932
rect 113144 174494 113204 174931
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 177651
rect 117234 176600 117854 190338
rect 120954 230614 121574 238000
rect 124262 234565 124322 389811
rect 124446 379677 124506 485691
rect 126102 484397 126162 572731
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 126099 484396 126165 484397
rect 126099 484332 126100 484396
rect 126164 484332 126165 484396
rect 126099 484331 126165 484332
rect 127794 453454 128414 488898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 133827 461140 133893 461141
rect 133827 461076 133828 461140
rect 133892 461076 133893 461140
rect 133827 461075 133893 461076
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 129779 454068 129845 454069
rect 129779 454004 129780 454068
rect 129844 454004 129845 454068
rect 129779 454003 129845 454004
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 125731 439516 125797 439517
rect 125731 439452 125732 439516
rect 125796 439452 125797 439516
rect 125731 439451 125797 439452
rect 124443 379676 124509 379677
rect 124443 379612 124444 379676
rect 124508 379612 124509 379676
rect 124443 379611 124509 379612
rect 125734 328405 125794 439451
rect 127794 417454 128414 452898
rect 128859 445092 128925 445093
rect 128859 445028 128860 445092
rect 128924 445028 128925 445092
rect 128859 445027 128925 445028
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 125731 328404 125797 328405
rect 125731 328340 125732 328404
rect 125796 328340 125797 328404
rect 125731 328339 125797 328340
rect 127794 309454 128414 344898
rect 128862 335341 128922 445027
rect 129782 342957 129842 454003
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 133830 353701 133890 461075
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 133827 353700 133893 353701
rect 133827 353636 133828 353700
rect 133892 353636 133893 353700
rect 133827 353635 133893 353636
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 129779 342956 129845 342957
rect 129779 342892 129780 342956
rect 129844 342892 129845 342956
rect 129779 342891 129845 342892
rect 128859 335340 128925 335341
rect 128859 335276 128860 335340
rect 128924 335276 128925 335340
rect 128859 335275 128925 335276
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 129782 237285 129842 342891
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 129779 237284 129845 237285
rect 129779 237220 129780 237284
rect 129844 237220 129845 237284
rect 129779 237219 129845 237220
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 124259 234564 124325 234565
rect 124259 234500 124260 234564
rect 124324 234500 124325 234564
rect 124259 234499 124325 234500
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 119475 177716 119541 177717
rect 119475 177652 119476 177716
rect 119540 177652 119541 177716
rect 119475 177651 119541 177652
rect 118371 176764 118437 176765
rect 118371 176700 118372 176764
rect 118436 176700 118437 176764
rect 118371 176699 118437 176700
rect 118374 175130 118434 176699
rect 119478 175130 119538 177651
rect 120763 177172 120829 177173
rect 120763 177108 120764 177172
rect 120828 177108 120829 177172
rect 120763 177107 120829 177108
rect 120766 175130 120826 177107
rect 120954 176600 121574 194058
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 121867 177716 121933 177717
rect 121867 177652 121868 177716
rect 121932 177652 121933 177716
rect 121867 177651 121933 177652
rect 121870 175130 121930 177651
rect 124443 176764 124509 176765
rect 124443 176700 124444 176764
rect 124508 176700 124509 176764
rect 124443 176699 124509 176700
rect 125731 176764 125797 176765
rect 125731 176700 125732 176764
rect 125796 176700 125797 176764
rect 125731 176699 125797 176700
rect 127019 176764 127085 176765
rect 127019 176700 127020 176764
rect 127084 176700 127085 176764
rect 127019 176699 127085 176700
rect 124446 175130 124506 176699
rect 125734 175130 125794 176699
rect 127022 175130 127082 176699
rect 127794 176600 128414 200898
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 129411 177716 129477 177717
rect 129411 177652 129412 177716
rect 129476 177652 129477 177716
rect 129411 177651 129477 177652
rect 130699 177716 130765 177717
rect 130699 177652 130700 177716
rect 130764 177652 130765 177716
rect 130699 177651 130765 177652
rect 128123 175404 128189 175405
rect 128123 175340 128124 175404
rect 128188 175340 128189 175404
rect 128123 175339 128189 175340
rect 128126 175130 128186 175339
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 177651
rect 130702 175130 130762 177651
rect 131514 176600 132134 204618
rect 135234 352894 135854 388338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 137139 387972 137205 387973
rect 137139 387908 137140 387972
rect 137204 387908 137205 387972
rect 137139 387907 137205 387908
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 137142 301477 137202 387907
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 137139 301476 137205 301477
rect 137139 301412 137140 301476
rect 137204 301412 137205 301476
rect 137139 301411 137205 301412
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 132355 177716 132421 177717
rect 132355 177652 132356 177716
rect 132420 177652 132421 177716
rect 132355 177651 132421 177652
rect 132358 175130 132418 177651
rect 133091 177172 133157 177173
rect 133091 177108 133092 177172
rect 133156 177108 133157 177172
rect 133091 177107 133157 177108
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123069 174996 123135 174997
rect 123069 174932 123070 174996
rect 123134 174932 123135 174996
rect 123069 174931 123135 174932
rect 123072 174494 123132 174931
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 177107
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 134382 175130 134442 176699
rect 135234 176600 135854 208338
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176600 139574 212058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 135667 175540 135733 175541
rect 135667 175476 135668 175540
rect 135732 175476 135733 175540
rect 135667 175475 135733 175476
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135670 175130 135730 175475
rect 148182 175130 148242 176699
rect 149514 176600 150134 186618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 176600 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 170259 239460 170325 239461
rect 170259 239396 170260 239460
rect 170324 239396 170325 239460
rect 170259 239395 170325 239396
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 166211 176900 166277 176901
rect 166211 176836 166212 176900
rect 166276 176836 166277 176900
rect 166211 176835 166277 176836
rect 158851 175404 158917 175405
rect 158851 175340 158852 175404
rect 158916 175340 158917 175404
rect 158851 175339 158917 175340
rect 158854 175130 158914 175339
rect 135670 175070 135780 175130
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 166214 160173 166274 176835
rect 167514 169174 168134 204618
rect 168235 177036 168301 177037
rect 168235 176972 168236 177036
rect 168300 176972 168301 177036
rect 168235 176971 168301 176972
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 166211 160172 166277 160173
rect 166211 160108 166212 160172
rect 166276 160108 166277 160172
rect 166211 160107 166277 160108
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 166395 134196 166461 134197
rect 166395 134132 166396 134196
rect 166460 134132 166461 134196
rect 166395 134131 166461 134132
rect 166211 130116 166277 130117
rect 166211 130052 166212 130116
rect 166276 130052 166277 130116
rect 166211 130051 166277 130052
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 61883 68916 61949 68917
rect 61883 68852 61884 68916
rect 61948 68852 61949 68916
rect 61883 68851 61949 68852
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 64894 63854 100338
rect 74656 94890 74716 95200
rect 74656 94830 74826 94890
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 93100
rect 74766 92445 74826 94830
rect 84312 94754 84372 95200
rect 85536 94754 85596 95200
rect 86624 94754 86684 95200
rect 87984 94754 88044 95200
rect 88936 94754 88996 95200
rect 84312 94694 84394 94754
rect 85536 94694 85866 94754
rect 86624 94694 86786 94754
rect 87984 94694 88074 94754
rect 74763 92444 74829 92445
rect 74763 92380 74764 92444
rect 74828 92380 74829 92444
rect 74763 92379 74829 92380
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 92445 84394 94694
rect 84331 92444 84397 92445
rect 84331 92380 84332 92444
rect 84396 92380 84397 92444
rect 84331 92379 84397 92380
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 85806 91221 85866 94694
rect 86726 91221 86786 94694
rect 88014 91221 88074 94694
rect 88934 94694 88996 94754
rect 90160 94754 90220 95200
rect 91384 94754 91444 95200
rect 90160 94694 90282 94754
rect 88934 92445 88994 94694
rect 88931 92444 88997 92445
rect 88931 92380 88932 92444
rect 88996 92380 88997 92444
rect 88931 92379 88997 92380
rect 90222 91221 90282 94694
rect 91326 94694 91444 94754
rect 92472 94754 92532 95200
rect 93832 94757 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 93829 94756 93895 94757
rect 92472 94694 92674 94754
rect 91326 91221 91386 94694
rect 85803 91220 85869 91221
rect 85803 91156 85804 91220
rect 85868 91156 85869 91220
rect 85803 91155 85869 91156
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 88011 91220 88077 91221
rect 88011 91156 88012 91220
rect 88076 91156 88077 91220
rect 88011 91155 88077 91156
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94694
rect 93829 94692 93830 94756
rect 93894 94692 93895 94756
rect 93829 94691 93895 94692
rect 95006 91221 95066 94830
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91357 96722 94830
rect 96659 91356 96725 91357
rect 96659 91292 96660 91356
rect 96724 91292 96725 91356
rect 96659 91291 96725 91292
rect 97214 91221 97274 94830
rect 98134 92445 98194 94830
rect 98131 92444 98197 92445
rect 98131 92380 98132 92444
rect 98196 92380 98197 92444
rect 98131 92379 98197 92380
rect 98502 91357 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 99544 94830 100034 94890
rect 98499 91356 98565 91357
rect 98499 91292 98500 91356
rect 98564 91292 98565 91356
rect 98499 91291 98565 91292
rect 99054 91221 99114 94830
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 99051 91220 99117 91221
rect 99051 91156 99052 91220
rect 99116 91156 99117 91220
rect 99051 91155 99117 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 91765 100034 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 99971 91764 100037 91765
rect 99971 91700 99972 91764
rect 100036 91700 100037 91764
rect 99971 91699 100037 91700
rect 100526 91221 100586 94830
rect 100894 91221 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 101814 91357 101874 94830
rect 101998 91493 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 102918 93870 102978 94830
rect 102734 93810 102978 93870
rect 102734 91765 102794 93810
rect 103286 93261 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 103283 93260 103349 93261
rect 103283 93196 103284 93260
rect 103348 93196 103349 93260
rect 103283 93195 103349 93196
rect 102731 91764 102797 91765
rect 102731 91700 102732 91764
rect 102796 91700 102797 91764
rect 102731 91699 102797 91700
rect 101995 91492 102061 91493
rect 101995 91428 101996 91492
rect 102060 91428 102061 91492
rect 101995 91427 102061 91428
rect 101811 91356 101877 91357
rect 101811 91292 101812 91356
rect 101876 91292 101877 91356
rect 101811 91291 101877 91292
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 100891 91220 100957 91221
rect 100891 91156 100892 91220
rect 100956 91156 100957 91220
rect 100891 91155 100957 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 91357 104266 94830
rect 104203 91356 104269 91357
rect 104203 91292 104204 91356
rect 104268 91292 104269 91356
rect 104203 91291 104269 91292
rect 104574 91221 104634 94830
rect 105494 91221 105554 94830
rect 105678 92445 105738 94830
rect 106414 94830 106540 94890
rect 105675 92444 105741 92445
rect 105675 92380 105676 92444
rect 105740 92380 105741 92444
rect 105675 92379 105741 92380
rect 106414 91221 106474 94830
rect 106616 94757 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 106613 94756 106679 94757
rect 106613 94692 106614 94756
rect 106678 94692 106679 94756
rect 106613 94691 106679 94692
rect 107702 91357 107762 94830
rect 107699 91356 107765 91357
rect 107699 91292 107700 91356
rect 107764 91292 107765 91356
rect 107699 91291 107765 91292
rect 108070 91221 108130 94830
rect 109174 91357 109234 94830
rect 109171 91356 109237 91357
rect 109171 91292 109172 91356
rect 109236 91292 109237 91356
rect 109171 91291 109237 91292
rect 109542 91221 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 111920 94830 111994 94890
rect 110094 93261 110154 94830
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105491 91220 105557 91221
rect 105491 91156 105492 91220
rect 105556 91156 105557 91220
rect 105491 91155 105557 91156
rect 106411 91220 106477 91221
rect 106411 91156 106412 91220
rect 106476 91156 106477 91220
rect 106411 91155 106477 91156
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 91221 110706 94830
rect 111198 92445 111258 94830
rect 111195 92444 111261 92445
rect 111195 92380 111196 92444
rect 111260 92380 111261 92444
rect 111195 92379 111261 92380
rect 111934 91357 111994 94830
rect 112302 94830 112388 94890
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 113144 94830 113282 94890
rect 113688 94830 113834 94890
rect 111931 91356 111997 91357
rect 111931 91292 111932 91356
rect 111996 91292 111997 91356
rect 111931 91291 111997 91292
rect 112302 91221 112362 94830
rect 113222 92309 113282 94830
rect 113774 93533 113834 94830
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 114326 93669 114386 94830
rect 114323 93668 114389 93669
rect 114323 93604 114324 93668
rect 114388 93604 114389 93668
rect 114323 93603 114389 93604
rect 113771 93532 113837 93533
rect 113771 93468 113772 93532
rect 113836 93468 113837 93532
rect 113771 93467 113837 93468
rect 113219 92308 113285 92309
rect 113219 92244 113220 92308
rect 113284 92244 113285 92308
rect 113219 92243 113285 92244
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 112299 91220 112365 91221
rect 112299 91156 112300 91220
rect 112364 91156 112365 91220
rect 112299 91155 112365 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114878 91629 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115430 92445 115490 94830
rect 115427 92444 115493 92445
rect 115427 92380 115428 92444
rect 115492 92380 115493 92444
rect 115427 92379 115493 92380
rect 114875 91628 114941 91629
rect 114875 91564 114876 91628
rect 114940 91564 114941 91628
rect 114875 91563 114941 91564
rect 115798 91221 115858 94830
rect 116718 91221 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 117904 94830 118066 94890
rect 117086 91357 117146 94830
rect 117083 91356 117149 91357
rect 117083 91292 117084 91356
rect 117148 91292 117149 91356
rect 117083 91291 117149 91292
rect 115795 91220 115861 91221
rect 115795 91156 115796 91220
rect 115860 91156 115861 91220
rect 115795 91155 115861 91156
rect 116715 91220 116781 91221
rect 116715 91156 116716 91220
rect 116780 91156 116781 91220
rect 116715 91155 116781 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 91221 118066 94830
rect 118176 94757 118236 95200
rect 119400 94890 119460 95200
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 119536 94830 119722 94890
rect 118173 94756 118239 94757
rect 118173 94692 118174 94756
rect 118238 94692 118239 94756
rect 118173 94691 118239 94692
rect 119294 92173 119354 94830
rect 119291 92172 119357 92173
rect 119291 92108 119292 92172
rect 119356 92108 119357 92172
rect 119291 92107 119357 92108
rect 119662 91221 119722 94830
rect 120214 94830 120276 94890
rect 120214 91901 120274 94830
rect 120624 94757 120684 95200
rect 121712 94890 121772 95200
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 120621 94756 120687 94757
rect 120621 94692 120622 94756
rect 120686 94692 120687 94756
rect 120621 94691 120687 94692
rect 120211 91900 120277 91901
rect 120211 91836 120212 91900
rect 120276 91836 120277 91900
rect 120211 91835 120277 91836
rect 118003 91220 118069 91221
rect 118003 91156 118004 91220
rect 118068 91156 118069 91220
rect 118003 91155 118069 91156
rect 119659 91220 119725 91221
rect 119659 91156 119660 91220
rect 119724 91156 119725 91220
rect 119659 91155 119725 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 121686 91357 121746 94830
rect 121683 91356 121749 91357
rect 121683 91292 121684 91356
rect 121748 91292 121749 91356
rect 121683 91291 121749 91292
rect 122054 91221 122114 94830
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122606 91354 122666 93810
rect 123158 91357 123218 94830
rect 123155 91356 123221 91357
rect 122606 91294 122850 91354
rect 122790 91221 122850 91294
rect 123155 91292 123156 91356
rect 123220 91292 123221 91356
rect 123155 91291 123221 91292
rect 124078 91221 124138 94830
rect 124446 92445 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125978 94890
rect 124443 92444 124509 92445
rect 124443 92380 124444 92444
rect 124508 92380 124509 92444
rect 124443 92379 124509 92380
rect 125366 91221 125426 94830
rect 125918 92445 125978 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 126470 92445 126530 94830
rect 125915 92444 125981 92445
rect 125915 92380 125916 92444
rect 125980 92380 125981 92444
rect 125915 92379 125981 92380
rect 126467 92444 126533 92445
rect 126467 92380 126468 92444
rect 126532 92380 126533 92444
rect 126467 92379 126533 92380
rect 126654 91221 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 127574 91221 127634 94830
rect 129414 93533 129474 94830
rect 129411 93532 129477 93533
rect 129411 93468 129412 93532
rect 129476 93468 129477 93532
rect 129411 93467 129477 93468
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 122787 91220 122853 91221
rect 122787 91156 122788 91220
rect 122852 91156 122853 91220
rect 122787 91155 122853 91156
rect 124075 91220 124141 91221
rect 124075 91156 124076 91220
rect 124140 91156 124141 91220
rect 124075 91155 124141 91156
rect 125363 91220 125429 91221
rect 125363 91156 125364 91220
rect 125428 91156 125429 91220
rect 125363 91155 125429 91156
rect 126651 91220 126717 91221
rect 126651 91156 126652 91220
rect 126716 91156 126717 91220
rect 126651 91155 126717 91156
rect 127571 91220 127637 91221
rect 127571 91156 127572 91220
rect 127636 91156 127637 91220
rect 127571 91155 127637 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 130702 91221 130762 94830
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 91629 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 133094 92445 133154 94830
rect 133091 92444 133157 92445
rect 133091 92380 133092 92444
rect 133156 92380 133157 92444
rect 133091 92379 133157 92380
rect 132355 91628 132421 91629
rect 132355 91564 132356 91628
rect 132420 91564 132421 91628
rect 132355 91563 132421 91564
rect 134382 91221 134442 94830
rect 134379 91220 134445 91221
rect 134379 91156 134380 91220
rect 134444 91156 134445 91220
rect 134379 91155 134445 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 92445 136098 94830
rect 151310 94830 151556 94890
rect 136035 92444 136101 92445
rect 136035 92380 136036 92444
rect 136100 92380 136101 92444
rect 136035 92379 136101 92380
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151310 91221 151370 94830
rect 151491 94756 151557 94757
rect 151491 94692 151492 94756
rect 151556 94692 151557 94756
rect 151491 94691 151557 94692
rect 151494 92445 151554 94691
rect 151632 94210 151692 95200
rect 151768 94757 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151765 94756 151831 94757
rect 151765 94692 151766 94756
rect 151830 94692 151831 94756
rect 151765 94691 151831 94692
rect 151632 94150 151738 94210
rect 151678 93669 151738 94150
rect 151675 93668 151741 93669
rect 151675 93604 151676 93668
rect 151740 93604 151741 93668
rect 151675 93603 151741 93604
rect 152046 92445 152106 94830
rect 151491 92444 151557 92445
rect 151491 92380 151492 92444
rect 151556 92380 151557 92444
rect 151491 92379 151557 92380
rect 152043 92444 152109 92445
rect 152043 92380 152044 92444
rect 152108 92380 152109 92444
rect 152043 92379 152109 92380
rect 151307 91220 151373 91221
rect 151307 91156 151308 91220
rect 151372 91156 151373 91220
rect 151307 91155 151373 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 82789 166274 130051
rect 166398 88229 166458 134131
rect 167514 133174 168134 168618
rect 168238 157997 168298 176971
rect 168235 157996 168301 157997
rect 168235 157932 168236 157996
rect 168300 157932 168301 157996
rect 168235 157931 168301 157932
rect 168235 139500 168301 139501
rect 168235 139436 168236 139500
rect 168300 139436 168301 139500
rect 168235 139435 168301 139436
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166395 88228 166461 88229
rect 166395 88164 166396 88228
rect 166460 88164 166461 88228
rect 166395 88163 166461 88164
rect 166211 82788 166277 82789
rect 166211 82724 166212 82788
rect 166276 82724 166277 82788
rect 166211 82723 166277 82724
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 96618
rect 168238 89725 168298 139435
rect 168971 136916 169037 136917
rect 168971 136852 168972 136916
rect 169036 136852 169037 136916
rect 168971 136851 169037 136852
rect 168235 89724 168301 89725
rect 168235 89660 168236 89724
rect 168300 89660 168301 89724
rect 168235 89659 168301 89660
rect 168974 82653 169034 136851
rect 169155 129980 169221 129981
rect 169155 129916 169156 129980
rect 169220 129916 169221 129980
rect 169155 129915 169221 129916
rect 169158 85509 169218 129915
rect 170262 95573 170322 239395
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 170443 127260 170509 127261
rect 170443 127196 170444 127260
rect 170508 127196 170509 127260
rect 170443 127195 170509 127196
rect 170259 95572 170325 95573
rect 170259 95508 170260 95572
rect 170324 95508 170325 95572
rect 170259 95507 170325 95508
rect 169155 85508 169221 85509
rect 169155 85444 169156 85508
rect 169220 85444 169221 85508
rect 169155 85443 169221 85444
rect 168971 82652 169037 82653
rect 168971 82588 168972 82652
rect 169036 82588 169037 82652
rect 168971 82587 169037 82588
rect 170446 81429 170506 127195
rect 171234 100894 171854 136338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 177251 294132 177317 294133
rect 177251 294068 177252 294132
rect 177316 294068 177317 294132
rect 177251 294067 177317 294068
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 173019 131204 173085 131205
rect 173019 131140 173020 131204
rect 173084 131140 173085 131204
rect 173019 131139 173085 131140
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 170443 81428 170509 81429
rect 170443 81364 170444 81428
rect 170508 81364 170509 81428
rect 170443 81363 170509 81364
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 100338
rect 173022 81293 173082 131139
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 173019 81292 173085 81293
rect 173019 81228 173020 81292
rect 173084 81228 173085 81292
rect 173019 81227 173085 81228
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 68614 175574 104058
rect 177254 95165 177314 294067
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 177251 95164 177317 95165
rect 177251 95100 177252 95164
rect 177316 95100 177317 95164
rect 177251 95099 177317 95100
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 227667 281892 227733 281893
rect 227667 281828 227668 281892
rect 227732 281828 227733 281892
rect 227667 281827 227733 281828
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 227670 175130 227730 281827
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 241835 334660 241901 334661
rect 241835 334596 241836 334660
rect 241900 334596 241901 334660
rect 241835 334595 241901 334596
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 236499 296988 236565 296989
rect 236499 296924 236500 296988
rect 236564 296924 236565 296988
rect 236499 296923 236565 296924
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 233187 216068 233253 216069
rect 233187 216004 233188 216068
rect 233252 216004 233253 216068
rect 233187 216003 233253 216004
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 178000 229574 194058
rect 231899 180028 231965 180029
rect 231899 179964 231900 180028
rect 231964 179964 231965 180028
rect 231899 179963 231965 179964
rect 228955 177852 229021 177853
rect 228955 177788 228956 177852
rect 229020 177788 229021 177852
rect 228955 177787 229021 177788
rect 228958 175810 229018 177787
rect 228958 175750 229202 175810
rect 229142 175269 229202 175750
rect 229139 175268 229205 175269
rect 229139 175204 229140 175268
rect 229204 175204 229205 175268
rect 229139 175203 229205 175204
rect 227670 175070 229202 175130
rect 229142 174725 229202 175070
rect 229139 174724 229205 174725
rect 229139 174660 229140 174724
rect 229204 174660 229205 174724
rect 229139 174659 229205 174660
rect 221207 165454 221527 165486
rect 221207 165218 221249 165454
rect 221485 165218 221527 165454
rect 221207 165134 221527 165218
rect 221207 164898 221249 165134
rect 221485 164898 221527 165134
rect 221207 164866 221527 164898
rect 224471 165454 224791 165486
rect 224471 165218 224513 165454
rect 224749 165218 224791 165454
rect 224471 165134 224791 165218
rect 224471 164898 224513 165134
rect 224749 164898 224791 165134
rect 224471 164866 224791 164898
rect 231163 154596 231229 154597
rect 231163 154532 231164 154596
rect 231228 154532 231229 154596
rect 231163 154531 231229 154532
rect 219575 147454 219895 147486
rect 219575 147218 219617 147454
rect 219853 147218 219895 147454
rect 219575 147134 219895 147218
rect 219575 146898 219617 147134
rect 219853 146898 219895 147134
rect 219575 146866 219895 146898
rect 222839 147454 223159 147486
rect 222839 147218 222881 147454
rect 223117 147218 223159 147454
rect 222839 147134 223159 147218
rect 222839 146898 222881 147134
rect 223117 146898 223159 147134
rect 222839 146866 223159 146898
rect 226103 147454 226423 147486
rect 226103 147218 226145 147454
rect 226381 147218 226423 147454
rect 226103 147134 226423 147218
rect 226103 146898 226145 147134
rect 226381 146898 226423 147134
rect 226103 146866 226423 146898
rect 230979 142764 231045 142765
rect 230979 142700 230980 142764
rect 231044 142700 231045 142764
rect 230979 142699 231045 142700
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 221207 129454 221527 129486
rect 221207 129218 221249 129454
rect 221485 129218 221527 129454
rect 221207 129134 221527 129218
rect 221207 128898 221249 129134
rect 221485 128898 221527 129134
rect 221207 128866 221527 128898
rect 224471 129454 224791 129486
rect 224471 129218 224513 129454
rect 224749 129218 224791 129454
rect 224471 129134 224791 129218
rect 224471 128898 224513 129134
rect 224749 128898 224791 129134
rect 224471 128866 224791 128898
rect 219575 111454 219895 111486
rect 219575 111218 219617 111454
rect 219853 111218 219895 111454
rect 219575 111134 219895 111218
rect 219575 110898 219617 111134
rect 219853 110898 219895 111134
rect 219575 110866 219895 110898
rect 222839 111454 223159 111486
rect 222839 111218 222881 111454
rect 223117 111218 223159 111454
rect 222839 111134 223159 111218
rect 222839 110898 222881 111134
rect 223117 110898 223159 111134
rect 222839 110866 223159 110898
rect 226103 111454 226423 111486
rect 226103 111218 226145 111454
rect 226381 111218 226423 111454
rect 226103 111134 226423 111218
rect 226103 110898 226145 111134
rect 226381 110898 226423 111134
rect 226103 110866 226423 110898
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 214419 102508 214485 102509
rect 214419 102444 214420 102508
rect 214484 102444 214485 102508
rect 214419 102443 214485 102444
rect 214422 91085 214482 102443
rect 230982 102373 231042 142699
rect 231166 117061 231226 154531
rect 231902 136373 231962 179963
rect 233190 153373 233250 216003
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 233371 185604 233437 185605
rect 233371 185540 233372 185604
rect 233436 185540 233437 185604
rect 233371 185539 233437 185540
rect 233187 153372 233253 153373
rect 233187 153308 233188 153372
rect 233252 153308 233253 153372
rect 233187 153307 233253 153308
rect 233374 148749 233434 185539
rect 234659 177444 234725 177445
rect 234659 177380 234660 177444
rect 234724 177380 234725 177444
rect 234659 177379 234725 177380
rect 234662 150109 234722 177379
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 234659 150108 234725 150109
rect 234659 150044 234660 150108
rect 234724 150044 234725 150108
rect 234659 150043 234725 150044
rect 233371 148748 233437 148749
rect 233371 148684 233372 148748
rect 233436 148684 233437 148748
rect 233371 148683 233437 148684
rect 233739 146980 233805 146981
rect 233739 146916 233740 146980
rect 233804 146916 233805 146980
rect 233739 146915 233805 146916
rect 231899 136372 231965 136373
rect 231899 136308 231900 136372
rect 231964 136308 231965 136372
rect 231899 136307 231965 136308
rect 232451 125900 232517 125901
rect 232451 125836 232452 125900
rect 232516 125836 232517 125900
rect 232451 125835 232517 125836
rect 231163 117060 231229 117061
rect 231163 116996 231164 117060
rect 231228 116996 231229 117060
rect 231163 116995 231229 116996
rect 230979 102372 231045 102373
rect 230979 102308 230980 102372
rect 231044 102308 231045 102372
rect 230979 102307 231045 102308
rect 229139 97204 229205 97205
rect 229139 97140 229140 97204
rect 229204 97140 229205 97204
rect 229139 97139 229205 97140
rect 229142 96930 229202 97139
rect 228590 96870 229202 96930
rect 227667 95300 227733 95301
rect 227667 95236 227668 95300
rect 227732 95236 227733 95300
rect 227667 95235 227733 95236
rect 214419 91084 214485 91085
rect 214419 91020 214420 91084
rect 214484 91020 214485 91084
rect 214419 91019 214485 91020
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 227670 70277 227730 95235
rect 228590 84210 228650 96870
rect 229139 96660 229205 96661
rect 229139 96630 229140 96660
rect 228958 96596 229140 96630
rect 229204 96596 229205 96660
rect 228958 96595 229205 96596
rect 228958 96570 229202 96595
rect 228958 95301 229018 96570
rect 228955 95300 229021 95301
rect 228955 95236 228956 95300
rect 229020 95236 229021 95300
rect 228955 95235 229021 95236
rect 228222 84150 228650 84210
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 227667 70276 227733 70277
rect 227667 70212 227668 70276
rect 227732 70212 227733 70276
rect 227667 70211 227733 70212
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 228222 17237 228282 84150
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228219 17236 228285 17237
rect 228219 17172 228220 17236
rect 228284 17172 228285 17236
rect 228219 17171 228285 17172
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 232454 14517 232514 125835
rect 233742 105637 233802 146915
rect 235794 129454 236414 164898
rect 236502 142085 236562 296923
rect 239514 277174 240134 312618
rect 240363 312492 240429 312493
rect 240363 312428 240364 312492
rect 240428 312428 240429 312492
rect 240363 312427 240429 312428
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 238523 198116 238589 198117
rect 238523 198052 238524 198116
rect 238588 198052 238589 198116
rect 238523 198051 238589 198052
rect 237419 195260 237485 195261
rect 237419 195196 237420 195260
rect 237484 195196 237485 195260
rect 237419 195195 237485 195196
rect 237422 164797 237482 195195
rect 237603 178668 237669 178669
rect 237603 178604 237604 178668
rect 237668 178604 237669 178668
rect 237603 178603 237669 178604
rect 237419 164796 237485 164797
rect 237419 164732 237420 164796
rect 237484 164732 237485 164796
rect 237419 164731 237485 164732
rect 237606 157453 237666 178603
rect 238526 168330 238586 198051
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 238707 168332 238773 168333
rect 238707 168330 238708 168332
rect 238526 168270 238708 168330
rect 238707 168268 238708 168270
rect 238772 168268 238773 168332
rect 238707 168267 238773 168268
rect 239259 164524 239325 164525
rect 239259 164460 239260 164524
rect 239324 164460 239325 164524
rect 239259 164459 239325 164460
rect 237603 157452 237669 157453
rect 237603 157388 237604 157452
rect 237668 157388 237669 157452
rect 237603 157387 237669 157388
rect 237971 152420 238037 152421
rect 237971 152356 237972 152420
rect 238036 152356 238037 152420
rect 237971 152355 238037 152356
rect 236499 142084 236565 142085
rect 236499 142020 236500 142084
rect 236564 142020 236565 142084
rect 236499 142019 236565 142020
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 233739 105636 233805 105637
rect 233739 105572 233740 105636
rect 233804 105572 233805 105636
rect 233739 105571 233805 105572
rect 235794 93454 236414 128898
rect 237974 111757 238034 152355
rect 239262 124813 239322 164459
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239259 124812 239325 124813
rect 239259 124748 239260 124812
rect 239324 124748 239325 124812
rect 239259 124747 239325 124748
rect 237971 111756 238037 111757
rect 237971 111692 237972 111756
rect 238036 111692 238037 111756
rect 237971 111691 238037 111692
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 232451 14516 232517 14517
rect 232451 14452 232452 14516
rect 232516 14452 232517 14516
rect 232451 14451 232517 14452
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 240366 43621 240426 312427
rect 241651 296852 241717 296853
rect 241651 296788 241652 296852
rect 241716 296788 241717 296852
rect 241651 296787 241717 296788
rect 240547 177308 240613 177309
rect 240547 177244 240548 177308
rect 240612 177244 240613 177308
rect 240547 177243 240613 177244
rect 240550 167653 240610 177243
rect 240547 167652 240613 167653
rect 240547 167588 240548 167652
rect 240612 167588 240613 167652
rect 240547 167587 240613 167588
rect 241654 152557 241714 296787
rect 241651 152556 241717 152557
rect 241651 152492 241652 152556
rect 241716 152492 241717 152556
rect 241651 152491 241717 152492
rect 240363 43620 240429 43621
rect 240363 43556 240364 43620
rect 240428 43556 240429 43620
rect 240363 43555 240429 43556
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 240366 11797 240426 43555
rect 241838 35189 241898 334595
rect 243234 316894 243854 352338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 252875 376004 252941 376005
rect 252875 375940 252876 376004
rect 252940 375940 252941 376004
rect 252875 375939 252941 375940
rect 251219 367708 251285 367709
rect 251219 367644 251220 367708
rect 251284 367644 251285 367708
rect 251219 367643 251285 367644
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 245699 330444 245765 330445
rect 245699 330380 245700 330444
rect 245764 330380 245765 330444
rect 245699 330379 245765 330380
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 242939 308412 243005 308413
rect 242939 308348 242940 308412
rect 243004 308348 243005 308412
rect 242939 308347 243005 308348
rect 242942 46341 243002 308347
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 244227 186964 244293 186965
rect 244227 186900 244228 186964
rect 244292 186900 244293 186964
rect 244227 186899 244293 186900
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 244230 147253 244290 186899
rect 244227 147252 244293 147253
rect 244227 147188 244228 147252
rect 244292 147188 244293 147252
rect 244227 147187 244293 147188
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 244779 129028 244845 129029
rect 244779 128964 244780 129028
rect 244844 128964 244845 129028
rect 244779 128963 244845 128964
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 242939 46340 243005 46341
rect 242939 46276 242940 46340
rect 243004 46276 243005 46340
rect 242939 46275 243005 46276
rect 241835 35188 241901 35189
rect 241835 35124 241836 35188
rect 241900 35124 241901 35188
rect 241835 35123 241901 35124
rect 241838 11797 241898 35123
rect 242942 11797 243002 46275
rect 243234 28894 243854 64338
rect 244782 32469 244842 128963
rect 244779 32468 244845 32469
rect 244779 32404 244780 32468
rect 244844 32404 244845 32468
rect 244779 32403 244845 32404
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 240363 11796 240429 11797
rect 240363 11732 240364 11796
rect 240428 11732 240429 11796
rect 240363 11731 240429 11732
rect 241835 11796 241901 11797
rect 241835 11732 241836 11796
rect 241900 11732 241901 11796
rect 241835 11731 241901 11732
rect 242939 11796 243005 11797
rect 242939 11732 242940 11796
rect 243004 11732 243005 11796
rect 242939 11731 243005 11732
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 28338
rect 245702 22677 245762 330379
rect 246954 320614 247574 356058
rect 250299 333300 250365 333301
rect 250299 333236 250300 333300
rect 250364 333236 250365 333300
rect 250299 333235 250365 333236
rect 248459 331804 248525 331805
rect 248459 331740 248460 331804
rect 248524 331740 248525 331804
rect 248459 331739 248525 331740
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 247723 309772 247789 309773
rect 247723 309708 247724 309772
rect 247788 309708 247789 309772
rect 247723 309707 247789 309708
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 245883 182884 245949 182885
rect 245883 182820 245884 182884
rect 245948 182820 245949 182884
rect 245883 182819 245949 182820
rect 245886 144941 245946 182819
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 245883 144940 245949 144941
rect 245883 144876 245884 144940
rect 245948 144876 245949 144940
rect 245883 144875 245949 144876
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 247726 48381 247786 309707
rect 247723 48380 247789 48381
rect 247723 48316 247724 48380
rect 247788 48316 247789 48380
rect 247723 48315 247789 48316
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 245699 22676 245765 22677
rect 245699 22612 245700 22676
rect 245764 22612 245765 22676
rect 245699 22611 245765 22612
rect 245702 11797 245762 22611
rect 245699 11796 245765 11797
rect 245699 11732 245700 11796
rect 245764 11732 245765 11796
rect 245699 11731 245765 11732
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 247726 3501 247786 48315
rect 248462 37909 248522 331739
rect 249011 127668 249077 127669
rect 249011 127604 249012 127668
rect 249076 127604 249077 127668
rect 249011 127603 249077 127604
rect 249014 42125 249074 127603
rect 249011 42124 249077 42125
rect 249011 42060 249012 42124
rect 249076 42060 249077 42124
rect 249011 42059 249077 42060
rect 248459 37908 248525 37909
rect 248459 37844 248460 37908
rect 248524 37844 248525 37908
rect 248459 37843 248525 37844
rect 248462 15605 248522 37843
rect 248459 15604 248525 15605
rect 248459 15540 248460 15604
rect 248524 15540 248525 15604
rect 248459 15539 248525 15540
rect 250302 3909 250362 333235
rect 251222 8261 251282 367643
rect 252691 302292 252757 302293
rect 252691 302228 252692 302292
rect 252756 302228 252757 302292
rect 252691 302227 252757 302228
rect 252694 140181 252754 302227
rect 252691 140180 252757 140181
rect 252691 140116 252692 140180
rect 252756 140116 252757 140180
rect 252691 140115 252757 140116
rect 252878 24309 252938 375939
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 255267 360908 255333 360909
rect 255267 360844 255268 360908
rect 255332 360844 255333 360908
rect 255267 360843 255333 360844
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 255270 39405 255330 360843
rect 257514 331174 258134 366618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 258395 336020 258461 336021
rect 258395 335956 258396 336020
rect 258460 335956 258461 336020
rect 258395 335955 258461 335956
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 258398 316050 258458 335955
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257291 130252 257357 130253
rect 257291 130188 257292 130252
rect 257356 130188 257357 130252
rect 257291 130187 257357 130188
rect 257294 72453 257354 130187
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257291 72452 257357 72453
rect 257291 72388 257292 72452
rect 257356 72388 257357 72452
rect 257291 72387 257357 72388
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 255267 39404 255333 39405
rect 255267 39340 255268 39404
rect 255332 39340 255333 39404
rect 255267 39339 255333 39340
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 252875 24308 252941 24309
rect 252875 24244 252876 24308
rect 252940 24244 252941 24308
rect 252875 24243 252941 24244
rect 252878 11797 252938 24243
rect 252875 11796 252941 11797
rect 252875 11732 252876 11796
rect 252940 11732 252941 11796
rect 252875 11731 252941 11732
rect 251219 8260 251285 8261
rect 251219 8196 251220 8260
rect 251284 8196 251285 8260
rect 251219 8195 251285 8196
rect 250299 3908 250365 3909
rect 250299 3844 250300 3908
rect 250364 3844 250365 3908
rect 250299 3843 250365 3844
rect 247723 3500 247789 3501
rect 247723 3436 247724 3500
rect 247788 3436 247789 3500
rect 247723 3435 247789 3436
rect 253794 3454 254414 38898
rect 255270 11797 255330 39339
rect 255267 11796 255333 11797
rect 255267 11732 255268 11796
rect 255332 11732 255333 11796
rect 255267 11731 255333 11732
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 42618
rect 258214 315990 258458 316050
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 258214 16590 258274 315990
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 260051 126444 260117 126445
rect 260051 126380 260052 126444
rect 260116 126380 260117 126444
rect 260051 126379 260117 126380
rect 260054 73813 260114 126379
rect 261234 118894 261854 154338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 268331 385388 268397 385389
rect 268331 385324 268332 385388
rect 268396 385324 268397 385388
rect 268331 385323 268397 385324
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264099 139500 264165 139501
rect 264099 139436 264100 139500
rect 264164 139436 264165 139500
rect 264099 139435 264165 139436
rect 262811 129844 262877 129845
rect 262811 129780 262812 129844
rect 262876 129780 262877 129844
rect 262811 129779 262877 129780
rect 262075 119100 262141 119101
rect 262075 119036 262076 119100
rect 262140 119036 262141 119100
rect 262075 119035 262141 119036
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 260051 73812 260117 73813
rect 260051 73748 260052 73812
rect 260116 73748 260117 73812
rect 260051 73747 260117 73748
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 258214 16530 258458 16590
rect 258398 10981 258458 16530
rect 258395 10980 258461 10981
rect 258395 10916 258396 10980
rect 258460 10916 258461 10980
rect 258395 10915 258461 10916
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 262078 2005 262138 119035
rect 262814 26893 262874 129779
rect 262995 112708 263061 112709
rect 262995 112644 262996 112708
rect 263060 112644 263061 112708
rect 262995 112643 263061 112644
rect 262998 36549 263058 112643
rect 262995 36548 263061 36549
rect 262995 36484 262996 36548
rect 263060 36484 263061 36548
rect 262995 36483 263061 36484
rect 262811 26892 262877 26893
rect 262811 26828 262812 26892
rect 262876 26828 262877 26892
rect 262811 26827 262877 26828
rect 264102 25533 264162 139435
rect 264954 122614 265574 158058
rect 265755 150516 265821 150517
rect 265755 150452 265756 150516
rect 265820 150452 265821 150516
rect 265755 150451 265821 150452
rect 265758 146437 265818 150451
rect 265755 146436 265821 146437
rect 265755 146372 265756 146436
rect 265820 146372 265821 146436
rect 265755 146371 265821 146372
rect 265755 129028 265821 129029
rect 265755 128964 265756 129028
rect 265820 128964 265821 129028
rect 265755 128963 265821 128964
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264283 107132 264349 107133
rect 264283 107068 264284 107132
rect 264348 107068 264349 107132
rect 264283 107067 264349 107068
rect 264286 50285 264346 107067
rect 264954 86614 265574 122058
rect 265758 90405 265818 128963
rect 265755 90404 265821 90405
rect 265755 90340 265756 90404
rect 265820 90340 265821 90404
rect 265755 90339 265821 90340
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264283 50284 264349 50285
rect 264283 50220 264284 50284
rect 264348 50220 264349 50284
rect 264283 50219 264349 50220
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264099 25532 264165 25533
rect 264099 25468 264100 25532
rect 264164 25468 264165 25532
rect 264099 25467 264165 25468
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 262075 2004 262141 2005
rect 262075 1940 262076 2004
rect 262140 1940 262141 2004
rect 262075 1939 262141 1940
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 268334 4045 268394 385323
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 178000 272414 200898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 178000 276134 204618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279003 178668 279069 178669
rect 279003 178604 279004 178668
rect 279068 178604 279069 178668
rect 279003 178603 279069 178604
rect 279006 173770 279066 178603
rect 279234 178000 279854 208338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 285627 286516 285693 286517
rect 285627 286452 285628 286516
rect 285692 286452 285693 286516
rect 285627 286451 285693 286452
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 280291 199340 280357 199341
rect 280291 199276 280292 199340
rect 280356 199276 280357 199340
rect 280291 199275 280357 199276
rect 279371 173772 279437 173773
rect 279371 173770 279372 173772
rect 279006 173710 279372 173770
rect 279371 173708 279372 173710
rect 279436 173708 279437 173772
rect 279371 173707 279437 173708
rect 272207 165454 272527 165486
rect 272207 165218 272249 165454
rect 272485 165218 272527 165454
rect 272207 165134 272527 165218
rect 272207 164898 272249 165134
rect 272485 164898 272527 165134
rect 272207 164866 272527 164898
rect 275471 165454 275791 165486
rect 275471 165218 275513 165454
rect 275749 165218 275791 165454
rect 275471 165134 275791 165218
rect 275471 164898 275513 165134
rect 275749 164898 275791 165134
rect 275471 164866 275791 164898
rect 268515 161668 268581 161669
rect 268515 161604 268516 161668
rect 268580 161604 268581 161668
rect 268515 161603 268581 161604
rect 268518 161261 268578 161603
rect 268515 161260 268581 161261
rect 268515 161196 268516 161260
rect 268580 161196 268581 161260
rect 268515 161195 268581 161196
rect 268515 147932 268581 147933
rect 268515 147868 268516 147932
rect 268580 147868 268581 147932
rect 268515 147867 268581 147868
rect 268518 146165 268578 147867
rect 270575 147454 270895 147486
rect 270575 147218 270617 147454
rect 270853 147218 270895 147454
rect 270575 147134 270895 147218
rect 270575 146898 270617 147134
rect 270853 146898 270895 147134
rect 270575 146866 270895 146898
rect 273839 147454 274159 147486
rect 273839 147218 273881 147454
rect 274117 147218 274159 147454
rect 273839 147134 274159 147218
rect 273839 146898 273881 147134
rect 274117 146898 274159 147134
rect 273839 146866 274159 146898
rect 277103 147454 277423 147486
rect 277103 147218 277145 147454
rect 277381 147218 277423 147454
rect 277103 147134 277423 147218
rect 277103 146898 277145 147134
rect 277381 146898 277423 147134
rect 277103 146866 277423 146898
rect 268515 146164 268581 146165
rect 268515 146100 268516 146164
rect 268580 146100 268581 146164
rect 268515 146099 268581 146100
rect 268515 141948 268581 141949
rect 268515 141884 268516 141948
rect 268580 141884 268581 141948
rect 268515 141883 268581 141884
rect 268518 140589 268578 141883
rect 268515 140588 268581 140589
rect 268515 140524 268516 140588
rect 268580 140524 268581 140588
rect 268515 140523 268581 140524
rect 272207 129454 272527 129486
rect 272207 129218 272249 129454
rect 272485 129218 272527 129454
rect 272207 129134 272527 129218
rect 272207 128898 272249 129134
rect 272485 128898 272527 129134
rect 272207 128866 272527 128898
rect 275471 129454 275791 129486
rect 275471 129218 275513 129454
rect 275749 129218 275791 129454
rect 275471 129134 275791 129218
rect 275471 128898 275513 129134
rect 275749 128898 275791 129134
rect 275471 128866 275791 128898
rect 268515 128620 268581 128621
rect 268515 128556 268516 128620
rect 268580 128556 268581 128620
rect 268515 128555 268581 128556
rect 268518 128213 268578 128555
rect 268515 128212 268581 128213
rect 268515 128148 268516 128212
rect 268580 128148 268581 128212
rect 268515 128147 268581 128148
rect 268515 127260 268581 127261
rect 268515 127196 268516 127260
rect 268580 127196 268581 127260
rect 268515 127195 268581 127196
rect 268518 126853 268578 127195
rect 268515 126852 268581 126853
rect 268515 126788 268516 126852
rect 268580 126788 268581 126852
rect 268515 126787 268581 126788
rect 268515 123044 268581 123045
rect 268515 122980 268516 123044
rect 268580 122980 268581 123044
rect 268515 122979 268581 122980
rect 268518 122637 268578 122979
rect 268515 122636 268581 122637
rect 268515 122572 268516 122636
rect 268580 122572 268581 122636
rect 268515 122571 268581 122572
rect 268515 121684 268581 121685
rect 268515 121620 268516 121684
rect 268580 121620 268581 121684
rect 268515 121619 268581 121620
rect 268518 121277 268578 121619
rect 268515 121276 268581 121277
rect 268515 121212 268516 121276
rect 268580 121212 268581 121276
rect 268515 121211 268581 121212
rect 268515 117332 268581 117333
rect 268515 117268 268516 117332
rect 268580 117268 268581 117332
rect 268515 117267 268581 117268
rect 268518 116517 268578 117267
rect 280294 117061 280354 199275
rect 282954 176614 283574 212058
rect 284339 192540 284405 192541
rect 284339 192476 284340 192540
rect 284404 192476 284405 192540
rect 284339 192475 284405 192476
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 280291 117060 280357 117061
rect 280291 116996 280292 117060
rect 280356 116996 280357 117060
rect 280291 116995 280357 116996
rect 268515 116516 268581 116517
rect 268515 116452 268516 116516
rect 268580 116452 268581 116516
rect 268515 116451 268581 116452
rect 270575 111454 270895 111486
rect 270575 111218 270617 111454
rect 270853 111218 270895 111454
rect 270575 111134 270895 111218
rect 270575 110898 270617 111134
rect 270853 110898 270895 111134
rect 270575 110866 270895 110898
rect 273839 111454 274159 111486
rect 273839 111218 273881 111454
rect 274117 111218 274159 111454
rect 273839 111134 274159 111218
rect 273839 110898 273881 111134
rect 274117 110898 274159 111134
rect 273839 110866 274159 110898
rect 277103 111454 277423 111486
rect 277103 111218 277145 111454
rect 277381 111218 277423 111454
rect 277103 111134 277423 111218
rect 277103 110898 277145 111134
rect 277381 110898 277423 111134
rect 277103 110866 277423 110898
rect 282954 104614 283574 140058
rect 284342 106317 284402 192475
rect 285630 124813 285690 286451
rect 285811 280532 285877 280533
rect 285811 280468 285812 280532
rect 285876 280468 285877 280532
rect 285811 280467 285877 280468
rect 285627 124812 285693 124813
rect 285627 124748 285628 124812
rect 285692 124748 285693 124812
rect 285627 124747 285693 124748
rect 285814 123997 285874 280467
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 287099 222868 287165 222869
rect 287099 222804 287100 222868
rect 287164 222804 287165 222868
rect 287099 222803 287165 222804
rect 285811 123996 285877 123997
rect 285811 123932 285812 123996
rect 285876 123932 285877 123996
rect 285811 123931 285877 123932
rect 284339 106316 284405 106317
rect 284339 106252 284340 106316
rect 284404 106252 284405 106316
rect 284339 106251 284405 106252
rect 287102 104957 287162 222803
rect 289794 219454 290414 254898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 295379 387020 295445 387021
rect 295379 386956 295380 387020
rect 295444 386956 295445 387020
rect 295379 386955 295445 386956
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 291883 233884 291949 233885
rect 291883 233820 291884 233884
rect 291948 233820 291949 233884
rect 291883 233819 291949 233820
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 287283 215932 287349 215933
rect 287283 215868 287284 215932
rect 287348 215868 287349 215932
rect 287283 215867 287349 215868
rect 287099 104956 287165 104957
rect 287099 104892 287100 104956
rect 287164 104892 287165 104956
rect 287099 104891 287165 104892
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 268515 102372 268581 102373
rect 268515 102308 268516 102372
rect 268580 102308 268581 102372
rect 268515 102307 268581 102308
rect 268518 101965 268578 102307
rect 268515 101964 268581 101965
rect 268515 101900 268516 101964
rect 268580 101900 268581 101964
rect 268515 101899 268581 101900
rect 281579 99380 281645 99381
rect 281579 99316 281580 99380
rect 281644 99316 281645 99380
rect 281579 99315 281645 99316
rect 279371 98292 279437 98293
rect 279371 98290 279372 98292
rect 278822 98230 279372 98290
rect 271794 93454 272414 94000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 268331 4044 268397 4045
rect 268331 3980 268332 4044
rect 268396 3980 268397 4044
rect 268331 3979 268397 3980
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 94000
rect 278822 93805 278882 98230
rect 279371 98228 279372 98230
rect 279436 98228 279437 98292
rect 279371 98227 279437 98228
rect 281582 95029 281642 99315
rect 281579 95028 281645 95029
rect 281579 94964 281580 95028
rect 281644 94964 281645 95028
rect 281579 94963 281645 94964
rect 278819 93804 278885 93805
rect 278819 93740 278820 93804
rect 278884 93740 278885 93804
rect 278819 93739 278885 93740
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 94000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 104058
rect 287286 102645 287346 215867
rect 288387 208996 288453 208997
rect 288387 208932 288388 208996
rect 288452 208932 288453 208996
rect 288387 208931 288453 208932
rect 288390 128757 288450 208931
rect 289794 183454 290414 218898
rect 290595 197980 290661 197981
rect 290595 197916 290596 197980
rect 290660 197916 290661 197980
rect 290595 197915 290661 197916
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 288571 177444 288637 177445
rect 288571 177380 288572 177444
rect 288636 177380 288637 177444
rect 288571 177379 288637 177380
rect 288574 171189 288634 177379
rect 288571 171188 288637 171189
rect 288571 171124 288572 171188
rect 288636 171124 288637 171188
rect 288571 171123 288637 171124
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 288387 128756 288453 128757
rect 288387 128692 288388 128756
rect 288452 128692 288453 128756
rect 288387 128691 288453 128692
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 287283 102644 287349 102645
rect 287283 102580 287284 102644
rect 287348 102580 287349 102644
rect 287283 102579 287349 102580
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 75454 290414 110898
rect 290598 110533 290658 197915
rect 291699 177308 291765 177309
rect 291699 177244 291700 177308
rect 291764 177244 291765 177308
rect 291699 177243 291765 177244
rect 290595 110532 290661 110533
rect 290595 110468 290596 110532
rect 290660 110468 290661 110532
rect 290595 110467 290661 110468
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 291702 31109 291762 177243
rect 291886 120189 291946 233819
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293171 218652 293237 218653
rect 293171 218588 293172 218652
rect 293236 218588 293237 218652
rect 293171 218587 293237 218588
rect 291883 120188 291949 120189
rect 291883 120124 291884 120188
rect 291948 120124 291949 120188
rect 291883 120123 291949 120124
rect 293174 111893 293234 218587
rect 293514 187174 294134 222618
rect 294459 220148 294525 220149
rect 294459 220084 294460 220148
rect 294524 220084 294525 220148
rect 294459 220083 294525 220084
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 294462 131069 294522 220083
rect 294459 131068 294525 131069
rect 294459 131004 294460 131068
rect 294524 131004 294525 131068
rect 294459 131003 294525 131004
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293171 111892 293237 111893
rect 293171 111828 293172 111892
rect 293236 111828 293237 111892
rect 293171 111827 293237 111828
rect 293514 79174 294134 114618
rect 295382 87005 295442 386955
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 305499 388380 305565 388381
rect 305499 388316 305500 388380
rect 305564 388316 305565 388380
rect 305499 388315 305565 388316
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 299611 370564 299677 370565
rect 299611 370500 299612 370564
rect 299676 370500 299677 370564
rect 299611 370499 299677 370500
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 298691 272508 298757 272509
rect 298691 272444 298692 272508
rect 298756 272444 298757 272508
rect 298691 272443 298757 272444
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 295931 211852 295997 211853
rect 295931 211788 295932 211852
rect 295996 211788 295997 211852
rect 295931 211787 295997 211788
rect 295934 98021 295994 211787
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 298139 189684 298205 189685
rect 298139 189620 298140 189684
rect 298204 189620 298205 189684
rect 298139 189619 298205 189620
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 295931 98020 295997 98021
rect 295931 97956 295932 98020
rect 295996 97956 295997 98020
rect 295931 97955 295997 97956
rect 295379 87004 295445 87005
rect 295379 86940 295380 87004
rect 295444 86940 295445 87004
rect 295379 86939 295445 86940
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 291699 31108 291765 31109
rect 291699 31044 291700 31108
rect 291764 31044 291765 31108
rect 291699 31043 291765 31044
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 295382 3501 295442 86939
rect 297234 82894 297854 118338
rect 298142 109173 298202 189619
rect 298694 122773 298754 272443
rect 298691 122772 298757 122773
rect 298691 122708 298692 122772
rect 298756 122708 298757 122772
rect 298691 122707 298757 122708
rect 298139 109172 298205 109173
rect 298139 109108 298140 109172
rect 298204 109108 298205 109172
rect 298139 109107 298205 109108
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 299614 66877 299674 370499
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 304211 282164 304277 282165
rect 304211 282100 304212 282164
rect 304276 282100 304277 282164
rect 304211 282099 304277 282100
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 302739 262852 302805 262853
rect 302739 262788 302740 262852
rect 302804 262788 302805 262852
rect 302739 262787 302805 262788
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 302742 113253 302802 262787
rect 302739 113252 302805 113253
rect 302739 113188 302740 113252
rect 302804 113188 302805 113252
rect 302739 113187 302805 113188
rect 304214 104957 304274 282099
rect 305502 134469 305562 388315
rect 306419 386476 306485 386477
rect 306419 386412 306420 386476
rect 306484 386412 306485 386476
rect 306419 386411 306485 386412
rect 306235 140044 306301 140045
rect 306235 139980 306236 140044
rect 306300 139980 306301 140044
rect 306235 139979 306301 139980
rect 305499 134468 305565 134469
rect 305499 134404 305500 134468
rect 305564 134404 305565 134468
rect 305499 134403 305565 134404
rect 304211 104956 304277 104957
rect 304211 104892 304212 104956
rect 304276 104892 304277 104956
rect 304211 104891 304277 104892
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 299611 66876 299677 66877
rect 299611 66812 299612 66876
rect 299676 66812 299677 66876
rect 299611 66811 299677 66812
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 295379 3500 295445 3501
rect 295379 3436 295380 3500
rect 295444 3436 295445 3500
rect 295379 3435 295445 3436
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 -4186 297854 10338
rect 299614 3501 299674 66811
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 299611 3500 299677 3501
rect 299611 3436 299612 3500
rect 299676 3436 299677 3500
rect 299611 3435 299677 3436
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 306238 3501 306298 139979
rect 306422 8261 306482 386411
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 309179 311132 309245 311133
rect 309179 311068 309180 311132
rect 309244 311068 309245 311132
rect 309179 311067 309245 311068
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 309182 49061 309242 311067
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 309179 49060 309245 49061
rect 309179 48996 309180 49060
rect 309244 48996 309245 49060
rect 309179 48995 309245 48996
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 306419 8260 306485 8261
rect 306419 8196 306420 8260
rect 306484 8196 306485 8260
rect 306419 8195 306485 8196
rect 306235 3500 306301 3501
rect 306235 3436 306236 3500
rect 306300 3436 306301 3500
rect 306235 3435 306301 3436
rect 307794 -1306 308414 20898
rect 309182 11797 309242 48995
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 309179 11796 309245 11797
rect 309179 11732 309180 11796
rect 309244 11732 309245 11796
rect 309179 11731 309245 11732
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 177600 348134 204618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 349107 188324 349173 188325
rect 349107 188260 349108 188324
rect 349172 188260 349173 188324
rect 349107 188259 349173 188260
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 349110 120189 349170 188259
rect 351234 177600 351854 208338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 177600 355574 212058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 177600 362414 182898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 177600 366134 186618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 177600 369854 190338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 177600 373574 194058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 177600 380414 200898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 177600 384134 204618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 177600 387854 208338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 177600 391574 212058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 177600 398414 182898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 177600 402134 186618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 177600 405854 190338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 177600 409574 194058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 177600 416414 200898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 177600 420134 204618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 177600 423854 208338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 436139 701724 436205 701725
rect 436139 701660 436140 701724
rect 436204 701660 436205 701724
rect 436139 701659 436205 701660
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 430619 258772 430685 258773
rect 430619 258708 430620 258772
rect 430684 258708 430685 258772
rect 430619 258707 430685 258708
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 427859 240820 427925 240821
rect 427859 240756 427860 240820
rect 427924 240756 427925 240820
rect 427859 240755 427925 240756
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 177600 427574 212058
rect 369568 165454 369888 165486
rect 369568 165218 369610 165454
rect 369846 165218 369888 165454
rect 369568 165134 369888 165218
rect 369568 164898 369610 165134
rect 369846 164898 369888 165134
rect 369568 164866 369888 164898
rect 400288 165454 400608 165486
rect 400288 165218 400330 165454
rect 400566 165218 400608 165454
rect 400288 165134 400608 165218
rect 400288 164898 400330 165134
rect 400566 164898 400608 165134
rect 400288 164866 400608 164898
rect 354208 147454 354528 147486
rect 354208 147218 354250 147454
rect 354486 147218 354528 147454
rect 354208 147134 354528 147218
rect 354208 146898 354250 147134
rect 354486 146898 354528 147134
rect 354208 146866 354528 146898
rect 384928 147454 385248 147486
rect 384928 147218 384970 147454
rect 385206 147218 385248 147454
rect 384928 147134 385248 147218
rect 384928 146898 384970 147134
rect 385206 146898 385248 147134
rect 384928 146866 385248 146898
rect 415648 147454 415968 147486
rect 415648 147218 415690 147454
rect 415926 147218 415968 147454
rect 415648 147134 415968 147218
rect 415648 146898 415690 147134
rect 415926 146898 415968 147134
rect 415648 146866 415968 146898
rect 369568 129454 369888 129486
rect 369568 129218 369610 129454
rect 369846 129218 369888 129454
rect 369568 129134 369888 129218
rect 369568 128898 369610 129134
rect 369846 128898 369888 129134
rect 369568 128866 369888 128898
rect 400288 129454 400608 129486
rect 400288 129218 400330 129454
rect 400566 129218 400608 129454
rect 400288 129134 400608 129218
rect 400288 128898 400330 129134
rect 400566 128898 400608 129134
rect 400288 128866 400608 128898
rect 427862 128349 427922 240755
rect 429147 206276 429213 206277
rect 429147 206212 429148 206276
rect 429212 206212 429213 206276
rect 429147 206211 429213 206212
rect 427859 128348 427925 128349
rect 427859 128284 427860 128348
rect 427924 128284 427925 128348
rect 427859 128283 427925 128284
rect 429150 126989 429210 206211
rect 430622 130797 430682 258707
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 430803 168876 430869 168877
rect 430803 168812 430804 168876
rect 430868 168812 430869 168876
rect 430803 168811 430869 168812
rect 430619 130796 430685 130797
rect 430619 130732 430620 130796
rect 430684 130732 430685 130796
rect 430619 130731 430685 130732
rect 429147 126988 429213 126989
rect 429147 126924 429148 126988
rect 429212 126924 429213 126988
rect 429147 126923 429213 126924
rect 349107 120188 349173 120189
rect 349107 120124 349108 120188
rect 349172 120124 349173 120188
rect 349107 120123 349173 120124
rect 354208 111454 354528 111486
rect 354208 111218 354250 111454
rect 354486 111218 354528 111454
rect 354208 111134 354528 111218
rect 354208 110898 354250 111134
rect 354486 110898 354528 111134
rect 354208 110866 354528 110898
rect 384928 111454 385248 111486
rect 384928 111218 384970 111454
rect 385206 111218 385248 111454
rect 384928 111134 385248 111218
rect 384928 110898 384970 111134
rect 385206 110898 385248 111134
rect 384928 110866 385248 110898
rect 415648 111454 415968 111486
rect 415648 111218 415690 111454
rect 415926 111218 415968 111454
rect 415648 111134 415968 111218
rect 415648 110898 415690 111134
rect 415926 110898 415968 111134
rect 415648 110866 415968 110898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 61174 348134 94000
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 64894 351854 94000
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 68614 355574 94000
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 75454 362414 94000
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 79174 366134 94000
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 82894 369854 94000
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 86614 373574 94000
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 93454 380414 94000
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 61174 384134 94000
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 64894 387854 94000
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 68614 391574 94000
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 75454 398414 94000
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 79174 402134 94000
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 82894 405854 94000
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 86614 409574 94000
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 93454 416414 94000
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 61174 420134 94000
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 64894 423854 94000
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 68614 427574 94000
rect 430806 90405 430866 168811
rect 433794 147454 434414 182898
rect 435035 176084 435101 176085
rect 435035 176020 435036 176084
rect 435100 176020 435101 176084
rect 435035 176019 435101 176020
rect 434851 171188 434917 171189
rect 434851 171124 434852 171188
rect 434916 171124 434917 171188
rect 434851 171123 434917 171124
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 430803 90404 430869 90405
rect 430803 90340 430804 90404
rect 430868 90340 430869 90404
rect 430803 90339 430869 90340
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 434854 47565 434914 171123
rect 435038 165069 435098 176019
rect 435035 165068 435101 165069
rect 435035 165004 435036 165068
rect 435100 165004 435101 165068
rect 435035 165003 435101 165004
rect 436142 107949 436202 701659
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 436139 107948 436205 107949
rect 436139 107884 436140 107948
rect 436204 107884 436205 107948
rect 436139 107883 436205 107884
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 434851 47564 434917 47565
rect 434851 47500 434852 47564
rect 434916 47500 434917 47564
rect 434851 47499 434917 47500
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 76618 579218 76854 579454
rect 76618 578898 76854 579134
rect 87882 579218 88118 579454
rect 87882 578898 88118 579134
rect 99146 579218 99382 579454
rect 99146 578898 99382 579134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 82250 561218 82486 561454
rect 82250 560898 82486 561134
rect 93514 561218 93750 561454
rect 93514 560898 93750 561134
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 76618 543218 76854 543454
rect 76618 542898 76854 543134
rect 87882 543218 88118 543454
rect 87882 542898 88118 543134
rect 99146 543218 99382 543454
rect 99146 542898 99382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 75618 471218 75854 471454
rect 75618 470898 75854 471134
rect 84882 471218 85118 471454
rect 84882 470898 85118 471134
rect 94146 471218 94382 471454
rect 94146 470898 94382 471134
rect 80250 453218 80486 453454
rect 80250 452898 80486 453134
rect 89514 453218 89750 453454
rect 89514 452898 89750 453134
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 89610 381218 89846 381454
rect 89610 380898 89846 381134
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 74250 363218 74486 363454
rect 74250 362898 74486 363134
rect 104970 363218 105206 363454
rect 104970 362898 105206 363134
rect 89610 345218 89846 345454
rect 89610 344898 89846 345134
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 89610 273218 89846 273454
rect 89610 272898 89846 273134
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 221249 165218 221485 165454
rect 221249 164898 221485 165134
rect 224513 165218 224749 165454
rect 224513 164898 224749 165134
rect 219617 147218 219853 147454
rect 219617 146898 219853 147134
rect 222881 147218 223117 147454
rect 222881 146898 223117 147134
rect 226145 147218 226381 147454
rect 226145 146898 226381 147134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 221249 129218 221485 129454
rect 221249 128898 221485 129134
rect 224513 129218 224749 129454
rect 224513 128898 224749 129134
rect 219617 111218 219853 111454
rect 219617 110898 219853 111134
rect 222881 111218 223117 111454
rect 222881 110898 223117 111134
rect 226145 111218 226381 111454
rect 226145 110898 226381 111134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 272249 165218 272485 165454
rect 272249 164898 272485 165134
rect 275513 165218 275749 165454
rect 275513 164898 275749 165134
rect 270617 147218 270853 147454
rect 270617 146898 270853 147134
rect 273881 147218 274117 147454
rect 273881 146898 274117 147134
rect 277145 147218 277381 147454
rect 277145 146898 277381 147134
rect 272249 129218 272485 129454
rect 272249 128898 272485 129134
rect 275513 129218 275749 129454
rect 275513 128898 275749 129134
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 270617 111218 270853 111454
rect 270617 110898 270853 111134
rect 273881 111218 274117 111454
rect 273881 110898 274117 111134
rect 277145 111218 277381 111454
rect 277145 110898 277381 111134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 369610 165218 369846 165454
rect 369610 164898 369846 165134
rect 400330 165218 400566 165454
rect 400330 164898 400566 165134
rect 354250 147218 354486 147454
rect 354250 146898 354486 147134
rect 384970 147218 385206 147454
rect 384970 146898 385206 147134
rect 415690 147218 415926 147454
rect 415690 146898 415926 147134
rect 369610 129218 369846 129454
rect 369610 128898 369846 129134
rect 400330 129218 400566 129454
rect 400330 128898 400566 129134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 354250 111218 354486 111454
rect 354250 110898 354486 111134
rect 384970 111218 385206 111454
rect 384970 110898 385206 111134
rect 415690 111218 415926 111454
rect 415690 110898 415926 111134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 76618 579454
rect 76854 579218 87882 579454
rect 88118 579218 99146 579454
rect 99382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 76618 579134
rect 76854 578898 87882 579134
rect 88118 578898 99146 579134
rect 99382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 82250 561454
rect 82486 561218 93514 561454
rect 93750 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 82250 561134
rect 82486 560898 93514 561134
rect 93750 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 76618 543454
rect 76854 543218 87882 543454
rect 88118 543218 99146 543454
rect 99382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 76618 543134
rect 76854 542898 87882 543134
rect 88118 542898 99146 543134
rect 99382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 75618 471454
rect 75854 471218 84882 471454
rect 85118 471218 94146 471454
rect 94382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 75618 471134
rect 75854 470898 84882 471134
rect 85118 470898 94146 471134
rect 94382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 80250 453454
rect 80486 453218 89514 453454
rect 89750 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 80250 453134
rect 80486 452898 89514 453134
rect 89750 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 89610 381454
rect 89846 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 89610 381134
rect 89846 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 74250 363454
rect 74486 363218 104970 363454
rect 105206 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 74250 363134
rect 74486 362898 104970 363134
rect 105206 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 89610 345454
rect 89846 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 89610 345134
rect 89846 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 89610 273454
rect 89846 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 89610 273134
rect 89846 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 221249 165454
rect 221485 165218 224513 165454
rect 224749 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 272249 165454
rect 272485 165218 275513 165454
rect 275749 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 369610 165454
rect 369846 165218 400330 165454
rect 400566 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 221249 165134
rect 221485 164898 224513 165134
rect 224749 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 272249 165134
rect 272485 164898 275513 165134
rect 275749 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 369610 165134
rect 369846 164898 400330 165134
rect 400566 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 219617 147454
rect 219853 147218 222881 147454
rect 223117 147218 226145 147454
rect 226381 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 270617 147454
rect 270853 147218 273881 147454
rect 274117 147218 277145 147454
rect 277381 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 354250 147454
rect 354486 147218 384970 147454
rect 385206 147218 415690 147454
rect 415926 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 219617 147134
rect 219853 146898 222881 147134
rect 223117 146898 226145 147134
rect 226381 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 270617 147134
rect 270853 146898 273881 147134
rect 274117 146898 277145 147134
rect 277381 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 354250 147134
rect 354486 146898 384970 147134
rect 385206 146898 415690 147134
rect 415926 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 221249 129454
rect 221485 129218 224513 129454
rect 224749 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 272249 129454
rect 272485 129218 275513 129454
rect 275749 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 369610 129454
rect 369846 129218 400330 129454
rect 400566 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 221249 129134
rect 221485 128898 224513 129134
rect 224749 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 272249 129134
rect 272485 128898 275513 129134
rect 275749 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 369610 129134
rect 369846 128898 400330 129134
rect 400566 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 219617 111454
rect 219853 111218 222881 111454
rect 223117 111218 226145 111454
rect 226381 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 270617 111454
rect 270853 111218 273881 111454
rect 274117 111218 277145 111454
rect 277381 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 354250 111454
rect 354486 111218 384970 111454
rect 385206 111218 415690 111454
rect 415926 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 219617 111134
rect 219853 110898 222881 111134
rect 223117 110898 226145 111134
rect 226381 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 270617 111134
rect 270853 110898 273881 111134
rect 274117 110898 277145 111134
rect 277381 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 354250 111134
rect 354486 110898 384970 111134
rect 385206 110898 415690 111134
rect 415926 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 268000 0 1 96000
box 0 0 12000 79688
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 12000 79688
use wrapped_frequency_counter  wrapped_frequency_counter_2
timestamp 0
transform 1 0 70000 0 1 440000
box -10 -52 30000 50000
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
use wrapped_hack_soc_dffram  wrapped_hack_soc_dffram_11
timestamp 0
transform 1 0 350000 0 1 96000
box 0 0 78450 79600
use wrapped_rgb_mixer  wrapped_rgb_mixer_3
timestamp 0
transform 1 0 70000 0 1 540000
box -10 -52 36000 42000
use wrapped_vga_clock  wrapped_vga_clock_1
timestamp 0
transform 1 0 70000 0 1 340000
box -10 -52 46000 46000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 294000 74414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 294000 110414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 388000 74414 438000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 492000 74414 538000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 584000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 388000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 177600 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 177600 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 294000 78134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 294000 114134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 388000 78134 438000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 492000 78134 538000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 584000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 388000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 177600 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 177600 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 294000 81854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 294000 117854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 388000 81854 438000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 492000 81854 538000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 584000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 388000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 177600 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 177600 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 294000 85574 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 388000 85574 438000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 492000 85574 538000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 584000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 294000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 177600 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 177600 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 294000 99854 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 388000 99854 438000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 492000 99854 538000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 584000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 178000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 177600 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 177600 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 177600 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 294000 103574 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 388000 103574 538000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 584000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 177600 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 177600 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 177600 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 294000 92414 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 388000 92414 438000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 492000 92414 538000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 584000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 178000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 177600 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 177600 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 294000 96134 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 388000 96134 438000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 492000 96134 538000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 584000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 178000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 177600 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 177600 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 177600 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
